module real_jpeg_25634_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_292;
wire n_215;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_255;
wire n_243;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_293;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_305;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_240;
wire n_55;
wire n_185;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_295;
wire n_167;
wire n_213;
wire n_179;
wire n_133;
wire n_202;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_23),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_62),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_2),
.A2(n_54),
.B1(n_56),
.B2(n_62),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_2),
.A2(n_62),
.B1(n_75),
.B2(n_76),
.Y(n_197)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_15),
.B(n_304),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_4),
.B(n_305),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_6),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_8),
.A2(n_21),
.B1(n_24),
.B2(n_27),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_8),
.A2(n_27),
.B1(n_33),
.B2(n_35),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_8),
.A2(n_27),
.B1(n_54),
.B2(n_56),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_8),
.A2(n_27),
.B1(n_75),
.B2(n_76),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_9),
.A2(n_21),
.B1(n_24),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_9),
.A2(n_37),
.B1(n_54),
.B2(n_56),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_37),
.B1(n_75),
.B2(n_76),
.Y(n_91)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_10),
.A2(n_11),
.B1(n_21),
.B2(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_44),
.B1(n_54),
.B2(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_11),
.A2(n_33),
.B1(n_35),
.B2(n_44),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_11),
.A2(n_44),
.B1(n_75),
.B2(n_76),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_11),
.B(n_31),
.C(n_35),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_11),
.B(n_32),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_11),
.B(n_51),
.C(n_54),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_11),
.B(n_72),
.C(n_75),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_11),
.B(n_13),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_11),
.B(n_106),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_11),
.B(n_65),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_13),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_13),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_297),
.B(n_301),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_78),
.B(n_296),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_38),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_18),
.B(n_38),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_18),
.B(n_298),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_18),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_28),
.B1(n_32),
.B2(n_36),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_20),
.A2(n_41),
.B(n_42),
.Y(n_40)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_22),
.B(n_193),
.Y(n_192)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_28),
.A2(n_32),
.B1(n_43),
.B2(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_28),
.B(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

AO22x1_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_33),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_35),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx6p67_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_35),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_36),
.B(n_300),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_39),
.B(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_39),
.B(n_294),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_45),
.CI(n_57),
.CON(n_39),
.SN(n_39)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_41),
.A2(n_42),
.B(n_60),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_49),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_48),
.A2(n_53),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_49),
.A2(n_65),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_49),
.B(n_111),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

OA22x2_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_53),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_53),
.A2(n_110),
.B(n_121),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_54),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_56),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_54),
.B(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.C(n_66),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_SL g128 ( 
.A(n_58),
.B(n_129),
.C(n_137),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_58),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_58),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_58),
.A2(n_137),
.B1(n_138),
.B2(n_151),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_58),
.A2(n_108),
.B1(n_151),
.B2(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_58),
.B(n_108),
.C(n_190),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_63),
.A2(n_66),
.B1(n_118),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_63),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_66),
.A2(n_118),
.B1(n_119),
.B2(n_122),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_66),
.B(n_114),
.C(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_77),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_68),
.B(n_96),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_70),
.A2(n_96),
.B1(n_106),
.B2(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_74),
.A2(n_95),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_75),
.B(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_293),
.B(n_295),
.Y(n_78)
);

OAI211xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_139),
.B(n_153),
.C(n_292),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_123),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_81),
.B(n_123),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_101),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_103),
.C(n_112),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_92),
.B(n_97),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_83),
.A2(n_97),
.B1(n_98),
.B2(n_126),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_83),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_83),
.A2(n_93),
.B1(n_126),
.B2(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_85),
.B(n_198),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_86),
.A2(n_91),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_86),
.B(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_86),
.Y(n_196)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_92),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_93),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_99),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_112),
.B2(n_113),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_104),
.B(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_108),
.B(n_210),
.C(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_108),
.A2(n_200),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_111),
.Y(n_173)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_115),
.B1(n_147),
.B2(n_152),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_114),
.B(n_137),
.C(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_114),
.A2(n_115),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_114),
.A2(n_115),
.B1(n_172),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_163),
.C(n_172),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_115),
.B(n_143),
.C(n_147),
.Y(n_294)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.C(n_128),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_127),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_130),
.A2(n_134),
.B1(n_135),
.B2(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_130),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_134),
.A2(n_135),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_134),
.A2(n_135),
.B1(n_223),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_135),
.B(n_217),
.C(n_223),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_135),
.B(n_195),
.C(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_137),
.A2(n_138),
.B1(n_186),
.B2(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_137),
.A2(n_138),
.B1(n_170),
.B2(n_183),
.Y(n_260)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_138),
.B(n_170),
.C(n_261),
.Y(n_264)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_SL g153 ( 
.A(n_140),
.B(n_154),
.C(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_141),
.B(n_142),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_176),
.B(n_291),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_174),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_157),
.B(n_174),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_158),
.B(n_160),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_162),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_163),
.A2(n_164),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_170),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_168),
.A2(n_197),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_170),
.A2(n_183),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_170),
.B(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_172),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_286),
.B(n_290),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_213),
.B(n_272),
.C(n_285),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_202),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_179),
.B(n_202),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_189),
.B2(n_201),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_182),
.B(n_188),
.C(n_201),
.Y(n_273)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_199),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_194),
.A2(n_195),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_246),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.C(n_209),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_204),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_209),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_210),
.A2(n_212),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_210),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_212),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_271),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_232),
.B(n_270),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_229),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_216),
.B(n_229),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_217),
.A2(n_218),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_222),
.B(n_237),
.Y(n_248)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_263),
.B(n_269),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_257),
.B(n_262),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_249),
.B(n_256),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_241),
.B(n_248),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_238),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_245),
.B(n_247),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_250),
.B(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_258),
.B(n_259),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_264),
.B(n_265),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_266),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_274),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_284),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_281),
.B2(n_282),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_282),
.C(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_288),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);


endmodule