module fake_jpeg_4733_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_18),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_19),
.B(n_21),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_48),
.A2(n_21),
.B(n_19),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_51),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_62),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_28),
.B1(n_31),
.B2(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_57),
.A2(n_30),
.B1(n_24),
.B2(n_17),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_58),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_32),
.C(n_34),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_18),
.C(n_27),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_36),
.A2(n_28),
.B1(n_33),
.B2(n_26),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_28),
.B1(n_33),
.B2(n_18),
.Y(n_74)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_86),
.Y(n_124)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_78),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_28),
.B1(n_36),
.B2(n_40),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_81),
.B1(n_82),
.B2(n_88),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_38),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_76),
.B(n_47),
.Y(n_107)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_38),
.B1(n_36),
.B2(n_40),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_33),
.B1(n_34),
.B2(n_27),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_92),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_44),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_51),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_24),
.B1(n_52),
.B2(n_53),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_17),
.B1(n_30),
.B2(n_32),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_96),
.A2(n_24),
.B1(n_32),
.B2(n_53),
.Y(n_102)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_104),
.B1(n_98),
.B2(n_87),
.Y(n_133)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_53),
.B1(n_47),
.B2(n_70),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_107),
.A2(n_99),
.B(n_89),
.Y(n_156)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_112),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_116),
.B1(n_118),
.B2(n_122),
.Y(n_132)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_117),
.Y(n_138)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_115),
.Y(n_149)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_47),
.B1(n_52),
.B2(n_43),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_68),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_37),
.B1(n_43),
.B2(n_35),
.Y(n_118)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_37),
.B1(n_43),
.B2(n_35),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_81),
.A2(n_43),
.B1(n_29),
.B2(n_35),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_122),
.B1(n_118),
.B2(n_121),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_77),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_145),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_90),
.B(n_77),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_129),
.A2(n_141),
.B(n_143),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_81),
.B1(n_101),
.B2(n_76),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_114),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_76),
.B1(n_86),
.B2(n_91),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_143),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_75),
.B1(n_98),
.B2(n_87),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_154),
.B1(n_112),
.B2(n_23),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_75),
.B1(n_74),
.B2(n_88),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_151),
.B1(n_153),
.B2(n_123),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_74),
.B(n_84),
.C(n_96),
.D(n_71),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_22),
.C(n_19),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_82),
.B1(n_96),
.B2(n_84),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_23),
.B(n_20),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_85),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_102),
.B(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_147),
.Y(n_191)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_85),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_94),
.B1(n_78),
.B2(n_73),
.Y(n_153)
);

AO22x1_ASAP7_75t_SL g154 ( 
.A1(n_100),
.A2(n_79),
.B1(n_54),
.B2(n_67),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_103),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_22),
.B(n_19),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_109),
.B(n_89),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_157),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_68),
.C(n_58),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_58),
.Y(n_168)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_164),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_21),
.B(n_72),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_160),
.A2(n_165),
.B(n_175),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_161),
.A2(n_186),
.B1(n_29),
.B2(n_62),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_21),
.B(n_22),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_179),
.B1(n_132),
.B2(n_151),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_170),
.C(n_144),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_136),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_173),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_56),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_22),
.B(n_21),
.C(n_19),
.Y(n_175)
);

OAI31xp33_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_21),
.A3(n_20),
.B(n_35),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_178),
.B(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_182),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_145),
.B1(n_133),
.B2(n_158),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_0),
.B(n_1),
.Y(n_207)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_128),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_152),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_129),
.A2(n_22),
.B(n_19),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_56),
.B1(n_20),
.B2(n_29),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_155),
.B(n_147),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_22),
.B(n_20),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_189),
.A2(n_190),
.B(n_29),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_152),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_192),
.A2(n_175),
.B(n_162),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_210),
.C(n_167),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_202),
.B1(n_213),
.B2(n_219),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_0),
.Y(n_242)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_186),
.A2(n_140),
.B1(n_132),
.B2(n_139),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_184),
.B(n_190),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_218),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_138),
.C(n_142),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_67),
.B1(n_62),
.B2(n_54),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_164),
.B1(n_182),
.B2(n_177),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_54),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_215),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_8),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_220),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_8),
.B(n_15),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_161),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_245),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_238),
.C(n_209),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_174),
.B(n_173),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_225),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_189),
.B(n_160),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_168),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_236),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_197),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_233),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_180),
.B1(n_159),
.B2(n_165),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_232),
.A2(n_242),
.B1(n_217),
.B2(n_220),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_234),
.A2(n_2),
.B(n_3),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_180),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_243),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_163),
.C(n_169),
.Y(n_238)
);

INVxp33_ASAP7_75t_SL g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_162),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_196),
.Y(n_261)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_246),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_9),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_263),
.C(n_225),
.Y(n_273)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_202),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_251),
.A2(n_267),
.B(n_234),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_198),
.B1(n_206),
.B2(n_216),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_244),
.A2(n_201),
.B1(n_193),
.B2(n_200),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_254),
.A2(n_235),
.B1(n_9),
.B2(n_10),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_257),
.A2(n_3),
.B(n_4),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_214),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_261),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_192),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_266),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_193),
.C(n_192),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_238),
.B(n_212),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_224),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_257),
.B(n_254),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_251),
.B(n_226),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_227),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_279),
.C(n_280),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_260),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_274),
.Y(n_293)
);

NAND4xp25_ASAP7_75t_SL g276 ( 
.A(n_253),
.B(n_228),
.C(n_230),
.D(n_232),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_221),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_223),
.C(n_235),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_259),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_284),
.B(n_247),
.Y(n_290)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_9),
.Y(n_283)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_268),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_290),
.B(n_251),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

INVxp33_ASAP7_75t_SL g305 ( 
.A(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_259),
.C(n_263),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_258),
.C(n_255),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_255),
.C(n_265),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_269),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_299),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_293),
.A3(n_285),
.B1(n_298),
.B2(n_295),
.C1(n_291),
.C2(n_297),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_302),
.C(n_303),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_270),
.B1(n_279),
.B2(n_273),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_278),
.C(n_280),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_282),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_304),
.A2(n_306),
.B(n_286),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_292),
.C(n_294),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_277),
.B1(n_262),
.B2(n_12),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_310),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_11),
.B(n_13),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_285),
.B(n_11),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_290),
.B(n_11),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_318),
.B(n_16),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_16),
.C(n_6),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_305),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_315),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_4),
.Y(n_317)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_317),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_305),
.A2(n_12),
.B(n_13),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_316),
.A2(n_301),
.B1(n_309),
.B2(n_12),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_323),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_314),
.B(n_309),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_324),
.B(n_312),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_319),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_327),
.Y(n_329)
);

AOI322xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_322),
.A3(n_328),
.B1(n_16),
.B2(n_7),
.C1(n_5),
.C2(n_6),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_7),
.B(n_308),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_7),
.Y(n_332)
);


endmodule