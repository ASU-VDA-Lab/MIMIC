module fake_jpeg_25169_n_180 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_2),
.B(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g41 ( 
.A(n_27),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_28),
.B(n_30),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_51),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_38),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_57),
.Y(n_62)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_71),
.B1(n_28),
.B2(n_19),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_16),
.B1(n_41),
.B2(n_17),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_60),
.A2(n_65),
.B1(n_72),
.B2(n_29),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_30),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_67),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_38),
.C(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_77),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_17),
.B1(n_23),
.B2(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_75),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_79),
.B(n_81),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_20),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_40),
.C(n_27),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_19),
.C(n_29),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_81),
.CON(n_92),
.SN(n_92)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_15),
.B(n_26),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_29),
.B(n_19),
.C(n_23),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_81),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_103),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_15),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_65),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_63),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_18),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_24),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_76),
.B1(n_71),
.B2(n_65),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_115),
.B1(n_121),
.B2(n_96),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_90),
.Y(n_127)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_88),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_78),
.B1(n_81),
.B2(n_63),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_64),
.B1(n_20),
.B2(n_3),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_85),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_131),
.B1(n_123),
.B2(n_115),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_104),
.C(n_91),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_127),
.C(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_132),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_85),
.C(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_133),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_111),
.C(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_99),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_115),
.C(n_84),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_116),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_84),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_118),
.B1(n_108),
.B2(n_113),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_112),
.B1(n_103),
.B2(n_100),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_110),
.B1(n_113),
.B2(n_108),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_139),
.B1(n_147),
.B2(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_148),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_125),
.C(n_86),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_135),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_155),
.B(n_158),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_98),
.C(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_157),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_9),
.B(n_14),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_95),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_145),
.B(n_10),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_140),
.B(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_160),
.C(n_163),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_142),
.B(n_141),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_154),
.A2(n_141),
.B(n_100),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_1),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_1),
.C(n_2),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_154),
.B1(n_152),
.B2(n_151),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_164),
.B(n_7),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_167),
.B(n_170),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_169),
.B(n_3),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_98),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_172),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_170),
.C(n_5),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_6),
.B(n_4),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_173),
.B(n_5),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_178),
.B(n_4),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_5),
.Y(n_180)
);


endmodule