module fake_jpeg_22090_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_5),
.B(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_18),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_27),
.B1(n_25),
.B2(n_19),
.Y(n_49)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_31),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_60),
.B1(n_20),
.B2(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_52),
.B(n_63),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_27),
.B1(n_18),
.B2(n_26),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_40),
.B1(n_33),
.B2(n_30),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_30),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_32),
.B1(n_25),
.B2(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_19),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_68),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_15),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_21),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_85),
.B1(n_87),
.B2(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_79),
.Y(n_110)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_69),
.B(n_61),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_37),
.B1(n_2),
.B2(n_4),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_50),
.B1(n_66),
.B2(n_51),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_48),
.B(n_0),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_0),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_105),
.B(n_94),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_107),
.B1(n_82),
.B2(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_66),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_112),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_109),
.B(n_78),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_91),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_72),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_131),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_129),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_80),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_120),
.B(n_125),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_80),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_121),
.C(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_73),
.C(n_83),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_79),
.C(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_127),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_86),
.C(n_95),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_124),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_135),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_107),
.B(n_105),
.C(n_113),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_126),
.B1(n_57),
.B2(n_67),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_128),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NAND4xp25_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_81),
.C(n_84),
.D(n_108),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_138),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_96),
.C(n_97),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_13),
.B(n_14),
.Y(n_152)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_97),
.B(n_96),
.C(n_114),
.D(n_101),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_102),
.C(n_57),
.Y(n_153)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_136),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_119),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_149),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_131),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_134),
.A2(n_118),
.B1(n_101),
.B2(n_90),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_151),
.A2(n_152),
.B(n_154),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_140),
.C(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_132),
.C(n_144),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_150),
.B(n_138),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_161),
.C(n_67),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_134),
.C(n_140),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_154),
.B(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_146),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_158),
.Y(n_169)
);

NOR2x1_ASAP7_75t_SL g172 ( 
.A(n_164),
.B(n_165),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_148),
.B(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_4),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_169),
.B(n_11),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_166),
.B(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_175),
.C(n_4),
.Y(n_177)
);

AOI21x1_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_169),
.B(n_171),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_177),
.B1(n_6),
.B2(n_7),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_7),
.Y(n_179)
);


endmodule