module fake_jpeg_18545_n_35 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

AOI22xp33_ASAP7_75t_SL g8 ( 
.A1(n_6),
.A2(n_3),
.B1(n_4),
.B2(n_2),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_4),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

OR2x2_ASAP7_75t_SL g14 ( 
.A(n_2),
.B(n_1),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_0),
.C(n_1),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_20),
.C(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_12),
.B(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_3),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_10),
.C(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

XNOR2x1_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_7),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_12),
.B(n_9),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_25),
.B(n_27),
.C(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_26),
.Y(n_30)
);

AO221x1_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_21),
.B1(n_10),
.B2(n_11),
.C(n_13),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

NAND4xp25_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_31),
.C(n_28),
.D(n_25),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_18),
.B1(n_16),
.B2(n_21),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_34),
.C(n_32),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.C(n_29),
.Y(n_34)
);


endmodule