module fake_jpeg_13592_n_35 (n_3, n_2, n_1, n_0, n_4, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_SL g6 ( 
.A(n_0),
.Y(n_6)
);

INVx6_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NAND2xp33_ASAP7_75t_SL g8 ( 
.A(n_4),
.B(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_SL g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_SL g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_20),
.Y(n_26)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_1),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_6),
.A2(n_1),
.B1(n_5),
.B2(n_3),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_19),
.B1(n_22),
.B2(n_10),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_5),
.B(n_11),
.C(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_21),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_11),
.B1(n_7),
.B2(n_9),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_18),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_10),
.C(n_7),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_12),
.C(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

AOI322xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_30),
.A3(n_23),
.B1(n_31),
.B2(n_24),
.C1(n_29),
.C2(n_14),
.Y(n_33)
);

AOI21x1_ASAP7_75t_SL g34 ( 
.A1(n_33),
.A2(n_31),
.B(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_21),
.Y(n_35)
);


endmodule