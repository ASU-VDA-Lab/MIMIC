module fake_jpeg_10001_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_17),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_54),
.B(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_26),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_26),
.C(n_19),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_24),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_28),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_65),
.B(n_52),
.Y(n_109)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_78),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_29),
.B1(n_32),
.B2(n_31),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_74),
.A2(n_82),
.B1(n_90),
.B2(n_97),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_60),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_81),
.Y(n_129)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_49),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_29),
.B1(n_34),
.B2(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_84),
.Y(n_105)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_29),
.B1(n_34),
.B2(n_36),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_99),
.Y(n_117)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_62),
.B1(n_49),
.B2(n_67),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_109),
.A2(n_118),
.B(n_0),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_115),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_61),
.B1(n_50),
.B2(n_52),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_85),
.B1(n_97),
.B2(n_39),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_64),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_70),
.B(n_28),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_65),
.C(n_62),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_83),
.C(n_73),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_54),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_14),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_125),
.B1(n_95),
.B2(n_84),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_39),
.B1(n_38),
.B2(n_36),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_134),
.C(n_137),
.Y(n_165)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_133),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_81),
.C(n_62),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_101),
.C(n_43),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_74),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_148),
.C(n_149),
.Y(n_169)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_143),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_71),
.B1(n_80),
.B2(n_77),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_151),
.B1(n_103),
.B2(n_102),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_150),
.B1(n_158),
.B2(n_102),
.Y(n_176)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_152),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_45),
.C(n_44),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_33),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_89),
.B1(n_30),
.B2(n_21),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_79),
.B1(n_15),
.B2(n_16),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_157),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_35),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_127),
.C(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_130),
.A2(n_21),
.B1(n_30),
.B2(n_28),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_16),
.B(n_15),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_107),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_160),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_162),
.B(n_175),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_134),
.B1(n_137),
.B2(n_131),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_178),
.B1(n_180),
.B2(n_28),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_117),
.B(n_114),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_164),
.A2(n_171),
.B(n_174),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_168),
.A2(n_176),
.B1(n_185),
.B2(n_190),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_173),
.C(n_191),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_128),
.B(n_124),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_124),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_103),
.B(n_122),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

AO21x2_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_106),
.B(n_122),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_20),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_135),
.A2(n_106),
.B1(n_108),
.B2(n_120),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_108),
.B(n_35),
.Y(n_182)
);

XNOR2x2_ASAP7_75t_SL g207 ( 
.A(n_182),
.B(n_24),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_138),
.A2(n_116),
.B1(n_126),
.B2(n_113),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_186),
.A2(n_187),
.B(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_192),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_116),
.B1(n_113),
.B2(n_30),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_35),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_22),
.B1(n_30),
.B2(n_21),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_45),
.B(n_47),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_28),
.C(n_33),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_199),
.C(n_210),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_33),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_201),
.Y(n_241)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_20),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_203),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_205),
.A2(n_219),
.B1(n_192),
.B2(n_190),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_208),
.B1(n_193),
.B2(n_187),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_1),
.B(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_215),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_22),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_22),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_220),
.C(n_221),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_162),
.A2(n_28),
.B1(n_23),
.B2(n_20),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_23),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_23),
.C(n_20),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_223),
.Y(n_234)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_225),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_202),
.Y(n_230)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_240),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_181),
.B1(n_164),
.B2(n_176),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_235),
.A2(n_238),
.B1(n_245),
.B2(n_244),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_216),
.B1(n_225),
.B2(n_207),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_161),
.B1(n_177),
.B2(n_194),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_171),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_171),
.B(n_174),
.C(n_170),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_247),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_186),
.B1(n_174),
.B2(n_191),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_216),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_2),
.B(n_3),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_23),
.C(n_3),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_217),
.C(n_221),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_195),
.B(n_23),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_218),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_252),
.A2(n_261),
.B1(n_267),
.B2(n_246),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_256),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_263),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_251),
.C(n_226),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_259),
.C(n_265),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_198),
.C(n_220),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_235),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_210),
.B1(n_217),
.B2(n_208),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_262),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_199),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_2),
.C(n_3),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_4),
.C(n_5),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_228),
.C(n_237),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_231),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_11),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_232),
.Y(n_287)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_272),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_231),
.A2(n_4),
.B(n_7),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_254),
.B(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_269),
.B(n_227),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_274),
.B(n_267),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_276),
.A2(n_281),
.B1(n_283),
.B2(n_288),
.Y(n_293)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_230),
.C(n_243),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_282),
.C(n_255),
.Y(n_298)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_253),
.A2(n_248),
.B1(n_230),
.B2(n_243),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_229),
.C(n_233),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_259),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_287),
.B(n_9),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_242),
.B1(n_236),
.B2(n_246),
.Y(n_288)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_240),
.B(n_232),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_289),
.A2(n_232),
.B(n_261),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_271),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_260),
.B(n_252),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_291),
.A2(n_295),
.B(n_285),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_303),
.Y(n_315)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_265),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_300),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_301),
.C(n_273),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_287),
.B(n_7),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_275),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_9),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_9),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_286),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_277),
.Y(n_311)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_293),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_313),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_314),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_311),
.A2(n_299),
.B(n_12),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_282),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_275),
.C(n_11),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_316),
.B(n_305),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_10),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_10),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_309),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_291),
.Y(n_320)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_322),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_291),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_292),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_314),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_325),
.A2(n_306),
.B(n_312),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_330),
.C(n_323),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_331),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_316),
.Y(n_330)
);

XNOR2x2_ASAP7_75t_SL g333 ( 
.A(n_332),
.B(n_326),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_333),
.B(n_334),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_327),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_328),
.B(n_335),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_318),
.B(n_13),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_10),
.C(n_14),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_340),
.Y(n_341)
);


endmodule