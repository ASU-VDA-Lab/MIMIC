module fake_jpeg_30375_n_517 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_59),
.Y(n_106)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_56),
.B(n_89),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_67),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_64),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_15),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_73),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_72),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_14),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_74),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_75),
.B(n_77),
.Y(n_142)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_25),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_78),
.B(n_83),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_12),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_30),
.B(n_12),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_33),
.B(n_0),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_91),
.B(n_95),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_19),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_103),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_33),
.B(n_0),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_65),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_107),
.B(n_112),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_32),
.B1(n_37),
.B2(n_39),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_109),
.A2(n_140),
.B1(n_148),
.B2(n_157),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_47),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_113),
.B(n_30),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_58),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_137),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_62),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_138),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_32),
.B1(n_37),
.B2(n_39),
.Y(n_140)
);

BUFx16f_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_105),
.A2(n_38),
.B1(n_41),
.B2(n_31),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_101),
.A2(n_37),
.B1(n_32),
.B2(n_46),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_156),
.A2(n_43),
.B(n_71),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_169),
.B(n_183),
.Y(n_262)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_176),
.Y(n_224)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_114),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_174),
.B(n_178),
.Y(n_242)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_47),
.Y(n_176)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_106),
.B(n_46),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_121),
.A2(n_142),
.B(n_147),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_180),
.A2(n_2),
.B(n_3),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_76),
.C(n_81),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_38),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_184),
.B(n_201),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_55),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_185),
.B(n_189),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_66),
.B1(n_72),
.B2(n_60),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_196),
.B1(n_204),
.B2(n_213),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_34),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_154),
.B(n_51),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_191),
.B(n_211),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_27),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_192),
.B(n_207),
.Y(n_248)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_194),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_151),
.A2(n_93),
.B1(n_105),
.B2(n_70),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_197),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_27),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_202),
.Y(n_243)
);

NAND2x1_ASAP7_75t_L g201 ( 
.A(n_146),
.B(n_100),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_51),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_206),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_151),
.A2(n_70),
.B1(n_36),
.B2(n_49),
.Y(n_204)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_126),
.B(n_34),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_19),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_210),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_129),
.B(n_128),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_119),
.B(n_84),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_212),
.B(n_214),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_145),
.A2(n_36),
.B1(n_49),
.B2(n_31),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_129),
.B(n_41),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_215),
.B(n_217),
.Y(n_265)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_145),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_128),
.B(n_41),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_79),
.Y(n_237)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_219),
.B(n_220),
.Y(n_267)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_120),
.B1(n_125),
.B2(n_161),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_225),
.A2(n_233),
.B1(n_250),
.B2(n_268),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_172),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_226),
.B(n_227),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

OAI22x1_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_148),
.B1(n_155),
.B2(n_161),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_187),
.A2(n_110),
.B1(n_131),
.B2(n_133),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_235),
.A2(n_179),
.B1(n_195),
.B2(n_182),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_237),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_183),
.A2(n_133),
.B1(n_131),
.B2(n_61),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_239),
.A2(n_247),
.B1(n_177),
.B2(n_170),
.Y(n_278)
);

BUFx12_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_108),
.B1(n_132),
.B2(n_57),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_213),
.A2(n_120),
.B1(n_125),
.B2(n_155),
.Y(n_250)
);

AOI32xp33_ASAP7_75t_L g251 ( 
.A1(n_184),
.A2(n_88),
.A3(n_136),
.B1(n_53),
.B2(n_150),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_252),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_167),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_208),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_41),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_260),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_202),
.B(n_41),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_263),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_3),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_217),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_206),
.A2(n_136),
.B1(n_138),
.B2(n_150),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_270),
.Y(n_309)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_274),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_248),
.B(n_201),
.Y(n_274)
);

OA22x2_ASAP7_75t_SL g276 ( 
.A1(n_233),
.A2(n_204),
.B1(n_196),
.B2(n_181),
.Y(n_276)
);

OA22x2_ASAP7_75t_L g322 ( 
.A1(n_276),
.A2(n_278),
.B1(n_259),
.B2(n_244),
.Y(n_322)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_280),
.A2(n_301),
.B1(n_245),
.B2(n_265),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_293),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_257),
.A2(n_208),
.B(n_188),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_284),
.A2(n_236),
.B(n_134),
.Y(n_340)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_227),
.B(n_212),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_262),
.B(n_49),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_232),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_261),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_295),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_237),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_292),
.B(n_298),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_248),
.B(n_168),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_226),
.B(n_132),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_299),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_229),
.Y(n_297)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_234),
.B(n_216),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_249),
.A2(n_193),
.B1(n_186),
.B2(n_108),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_123),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_300),
.A2(n_188),
.B(n_232),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_249),
.A2(n_262),
.B1(n_228),
.B2(n_231),
.Y(n_301)
);

OAI32xp33_ASAP7_75t_L g302 ( 
.A1(n_228),
.A2(n_124),
.A3(n_138),
.B1(n_216),
.B2(n_7),
.Y(n_302)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_246),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_303),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_224),
.B(n_124),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_263),
.Y(n_331)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_229),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_308),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_251),
.A2(n_254),
.B1(n_230),
.B2(n_240),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_266),
.B(n_252),
.Y(n_318)
);

CKINVDCx12_ASAP7_75t_R g307 ( 
.A(n_246),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_307),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_243),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_310),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_283),
.A2(n_260),
.B1(n_258),
.B2(n_241),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_312),
.A2(n_321),
.B1(n_327),
.B2(n_342),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_285),
.B(n_242),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_314),
.B(n_336),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_242),
.C(n_269),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_308),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_318),
.A2(n_337),
.B(n_278),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_276),
.A2(n_230),
.B1(n_240),
.B2(n_255),
.Y(n_321)
);

OA22x2_ASAP7_75t_L g372 ( 
.A1(n_322),
.A2(n_271),
.B1(n_305),
.B2(n_297),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_293),
.B(n_269),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_334),
.Y(n_355)
);

OA21x2_ASAP7_75t_SL g325 ( 
.A1(n_279),
.A2(n_246),
.B(n_253),
.Y(n_325)
);

XOR2x1_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_328),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_276),
.A2(n_259),
.B1(n_244),
.B2(n_238),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_331),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_332),
.A2(n_273),
.B(n_300),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_254),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_279),
.B(n_254),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_291),
.A2(n_238),
.B(n_167),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_284),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_276),
.A2(n_236),
.B1(n_5),
.B2(n_6),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_285),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_346),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_347),
.A2(n_354),
.B(n_368),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_294),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_348),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_321),
.A2(n_292),
.B1(n_281),
.B2(n_299),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_350),
.A2(n_361),
.B1(n_365),
.B2(n_369),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_290),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_351),
.Y(n_387)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_353),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_313),
.A2(n_300),
.B(n_274),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_295),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_356),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_357),
.B(n_316),
.C(n_338),
.Y(n_394)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

INVx13_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_359),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_327),
.A2(n_342),
.B1(n_343),
.B2(n_322),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_362),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_367),
.Y(n_385)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_335),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_366),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_343),
.A2(n_322),
.B1(n_312),
.B2(n_310),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_334),
.Y(n_366)
);

OAI32xp33_ASAP7_75t_L g367 ( 
.A1(n_319),
.A2(n_282),
.A3(n_302),
.B1(n_304),
.B2(n_289),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_322),
.A2(n_280),
.B1(n_277),
.B2(n_270),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_311),
.B(n_286),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_371),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_296),
.Y(n_371)
);

AO22x1_ASAP7_75t_L g399 ( 
.A1(n_372),
.A2(n_324),
.B1(n_337),
.B2(n_340),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_341),
.B(n_296),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_375),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_322),
.A2(n_272),
.B1(n_271),
.B2(n_307),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_346),
.B(n_317),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_379),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_351),
.B(n_331),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_360),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_358),
.B(n_319),
.Y(n_382)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_382),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_328),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_395),
.C(n_349),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_330),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_387),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_333),
.Y(n_389)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_333),
.Y(n_391)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_391),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_344),
.A2(n_324),
.B1(n_323),
.B2(n_313),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_392),
.A2(n_375),
.B1(n_372),
.B2(n_355),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_394),
.B(n_360),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_338),
.C(n_318),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_399),
.A2(n_350),
.B1(n_369),
.B2(n_355),
.Y(n_412)
);

AO22x1_ASAP7_75t_L g401 ( 
.A1(n_372),
.A2(n_366),
.B1(n_367),
.B2(n_361),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_401),
.A2(n_372),
.B(n_272),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_345),
.B(n_326),
.Y(n_403)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_403),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_345),
.B(n_326),
.Y(n_404)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_404),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_309),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_405),
.B(n_374),
.Y(n_406)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_406),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_407),
.B(n_408),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_405),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_401),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_409),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_401),
.A2(n_344),
.B1(n_365),
.B2(n_352),
.Y(n_410)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_411),
.B(n_404),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_412),
.A2(n_392),
.B1(n_378),
.B2(n_399),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_383),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_421),
.Y(n_444)
);

NOR3xp33_ASAP7_75t_SL g415 ( 
.A(n_385),
.B(n_347),
.C(n_373),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_415),
.B(n_393),
.Y(n_449)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_416),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_347),
.C(n_368),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_420),
.C(n_427),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_353),
.C(n_373),
.Y(n_420)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_422),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_380),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_387),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_424),
.A2(n_399),
.B(n_388),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_372),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_429),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_330),
.C(n_339),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_386),
.B(n_309),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_433),
.A2(n_449),
.B1(n_413),
.B2(n_409),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_422),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_376),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_402),
.C(n_398),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_442),
.C(n_443),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_385),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_451),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_402),
.C(n_398),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_396),
.C(n_393),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g453 ( 
.A(n_445),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_378),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_450),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_448),
.A2(n_381),
.B(n_406),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_380),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_441),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_466),
.Y(n_482)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_438),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_457),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_446),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_465),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_447),
.B(n_430),
.Y(n_457)
);

INVx13_ASAP7_75t_L g458 ( 
.A(n_436),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_467),
.Y(n_468)
);

A2O1A1O1Ixp25_ASAP7_75t_L g459 ( 
.A1(n_439),
.A2(n_415),
.B(n_426),
.C(n_428),
.D(n_414),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_465),
.Y(n_472)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_463),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_376),
.Y(n_473)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_444),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_440),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_437),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_475),
.C(n_478),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_464),
.A2(n_443),
.B(n_431),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_471),
.A2(n_474),
.B(n_479),
.Y(n_484)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_472),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_473),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_464),
.A2(n_431),
.B(n_417),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_452),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_451),
.C(n_442),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_453),
.B(n_379),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_460),
.A2(n_419),
.B(n_396),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_377),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_467),
.B(n_377),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_481),
.B(n_469),
.C(n_476),
.Y(n_488)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_483),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_452),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_487),
.A2(n_397),
.B1(n_339),
.B2(n_359),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_488),
.A2(n_491),
.B(n_492),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_473),
.A2(n_433),
.B1(n_421),
.B2(n_390),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_490),
.A2(n_494),
.B1(n_382),
.B2(n_400),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_470),
.B(n_434),
.C(n_450),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_458),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_424),
.C(n_455),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_493),
.B(n_475),
.C(n_477),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_468),
.A2(n_412),
.B1(n_390),
.B2(n_459),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_499),
.C(n_320),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_498),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_484),
.A2(n_482),
.B(n_397),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_403),
.C(n_397),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_500),
.A2(n_501),
.B(n_320),
.Y(n_507)
);

OA21x2_ASAP7_75t_SL g501 ( 
.A1(n_485),
.A2(n_359),
.B(n_364),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_496),
.A2(n_489),
.B1(n_487),
.B2(n_492),
.Y(n_503)
);

NOR2x1_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_504),
.Y(n_510)
);

AOI322xp5_ASAP7_75t_L g504 ( 
.A1(n_499),
.A2(n_483),
.A3(n_493),
.B1(n_486),
.B2(n_320),
.C1(n_296),
.C2(n_275),
.Y(n_504)
);

OAI21xp33_ASAP7_75t_L g509 ( 
.A1(n_504),
.A2(n_506),
.B(n_303),
.Y(n_509)
);

O2A1O1Ixp33_ASAP7_75t_SL g508 ( 
.A1(n_507),
.A2(n_502),
.B(n_495),
.C(n_335),
.Y(n_508)
);

NAND4xp25_ASAP7_75t_L g511 ( 
.A(n_508),
.B(n_505),
.C(n_303),
.D(n_275),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_509),
.A2(n_510),
.B(n_275),
.Y(n_512)
);

AOI321xp33_ASAP7_75t_L g513 ( 
.A1(n_511),
.A2(n_512),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_513)
);

AOI322xp5_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_4),
.A3(n_5),
.B1(n_8),
.B2(n_9),
.C1(n_485),
.C2(n_435),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_514),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_4),
.B(n_8),
.C(n_9),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_9),
.Y(n_517)
);


endmodule