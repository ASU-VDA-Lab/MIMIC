module fake_jpeg_12417_n_523 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_523);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_523;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_50),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_51),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_9),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_52),
.B(n_67),
.Y(n_123)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_58),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_20),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g150 ( 
.A(n_61),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_16),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_98),
.Y(n_105)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_66),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_28),
.B(n_33),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_68),
.Y(n_132)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_28),
.B(n_9),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_76),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_29),
.B(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_84),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_94),
.Y(n_110)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_92),
.B(n_95),
.Y(n_128)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_96),
.B(n_97),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_37),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_106),
.B(n_89),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_48),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_107),
.B(n_143),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_56),
.A2(n_36),
.B1(n_37),
.B2(n_45),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_108),
.A2(n_111),
.B1(n_124),
.B2(n_155),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_65),
.A2(n_45),
.B1(n_26),
.B2(n_22),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_57),
.A2(n_26),
.B1(n_47),
.B2(n_42),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_112),
.A2(n_133),
.B1(n_141),
.B2(n_154),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_51),
.A2(n_26),
.B1(n_47),
.B2(n_42),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_114),
.A2(n_80),
.B(n_92),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_41),
.B1(n_47),
.B2(n_42),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_115),
.A2(n_121),
.B1(n_139),
.B2(n_147),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_54),
.A2(n_48),
.B1(n_29),
.B2(n_33),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_75),
.A2(n_45),
.B1(n_22),
.B2(n_47),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_38),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_129),
.B(n_135),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_58),
.A2(n_98),
.B1(n_97),
.B2(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_38),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_59),
.A2(n_41),
.B1(n_42),
.B2(n_22),
.Y(n_139)
);

AO22x2_ASAP7_75t_L g141 ( 
.A1(n_72),
.A2(n_44),
.B1(n_46),
.B2(n_43),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_35),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_73),
.A2(n_34),
.B1(n_43),
.B2(n_27),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_81),
.A2(n_34),
.B1(n_30),
.B2(n_44),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_84),
.A2(n_24),
.B1(n_30),
.B2(n_46),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_62),
.B(n_10),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_13),
.Y(n_192)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_150),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g270 ( 
.A(n_161),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_66),
.B(n_55),
.Y(n_162)
);

AOI32xp33_ASAP7_75t_L g246 ( 
.A1(n_162),
.A2(n_40),
.A3(n_10),
.B1(n_11),
.B2(n_16),
.Y(n_246)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_165),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_166),
.B(n_184),
.Y(n_254)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_170),
.Y(n_266)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_175),
.Y(n_227)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_180),
.Y(n_253)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_185),
.B(n_189),
.Y(n_257)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_186),
.B(n_187),
.Y(n_258)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_105),
.B(n_0),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_205),
.Y(n_236)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_191),
.B(n_193),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_192),
.B(n_194),
.Y(n_261)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_195),
.B(n_196),
.Y(n_268)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_101),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_108),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_197),
.Y(n_228)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_199),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_110),
.Y(n_200)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_201),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_239)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_203),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_146),
.A2(n_95),
.B1(n_91),
.B2(n_90),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_204),
.A2(n_46),
.B1(n_40),
.B2(n_2),
.Y(n_245)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_110),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_206),
.B(n_209),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_100),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_103),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.Y(n_241)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_141),
.B(n_132),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_146),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_125),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_131),
.A2(n_140),
.B1(n_119),
.B2(n_126),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_218),
.B(n_132),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_128),
.A2(n_46),
.B(n_9),
.C(n_12),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_145),
.A2(n_85),
.B1(n_87),
.B2(n_83),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_124),
.B1(n_111),
.B2(n_155),
.Y(n_223)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_221),
.B(n_264),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_223),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_114),
.B1(n_112),
.B2(n_141),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_238),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_141),
.B1(n_157),
.B2(n_102),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_167),
.A2(n_157),
.B1(n_102),
.B2(n_156),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_128),
.B1(n_160),
.B2(n_117),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_232),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_117),
.B1(n_160),
.B2(n_131),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_240),
.B(n_244),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_190),
.A2(n_140),
.B1(n_46),
.B2(n_40),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_245),
.B1(n_174),
.B2(n_188),
.Y(n_277)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_207),
.B1(n_166),
.B2(n_184),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_SL g308 ( 
.A(n_246),
.B(n_13),
.C(n_8),
.Y(n_308)
);

OA22x2_ASAP7_75t_L g251 ( 
.A1(n_191),
.A2(n_40),
.B1(n_1),
.B2(n_2),
.Y(n_251)
);

AO21x2_ASAP7_75t_L g293 ( 
.A1(n_251),
.A2(n_267),
.B(n_0),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_177),
.B(n_40),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_264),
.C(n_265),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_255),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_187),
.B(n_11),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_187),
.B(n_11),
.C(n_15),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g267 ( 
.A1(n_205),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_275),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_172),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_276),
.B(n_282),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_277),
.B(n_300),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_278),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_175),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_280),
.B(n_286),
.C(n_287),
.Y(n_350)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_261),
.B(n_161),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_240),
.A2(n_217),
.B(n_216),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_307),
.B(n_239),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_232),
.A2(n_181),
.B1(n_176),
.B2(n_164),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_284),
.A2(n_295),
.B1(n_310),
.B2(n_231),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_256),
.B(n_173),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_285),
.B(n_288),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_221),
.B(n_198),
.C(n_163),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_168),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_256),
.B(n_193),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_289),
.B(n_265),
.Y(n_320)
);

AOI32xp33_ASAP7_75t_L g290 ( 
.A1(n_228),
.A2(n_195),
.A3(n_208),
.B1(n_213),
.B2(n_183),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_290),
.A2(n_301),
.B(n_312),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_236),
.B(n_170),
.C(n_171),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_304),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_229),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_292),
.B(n_299),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_297),
.Y(n_321)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_244),
.A2(n_220),
.B1(n_201),
.B2(n_186),
.Y(n_295)
);

OAI32xp33_ASAP7_75t_L g296 ( 
.A1(n_257),
.A2(n_169),
.A3(n_212),
.B1(n_6),
.B2(n_7),
.Y(n_296)
);

XOR2x2_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_267),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_244),
.B(n_1),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_298),
.Y(n_342)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_263),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_254),
.A2(n_195),
.B(n_6),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_302),
.B(n_309),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_244),
.B(n_3),
.C(n_7),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_254),
.A2(n_3),
.B(n_8),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_315),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_268),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_254),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_317),
.B1(n_239),
.B2(n_241),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_SL g312 ( 
.A(n_258),
.B(n_269),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_222),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_313),
.B(n_248),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_258),
.B(n_3),
.C(n_14),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_272),
.Y(n_329)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_253),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_249),
.B(n_16),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_316),
.B(n_247),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_245),
.A2(n_228),
.B1(n_258),
.B2(n_249),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_318),
.A2(n_330),
.B(n_341),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_320),
.B(n_329),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_323),
.A2(n_348),
.B1(n_307),
.B2(n_278),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_281),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_331),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_271),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_336),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_306),
.A2(n_241),
.B(n_262),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_275),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_294),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_335),
.B(n_339),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_271),
.Y(n_336)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_298),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_267),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_345),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_297),
.A2(n_259),
.B(n_262),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_279),
.A2(n_253),
.B1(n_251),
.B2(n_234),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_343),
.A2(n_347),
.B1(n_351),
.B2(n_293),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_289),
.B(n_222),
.C(n_270),
.Y(n_344)
);

A2O1A1O1Ixp25_ASAP7_75t_L g383 ( 
.A1(n_344),
.A2(n_250),
.B(n_260),
.C(n_266),
.D(n_350),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_279),
.A2(n_251),
.B1(n_234),
.B2(n_267),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_295),
.A2(n_251),
.B1(n_248),
.B2(n_237),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_280),
.B(n_247),
.Y(n_352)
);

NAND3xp33_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_301),
.C(n_313),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_272),
.B(n_270),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_317),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_354),
.B(n_311),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_306),
.A2(n_230),
.B(n_233),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_356),
.A2(n_266),
.B(n_355),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_346),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_359),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_321),
.A2(n_274),
.B1(n_293),
.B2(n_304),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_360),
.A2(n_374),
.B1(n_375),
.B2(n_387),
.Y(n_409)
);

OAI32xp33_ASAP7_75t_L g361 ( 
.A1(n_321),
.A2(n_306),
.A3(n_336),
.B1(n_340),
.B2(n_327),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_361),
.B(n_362),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_345),
.Y(n_362)
);

AOI322xp5_ASAP7_75t_L g363 ( 
.A1(n_326),
.A2(n_274),
.A3(n_284),
.B1(n_296),
.B2(n_302),
.C1(n_283),
.C2(n_293),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_363),
.B(n_358),
.Y(n_414)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_377),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_349),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_379),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_319),
.C(n_329),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_347),
.A2(n_293),
.B1(n_277),
.B2(n_303),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_300),
.Y(n_376)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_376),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_335),
.B(n_314),
.Y(n_378)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_378),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_348),
.A2(n_303),
.B1(n_305),
.B2(n_308),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_328),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_382),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_348),
.A2(n_250),
.B1(n_260),
.B2(n_233),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_383),
.A2(n_385),
.B(n_388),
.Y(n_395)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_325),
.Y(n_384)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_384),
.Y(n_412)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_325),
.Y(n_386)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_351),
.A2(n_343),
.B1(n_337),
.B2(n_341),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_323),
.A2(n_355),
.B1(n_357),
.B2(n_322),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_334),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_391),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_318),
.A2(n_350),
.B1(n_332),
.B2(n_326),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_390),
.A2(n_342),
.B1(n_333),
.B2(n_357),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_338),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_334),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_392),
.B(n_324),
.Y(n_396)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_396),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_353),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_402),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_398),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_319),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_371),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_411),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_372),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_406),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_372),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_320),
.C(n_344),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_413),
.C(n_416),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_356),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_361),
.B(n_330),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_414),
.A2(n_422),
.B1(n_382),
.B2(n_380),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_359),
.B(n_354),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_415),
.B(n_417),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_358),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_381),
.B(n_322),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_376),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_366),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_370),
.B(n_358),
.C(n_342),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_420),
.B(n_365),
.C(n_367),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_424),
.B(n_435),
.Y(n_456)
);

XNOR2x1_ASAP7_75t_L g449 ( 
.A(n_425),
.B(n_439),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_378),
.C(n_365),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_437),
.C(n_440),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_391),
.Y(n_430)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_401),
.A2(n_369),
.B(n_385),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_431),
.A2(n_421),
.B(n_428),
.Y(n_461)
);

OAI22xp33_ASAP7_75t_L g432 ( 
.A1(n_409),
.A2(n_380),
.B1(n_362),
.B2(n_375),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_432),
.A2(n_446),
.B1(n_419),
.B2(n_412),
.Y(n_460)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_410),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_434),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_409),
.A2(n_379),
.B1(n_377),
.B2(n_366),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_420),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_402),
.B(n_383),
.C(n_387),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_416),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_438),
.B(n_445),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_404),
.B(n_383),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_360),
.C(n_384),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_393),
.B(n_389),
.C(n_392),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_443),
.C(n_444),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_393),
.B(n_386),
.C(n_333),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_374),
.C(n_363),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_405),
.B(n_406),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_407),
.B1(n_397),
.B2(n_399),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_430),
.A2(n_399),
.B(n_403),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_448),
.A2(n_449),
.B(n_466),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_413),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_450),
.B(n_463),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_444),
.A2(n_407),
.B1(n_395),
.B2(n_418),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_452),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_454),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_411),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_440),
.A2(n_395),
.B1(n_397),
.B2(n_394),
.Y(n_455)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_455),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_437),
.A2(n_419),
.B1(n_412),
.B2(n_421),
.Y(n_459)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_459),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_452),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_455),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_424),
.B(n_423),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_464),
.C(n_466),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_429),
.B(n_423),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_447),
.C(n_443),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_447),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_441),
.B(n_433),
.C(n_432),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_468),
.B(n_458),
.C(n_464),
.Y(n_475)
);

INVx11_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_469),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_448),
.A2(n_426),
.B1(n_442),
.B2(n_468),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_471),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_482),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_467),
.Y(n_476)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_476),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_453),
.C(n_451),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_477),
.B(n_478),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_462),
.C(n_456),
.Y(n_478)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_480),
.Y(n_495)
);

NOR2x1_ASAP7_75t_SL g489 ( 
.A(n_481),
.B(n_454),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_459),
.A2(n_449),
.B1(n_461),
.B2(n_465),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_484),
.B(n_450),
.Y(n_490)
);

XNOR2x1_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_490),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_480),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_491),
.B(n_492),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_469),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_484),
.B(n_463),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_493),
.B(n_496),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_482),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_478),
.A2(n_477),
.B(n_481),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_497),
.B(n_470),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_488),
.A2(n_483),
.B1(n_472),
.B2(n_479),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_501),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_488),
.A2(n_471),
.B1(n_472),
.B2(n_479),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_475),
.C(n_473),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_502),
.B(n_505),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_504),
.A2(n_470),
.B(n_489),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_495),
.A2(n_494),
.B1(n_485),
.B2(n_487),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_473),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_506),
.B(n_496),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_510),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_508),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_493),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_501),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_511),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_509),
.B(n_500),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_499),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_515),
.A2(n_512),
.B(n_499),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_517),
.A2(n_518),
.B(n_513),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_519),
.A2(n_514),
.B(n_516),
.Y(n_520)
);

NOR3xp33_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_503),
.C(n_490),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_521),
.B(n_503),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_474),
.Y(n_523)
);


endmodule