module fake_jpeg_6674_n_43 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_43);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_43;

wire n_33;
wire n_23;
wire n_27;
wire n_40;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_10),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_11),
.A2(n_1),
.B(n_21),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_33),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_14),
.B1(n_20),
.B2(n_3),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_2),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_34),
.A2(n_35),
.B1(n_27),
.B2(n_30),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_2),
.C(n_5),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_39),
.B(n_37),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_36),
.A3(n_38),
.B1(n_16),
.B2(n_17),
.C1(n_6),
.C2(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

NOR4xp25_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_7),
.C(n_18),
.D(n_22),
.Y(n_43)
);


endmodule