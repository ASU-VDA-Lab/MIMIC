module fake_jpeg_6623_n_95 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_95);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx6_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

AND2x4_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_27),
.Y(n_44)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_33),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_29),
.A2(n_22),
.B1(n_12),
.B2(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_13),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_37),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_26),
.B1(n_32),
.B2(n_31),
.Y(n_36)
);

OAI22x1_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_18),
.B1(n_2),
.B2(n_5),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_16),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_47),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_14),
.B(n_19),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_17),
.Y(n_59)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_16),
.Y(n_47)
);

AND2x6_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_22),
.Y(n_48)
);

AND2x6_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_21),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_12),
.B1(n_17),
.B2(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_18),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_26),
.B(n_1),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_19),
.B(n_17),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_48),
.B1(n_41),
.B2(n_36),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_12),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_51),
.C(n_45),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_61),
.B1(n_46),
.B2(n_37),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_50),
.B1(n_52),
.B2(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_66),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_77),
.Y(n_84)
);

AOI21x1_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_49),
.B(n_53),
.Y(n_72)
);

FAx1_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_61),
.CI(n_59),
.CON(n_81),
.SN(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_64),
.C(n_34),
.Y(n_82)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_35),
.C(n_45),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_65),
.C(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_82),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_74),
.C(n_69),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_40),
.C(n_38),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_73),
.B1(n_75),
.B2(n_67),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_72),
.B(n_77),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_87),
.B(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_78),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_91),
.A3(n_92),
.B1(n_89),
.B2(n_88),
.C1(n_85),
.C2(n_84),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_79),
.B(n_8),
.C(n_10),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_94),
.Y(n_95)
);


endmodule