module real_jpeg_29028_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_0),
.A2(n_26),
.B(n_129),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_1),
.A2(n_75),
.B1(n_76),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_1),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_1),
.A2(n_57),
.B1(n_59),
.B2(n_138),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_138),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_1),
.A2(n_28),
.B1(n_33),
.B2(n_138),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_59),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_3),
.A2(n_59),
.B(n_180),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_126),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_3),
.A2(n_10),
.B(n_28),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_3),
.B(n_60),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_3),
.A2(n_27),
.B1(n_100),
.B2(n_229),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_5),
.A2(n_75),
.B1(n_76),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_5),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_5),
.A2(n_57),
.B1(n_59),
.B2(n_112),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_112),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_5),
.A2(n_28),
.B1(n_33),
.B2(n_112),
.Y(n_221)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_7),
.A2(n_28),
.B1(n_33),
.B2(n_52),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_8),
.A2(n_28),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_8),
.A2(n_39),
.B1(n_75),
.B2(n_76),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_8),
.A2(n_39),
.B1(n_57),
.B2(n_59),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_8),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_9),
.A2(n_34),
.B1(n_57),
.B2(n_59),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_34),
.B1(n_43),
.B2(n_44),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_50),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_11),
.A2(n_28),
.B1(n_33),
.B2(n_50),
.Y(n_129)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_13),
.A2(n_57),
.B1(n_59),
.B2(n_64),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_14),
.A2(n_75),
.B1(n_76),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_14),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_14),
.A2(n_57),
.B1(n_59),
.B2(n_80),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_80),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_14),
.A2(n_28),
.B1(n_33),
.B2(n_80),
.Y(n_216)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_141),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_114),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_19),
.B(n_114),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_94),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_83),
.B2(n_84),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_24),
.B(n_40),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_35),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_27),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_27),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_27),
.A2(n_97),
.B1(n_100),
.B2(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_27),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_27),
.A2(n_35),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_27),
.A2(n_37),
.B1(n_221),
.B2(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_33),
.B1(n_46),
.B2(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_30),
.B(n_126),
.Y(n_233)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_32),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_33),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g87 ( 
.A(n_36),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_36),
.A2(n_178),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_38),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_38),
.A2(n_99),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_41),
.A2(n_51),
.B(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_41),
.A2(n_90),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_41),
.A2(n_47),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_41),
.A2(n_188),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_41),
.A2(n_47),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_41),
.A2(n_47),
.B1(n_187),
.B2(n_206),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_43),
.A2(n_57),
.A3(n_62),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_44),
.B(n_63),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_44),
.A2(n_46),
.B(n_126),
.C(n_208),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_47),
.A2(n_49),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_47),
.B(n_126),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_69),
.B2(n_70),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_65),
.Y(n_55)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_59),
.B1(n_73),
.B2(n_74),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_57),
.A2(n_77),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_59),
.B(n_73),
.Y(n_124)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_61),
.B(n_107),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_61),
.A2(n_67),
.B1(n_132),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_61),
.A2(n_67),
.B1(n_153),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_61),
.A2(n_67),
.B1(n_166),
.B2(n_184),
.Y(n_183)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_79),
.B(n_81),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_79),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_71),
.A2(n_111),
.B1(n_113),
.B2(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_72),
.A2(n_78),
.B1(n_125),
.B2(n_137),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B(n_77),
.C(n_78),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_75),
.Y(n_77)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g125 ( 
.A(n_75),
.B(n_126),
.CON(n_125),
.SN(n_125)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_93),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_92),
.B(n_150),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.C(n_109),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_101),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_101),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_109),
.B1(n_110),
.B2(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_108),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_131),
.B(n_133),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_113),
.B(n_126),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_120),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_115),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_120),
.A2(n_121),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_130),
.C(n_134),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_127),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_134),
.B1(n_135),
.B2(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_170),
.B(n_252),
.C(n_258),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_158),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_143),
.B(n_158),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_155),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_145),
.B(n_146),
.C(n_155),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_154),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_154),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_159),
.A2(n_160),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_164),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_168),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_193),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_167),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_251),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_244),
.B(n_250),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_199),
.B(n_243),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_189),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_174),
.B(n_189),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_182),
.C(n_185),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_175),
.A2(n_176),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_179),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_182),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_196),
.C(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_237),
.B(n_242),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_217),
.B(n_236),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_202),
.B(n_209),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_225),
.B(n_235),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_223),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_230),
.B(n_234),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_227),
.B(n_228),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_245),
.B(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);


endmodule