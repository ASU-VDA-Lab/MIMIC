module fake_jpeg_30626_n_222 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_56),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_58),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_26),
.C(n_21),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_55),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_34),
.B1(n_31),
.B2(n_49),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_33),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_36),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_35),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_32),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_38),
.A2(n_34),
.B1(n_20),
.B2(n_26),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_39),
.B1(n_44),
.B2(n_34),
.Y(n_94)
);

NOR2xp67_ASAP7_75t_SL g88 ( 
.A(n_42),
.B(n_32),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_80),
.B1(n_64),
.B2(n_53),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_80),
.B1(n_87),
.B2(n_85),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_69),
.Y(n_96)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_99),
.B(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_17),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_108),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_107),
.Y(n_120)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_100),
.B(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_17),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_76),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_87),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_69),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_61),
.A2(n_32),
.B1(n_18),
.B2(n_19),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_17),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_117),
.Y(n_135)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_30),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_23),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_130),
.B1(n_134),
.B2(n_106),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_114),
.B1(n_115),
.B2(n_92),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_79),
.B1(n_74),
.B2(n_66),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_108),
.B1(n_110),
.B2(n_117),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_32),
.B1(n_18),
.B2(n_66),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_106),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_94),
.A2(n_32),
.B1(n_18),
.B2(n_66),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_89),
.Y(n_149)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_153),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_151),
.B1(n_157),
.B2(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_150),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_121),
.B(n_78),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_149),
.B(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_103),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_101),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_97),
.Y(n_154)
);

NOR4xp25_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_158),
.C(n_159),
.D(n_23),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_90),
.B1(n_91),
.B2(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_156),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_129),
.A2(n_105),
.B1(n_74),
.B2(n_18),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_111),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_136),
.B(n_121),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_165),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_131),
.B(n_135),
.C(n_130),
.D(n_123),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_160),
.B(n_157),
.C(n_133),
.D(n_17),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_126),
.C(n_136),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_171),
.C(n_17),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_126),
.B(n_144),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_142),
.B1(n_147),
.B2(n_151),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_118),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_175),
.B(n_146),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_165),
.A2(n_143),
.B1(n_141),
.B2(n_150),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_181),
.B1(n_188),
.B2(n_173),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_178),
.A2(n_183),
.B1(n_186),
.B2(n_189),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_187),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_118),
.B1(n_133),
.B2(n_17),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_185),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_0),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_SL g190 ( 
.A1(n_180),
.A2(n_162),
.B(n_175),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_179),
.B(n_173),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_169),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_195),
.C(n_172),
.Y(n_205)
);

AOI321xp33_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_163),
.A3(n_164),
.B1(n_171),
.B2(n_170),
.C(n_161),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_161),
.B(n_167),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_161),
.C(n_167),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_182),
.C(n_183),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_203),
.C(n_204),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_191),
.C(n_197),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_201),
.B(n_202),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_189),
.C(n_186),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_195),
.C(n_193),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_16),
.C(n_14),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_211),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_14),
.B1(n_11),
.B2(n_10),
.Y(n_211)
);

AOI21x1_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_3),
.B(n_4),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_206),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_6),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_5),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_218),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_217),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_219),
.A2(n_213),
.B(n_212),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_220),
.Y(n_222)
);


endmodule