module real_jpeg_5892_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_313;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_1),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_1),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_1),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_1),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_1),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_1),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_1),
.B(n_261),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_1),
.B(n_367),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_2),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_2),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_2),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_2),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_2),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_2),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_2),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_2),
.B(n_294),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_3),
.Y(n_135)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_4),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_4),
.B(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_4),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_4),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_4),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_4),
.B(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_6),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_6),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_6),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_7),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_7),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_8),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_8),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_8),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_8),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_8),
.B(n_192),
.Y(n_191)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_10),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_10),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_10),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_11),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_11),
.B(n_79),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_11),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_12),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_12),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_12),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_12),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_12),
.B(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_13),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_14),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_14),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_14),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_14),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_14),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_15),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_15),
.B(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_15),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_15),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_15),
.B(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_208),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_207),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_168),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_19),
.B(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_19),
.B(n_211),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_19),
.B(n_211),
.Y(n_414)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_64),
.CI(n_126),
.CON(n_19),
.SN(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_53),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_34),
.B1(n_51),
.B2(n_52),
.Y(n_21)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_22),
.B(n_52),
.C(n_53),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.C(n_31),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_23),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_23),
.A2(n_31),
.B1(n_62),
.B2(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_23),
.B(n_55),
.C(n_59),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_23),
.A2(n_62),
.B1(n_274),
.B2(n_275),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_24),
.B(n_89),
.Y(n_88)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_24),
.B(n_105),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_24),
.B(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_26),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_28),
.Y(n_188)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_29),
.Y(n_148)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_31),
.B(n_179),
.C(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_31),
.A2(n_69),
.B1(n_178),
.B2(n_179),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_32),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g328 ( 
.A(n_33),
.Y(n_328)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_41),
.B2(n_50),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_35),
.A2(n_36),
.B1(n_146),
.B2(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_36),
.B(n_145),
.C(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_36),
.B(n_42),
.C(n_45),
.Y(n_183)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_40),
.Y(n_311)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_44),
.Y(n_277)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_48),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_48),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_48),
.Y(n_296)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_49),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_63),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_58),
.A2(n_59),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_58),
.A2(n_59),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_59),
.B(n_266),
.C(n_271),
.Y(n_351)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_62),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_96),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_65),
.B(n_97),
.C(n_115),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.C(n_86),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_66),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_71),
.B(n_86),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.C(n_82),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_72),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_77),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_82),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_78),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_78),
.Y(n_190)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_85),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_95),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_124),
.C(n_125),
.Y(n_123)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_93),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_115),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.C(n_112),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_99),
.B(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.C(n_107),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_100),
.A2(n_107),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_100),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_100),
.A2(n_240),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_104),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_104),
.Y(n_236)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_105),
.Y(n_268)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_107),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_112),
.Y(n_167)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_123),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_121),
.C(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_119),
.A2(n_122),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_149),
.C(n_166),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_127),
.B(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.C(n_144),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_128),
.B(n_144),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_130),
.B(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.C(n_140),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_131),
.B(n_140),
.Y(n_220)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_134),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_135),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_136),
.B(n_220),
.Y(n_219)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_139),
.Y(n_369)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_145),
.A2(n_382),
.B1(n_383),
.B2(n_385),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_145),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_146),
.Y(n_384)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_166),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.C(n_161),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_150),
.B(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_150),
.A2(n_151),
.B(n_153),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_157),
.B(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_158),
.B(n_161),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_162),
.B(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_162),
.B(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_162),
.B(n_318),
.Y(n_317)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_194),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_182),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_191),
.B2(n_193),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_188),
.Y(n_365)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_206),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_243),
.B(n_414),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.C(n_217),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_215),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_217),
.B(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_235),
.C(n_241),
.Y(n_217)
);

FAx1_ASAP7_75t_L g399 ( 
.A(n_218),
.B(n_235),
.CI(n_241),
.CON(n_399),
.SN(n_399)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.C(n_227),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_219),
.B(n_391),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_221),
.A2(n_227),
.B1(n_228),
.B2(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_221),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_222),
.B(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_229),
.A2(n_230),
.B1(n_233),
.B2(n_234),
.Y(n_352)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_232),
.Y(n_320)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_240),
.B(n_284),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_395),
.B(n_410),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_373),
.B(n_394),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_343),
.B(n_372),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_298),
.B(n_342),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_289),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_249),
.B(n_289),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_272),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_263),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_251),
.B(n_263),
.C(n_272),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.C(n_259),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_291)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_259),
.B(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_271),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_273),
.B(n_356),
.C(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_283),
.Y(n_278)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_279),
.Y(n_356)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_283),
.Y(n_357)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.C(n_297),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_290),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_292),
.A2(n_297),
.B1(n_334),
.B2(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_336),
.B(n_341),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_322),
.B(n_335),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_307),
.B(n_321),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_317),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_317),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_312),
.B(n_316),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_312),
.Y(n_316)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_324),
.B1(n_329),
.B2(n_330),
.Y(n_323)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx8_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_331),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_324),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_325),
.A2(n_326),
.B(n_329),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_333),
.B(n_334),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_337),
.B(n_338),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_345),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_353),
.B2(n_354),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_355),
.C(n_358),
.Y(n_374)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_348),
.B(n_351),
.C(n_352),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_361),
.B2(n_371),
.Y(n_358)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_359),
.Y(n_371)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_366),
.B2(n_370),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_370),
.C(n_371),
.Y(n_378)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_366),
.Y(n_370)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_375),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_388),
.B2(n_393),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_389),
.C(n_390),
.Y(n_404)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_381),
.C(n_386),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_381),
.B1(n_386),
.B2(n_387),
.Y(n_379)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_380),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_381),
.Y(n_387)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_383),
.Y(n_385)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_388),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_405),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_404),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_404),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_399),
.B(n_401),
.C(n_402),
.Y(n_406)
);

BUFx24_ASAP7_75t_SL g415 ( 
.A(n_399),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_405),
.A2(n_412),
.B(n_413),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_406),
.B(n_407),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);


endmodule