module real_jpeg_32931_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_0),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_0),
.Y(n_331)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_0),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_R g88 ( 
.A(n_1),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_1),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_1),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_1),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_1),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_2),
.B(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_2),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_2),
.A2(n_15),
.B1(n_201),
.B2(n_231),
.Y(n_230)
);

NAND2x1_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_3),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_3),
.B(n_29),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_3),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_3),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_3),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_4),
.B(n_212),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_4),
.Y(n_510)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_5),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_5),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_5),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_5),
.B(n_466),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_6),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_7),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_8),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_9),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_9),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_9),
.B(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_9),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_9),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_9),
.B(n_409),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_9),
.Y(n_435)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_10),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_11),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_12),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_12),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_12),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_12),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_12),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_12),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_12),
.B(n_191),
.Y(n_190)
);

NAND2x1_ASAP7_75t_L g274 ( 
.A(n_12),
.B(n_191),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_13),
.Y(n_203)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_14),
.Y(n_122)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_14),
.Y(n_242)
);

NAND2x1_ASAP7_75t_L g185 ( 
.A(n_15),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_15),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_15),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_15),
.B(n_367),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_15),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_15),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_15),
.B(n_482),
.Y(n_481)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_16),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_50),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_17),
.B(n_98),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_17),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_17),
.B(n_257),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_17),
.B(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_17),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_17),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_17),
.B(n_478),
.Y(n_477)
);

OAI211xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_213),
.B(n_509),
.C(n_511),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_210),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_20),
.B(n_211),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_208),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_152),
.Y(n_21)
);

NOR2xp67_ASAP7_75t_SL g209 ( 
.A(n_22),
.B(n_152),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_91),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_66),
.C(n_80),
.Y(n_23)
);

INVxp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_25),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.C(n_54),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_26),
.B(n_54),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_27),
.B(n_31),
.C(n_37),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_27),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_27),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_27),
.B(n_117),
.C(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_27),
.B(n_194),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_27),
.A2(n_118),
.B1(n_194),
.B2(n_195),
.Y(n_414)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_28),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_29),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_29),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_35),
.Y(n_178)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_39),
.Y(n_198)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_40),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_40),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_40),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_41),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_42),
.A2(n_43),
.B1(n_256),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_49),
.C(n_52),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_43),
.B(n_256),
.C(n_260),
.Y(n_255)
);

OR2x2_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_51),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_51),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_82),
.C(n_85),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_52),
.B(n_85),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_52),
.B(n_82),
.C(n_85),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_52),
.B(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_52),
.B(n_404),
.Y(n_440)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_53),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_62),
.Y(n_54)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_55),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_181)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_64),
.Y(n_494)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_67),
.A2(n_68),
.B1(n_80),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_69),
.B(n_71),
.C(n_77),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_75),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_76),
.A2(n_77),
.B1(n_86),
.B2(n_87),
.Y(n_207)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_81),
.C(n_86),
.Y(n_80)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_78),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_79),
.Y(n_298)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_82),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_82),
.A2(n_132),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_84),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_85),
.B(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_85),
.B(n_296),
.Y(n_380)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_138),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_125),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_111),
.C(n_112),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2x1_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_163),
.Y(n_162)
);

XOR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_101),
.C(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

NAND2x1_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_102),
.B(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_106),
.A2(n_107),
.B1(n_175),
.B2(n_176),
.Y(n_246)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_172),
.C(n_175),
.Y(n_171)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_124),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_119),
.B(n_290),
.C(n_294),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_119),
.A2(n_124),
.B1(n_294),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_122),
.Y(n_412)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_122),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

XOR2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_133),
.Y(n_126)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_148),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_140),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_140),
.A2(n_146),
.B1(n_252),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_146),
.B(n_248),
.C(n_252),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.C(n_164),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_154),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_313)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_165),
.B(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_182),
.C(n_204),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_166),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_179),
.Y(n_166)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_167),
.Y(n_302)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_170),
.A2(n_171),
.B1(n_179),
.B2(n_180),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_172),
.B(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_182),
.A2(n_183),
.B1(n_204),
.B2(n_205),
.Y(n_268)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_197),
.C(n_199),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_226),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.C(n_194),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_185),
.A2(n_194),
.B1(n_195),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_185),
.Y(n_277)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_193),
.Y(n_370)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_193),
.Y(n_428)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_196),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_197),
.A2(n_199),
.B1(n_200),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_198),
.Y(n_373)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_210),
.B(n_510),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_215),
.Y(n_513)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_388),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_314),
.B(n_384),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g388 ( 
.A(n_218),
.B(n_389),
.C(n_507),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_269),
.B1(n_308),
.B2(n_311),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_220),
.B(n_270),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_264),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_222),
.B(n_267),
.C(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.C(n_243),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_229),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.C(n_236),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_230),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_235),
.B(n_237),
.Y(n_282)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_242),
.Y(n_464)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_244),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.C(n_255),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_245),
.B(n_255),
.Y(n_351)
);

XOR2x2_ASAP7_75t_L g350 ( 
.A(n_247),
.B(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_287),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_251),
.Y(n_407)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

INVx3_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_256),
.Y(n_340)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_260),
.B(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

INVx3_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_263),
.B(n_488),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_263),
.B(n_493),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_265),
.Y(n_310)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_300),
.C(n_304),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_318),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_284),
.B(n_299),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_279),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_279),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_273),
.B(n_280),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_278),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OA21x2_ASAP7_75t_SL g341 ( 
.A1(n_281),
.A2(n_342),
.B(n_345),
.Y(n_341)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_282),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_284),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_289),
.C(n_295),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_286),
.B(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_289),
.B(n_295),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_290),
.B(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_292),
.Y(n_466)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_294),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_301),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_319),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_309),
.B(n_312),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_309),
.B(n_312),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_352),
.B(n_383),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_316),
.B(n_508),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_317),
.B(n_320),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.C(n_350),
.Y(n_320)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_321),
.Y(n_356)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_338),
.C(n_341),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.C(n_332),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_325),
.A2(n_326),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_327),
.A2(n_328),
.B1(n_332),
.B2(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_330),
.B(n_422),
.Y(n_486)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx12f_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_341),
.Y(n_359)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_350),
.B(n_355),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_357),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_353),
.B(n_357),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.C(n_381),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_381),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.C(n_379),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_361),
.B(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_364),
.A2(n_379),
.B1(n_380),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_364),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_371),
.C(n_374),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_365),
.A2(n_366),
.B1(n_374),
.B2(n_375),
.Y(n_448)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_371),
.B(n_448),
.Y(n_447)
);

INVx3_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_386),
.B(n_387),
.Y(n_384)
);

AO21x1_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_415),
.B(n_506),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_393),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_391),
.B(n_393),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_398),
.C(n_401),
.Y(n_393)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_395),
.B(n_504),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_398),
.B(n_401),
.Y(n_504)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_408),
.C(n_413),
.Y(n_401)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_402),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_406),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_408),
.A2(n_413),
.B1(n_414),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_416),
.A2(n_500),
.B(n_505),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_455),
.B(n_499),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_441),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g499 ( 
.A(n_418),
.B(n_441),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_432),
.C(n_440),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_419),
.B(n_468),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_429),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_425),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_429),
.C(n_445),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_432),
.A2(n_433),
.B1(n_440),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_434),
.A2(n_437),
.B1(n_438),
.B2(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_434),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_440),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_449),
.B1(n_453),
.B2(n_454),
.Y(n_441)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_442),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_444),
.B1(n_446),
.B2(n_447),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_444),
.B(n_454),
.C(n_502),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_446),
.Y(n_502)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_449),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_470),
.B(n_498),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_467),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_457),
.B(n_467),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_461),
.C(n_465),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_458),
.A2(n_459),
.B1(n_473),
.B2(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_461),
.B(n_465),
.Y(n_474)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_484),
.B(n_497),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_475),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_475),
.Y(n_497)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_480),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_476),
.A2(n_477),
.B1(n_480),
.B2(n_481),
.Y(n_495)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_491),
.B(n_496),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.Y(n_485)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_495),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_492),
.B(n_495),
.Y(n_496)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_503),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_501),
.B(n_503),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_512),
.B(n_513),
.Y(n_511)
);


endmodule