module fake_jpeg_6610_n_308 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_308);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_33),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_22),
.B(n_19),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_22),
.B1(n_19),
.B2(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_48),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_29),
.A2(n_33),
.B(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_59),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_38),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_70),
.Y(n_76)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_38),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_46),
.Y(n_79)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_47),
.B(n_22),
.C(n_32),
.D(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_79),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp67_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_45),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_24),
.B1(n_14),
.B2(n_18),
.Y(n_111)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_53),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_43),
.B1(n_54),
.B2(n_24),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_88),
.B1(n_66),
.B2(n_64),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_95),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_43),
.B1(n_31),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_43),
.B1(n_31),
.B2(n_14),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_63),
.B1(n_64),
.B2(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_23),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_23),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_17),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_74),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_36),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_106),
.B1(n_85),
.B2(n_57),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_102),
.Y(n_130)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_66),
.B1(n_56),
.B2(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_111),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_61),
.C(n_56),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_18),
.C(n_17),
.Y(n_142)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_113),
.Y(n_120)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_72),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_89),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_57),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_118),
.Y(n_144)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

OAI22x1_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_76),
.B1(n_77),
.B2(n_87),
.Y(n_121)
);

OAI22x1_ASAP7_75t_SL g154 ( 
.A1(n_121),
.A2(n_105),
.B1(n_99),
.B2(n_103),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_87),
.B(n_78),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_129),
.B(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_133),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_89),
.B(n_13),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_79),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_104),
.Y(n_153)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_101),
.A2(n_97),
.B(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_102),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_116),
.C(n_113),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_134),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

CKINVDCx10_ASAP7_75t_R g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_155),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_SL g184 ( 
.A1(n_154),
.A2(n_34),
.B(n_37),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_161),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_162),
.Y(n_194)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_121),
.A2(n_114),
.B1(n_103),
.B2(n_24),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_166),
.B(n_171),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_37),
.C(n_34),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_133),
.C(n_127),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_122),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_102),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_157),
.A2(n_139),
.B1(n_143),
.B2(n_131),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_172),
.A2(n_188),
.B1(n_67),
.B2(n_71),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_168),
.Y(n_202)
);

AOI321xp33_ASAP7_75t_SL g177 ( 
.A1(n_154),
.A2(n_170),
.A3(n_153),
.B1(n_167),
.B2(n_156),
.C(n_151),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_161),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_189),
.C(n_193),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_192),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_150),
.B1(n_169),
.B2(n_149),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_146),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_13),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_151),
.A2(n_135),
.B1(n_114),
.B2(n_128),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_147),
.C(n_148),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_144),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_128),
.C(n_141),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_109),
.Y(n_196)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_145),
.B(n_158),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_202),
.Y(n_230)
);

XNOR2x2_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_160),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_207),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_187),
.A2(n_141),
.B(n_34),
.C(n_37),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_200),
.A2(n_218),
.B1(n_178),
.B2(n_173),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_175),
.B(n_166),
.Y(n_204)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_185),
.B(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_168),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_212),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_168),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_209),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_36),
.C(n_141),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_179),
.B(n_94),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_58),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_36),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_23),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_169),
.B1(n_94),
.B2(n_13),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_235),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_191),
.C(n_183),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_225),
.C(n_233),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_208),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_200),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_181),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_234),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_191),
.C(n_174),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_180),
.B1(n_194),
.B2(n_188),
.Y(n_229)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_207),
.A2(n_173),
.B1(n_190),
.B2(n_27),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_190),
.C(n_58),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_201),
.A2(n_27),
.B1(n_18),
.B2(n_17),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

BUFx12_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_211),
.A2(n_27),
.B1(n_53),
.B2(n_20),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_200),
.B(n_8),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_242),
.A2(n_11),
.B(n_9),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_21),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_200),
.B(n_36),
.Y(n_247)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_16),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_251),
.C(n_252),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_69),
.B(n_11),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_0),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_16),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_227),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_11),
.C(n_9),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_255),
.C(n_0),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_16),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_219),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_256),
.A2(n_258),
.B(n_265),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_226),
.B1(n_236),
.B2(n_221),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_269),
.B1(n_246),
.B2(n_251),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_237),
.B(n_234),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_2),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_248),
.C(n_240),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_20),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_268),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_1),
.Y(n_269)
);

NAND2xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_254),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_277),
.B(n_259),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_240),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_280),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_3),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_269),
.C(n_266),
.Y(n_283)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_275),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_3),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_270),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_290),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_276),
.B(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_291),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_3),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_3),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_288),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_SL g301 ( 
.A1(n_293),
.A2(n_296),
.B(n_290),
.C(n_297),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_298),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_287),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g303 ( 
.A1(n_299),
.A2(n_301),
.A3(n_284),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_4),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_293),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.C(n_7),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_5),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_305),
.A2(n_5),
.B(n_6),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_306),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_307),
.B(n_6),
.CI(n_7),
.CON(n_308),
.SN(n_308)
);


endmodule