module fake_ariane_1328_n_105 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_4, n_10, n_105);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_4;
input n_10;

output n_105;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_18;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_17;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVxp67_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVxp33_ASAP7_75t_SL g28 ( 
.A(n_14),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

AND2x4_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_23),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

AND2x4_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_30),
.B1(n_20),
.B2(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_28),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_17),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_42),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_R g57 ( 
.A(n_48),
.B(n_37),
.Y(n_57)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_42),
.B1(n_37),
.B2(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_52),
.Y(n_59)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

OAI211xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_49),
.B(n_55),
.C(n_47),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_54),
.Y(n_66)
);

AOI222xp33_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_45),
.B1(n_33),
.B2(n_31),
.C1(n_38),
.C2(n_58),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_54),
.B1(n_52),
.B2(n_56),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

OAI221xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_67),
.B1(n_55),
.B2(n_65),
.C(n_44),
.Y(n_74)
);

OAI332xp33_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_39),
.A3(n_40),
.B1(n_51),
.B2(n_19),
.B3(n_53),
.C1(n_43),
.C2(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

OAI33xp33_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_46),
.A3(n_53),
.B1(n_63),
.B2(n_62),
.B3(n_69),
.Y(n_78)
);

AOI221xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_58),
.B1(n_36),
.B2(n_48),
.C(n_70),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_70),
.Y(n_80)
);

NAND2x1p5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_1),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_81),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_79),
.B1(n_72),
.B2(n_68),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_56),
.C(n_72),
.Y(n_89)
);

AND2x4_ASAP7_75t_SL g90 ( 
.A(n_87),
.B(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_86),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_89),
.B(n_85),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_61),
.C(n_52),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_54),
.B(n_56),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_92),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_3),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_93),
.B1(n_56),
.B2(n_5),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_98)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_96),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

XNOR2x1_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_7),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_99),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_100),
.A3(n_9),
.B1(n_10),
.B2(n_8),
.C1(n_13),
.C2(n_15),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_103),
.B(n_10),
.Y(n_105)
);


endmodule