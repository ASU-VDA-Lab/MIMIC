module real_aes_1259_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_626;
wire n_400;
wire n_539;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_755;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_0), .B(n_130), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_1), .A2(n_139), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_2), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_3), .B(n_146), .Y(n_209) );
INVx1_ASAP7_75t_L g137 ( .A(n_4), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_5), .B(n_146), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_6), .B(n_150), .Y(n_478) );
INVx1_ASAP7_75t_L g512 ( .A(n_7), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g812 ( .A1(n_8), .A2(n_813), .B1(n_816), .B2(n_817), .Y(n_812) );
INVx1_ASAP7_75t_L g816 ( .A(n_8), .Y(n_816) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_9), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_10), .Y(n_550) );
NAND2xp33_ASAP7_75t_L g147 ( .A(n_11), .B(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g127 ( .A(n_12), .Y(n_127) );
AOI221x1_ASAP7_75t_L g225 ( .A1(n_13), .A2(n_25), .B1(n_130), .B2(n_139), .C(n_226), .Y(n_225) );
AND3x1_ASAP7_75t_L g110 ( .A(n_14), .B(n_38), .C(n_111), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_14), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g129 ( .A(n_15), .B(n_130), .Y(n_129) );
AO21x2_ASAP7_75t_L g124 ( .A1(n_16), .A2(n_125), .B(n_128), .Y(n_124) );
INVx1_ASAP7_75t_L g487 ( .A(n_17), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_18), .B(n_164), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_19), .B(n_146), .Y(n_173) );
AO21x1_ASAP7_75t_L g204 ( .A1(n_20), .A2(n_130), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g109 ( .A(n_21), .Y(n_109) );
INVx1_ASAP7_75t_L g485 ( .A(n_22), .Y(n_485) );
INVx1_ASAP7_75t_SL g495 ( .A(n_23), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_24), .B(n_131), .Y(n_578) );
NAND2x1_ASAP7_75t_L g195 ( .A(n_26), .B(n_146), .Y(n_195) );
AOI33xp33_ASAP7_75t_L g524 ( .A1(n_27), .A2(n_55), .A3(n_462), .B1(n_467), .B2(n_525), .B3(n_526), .Y(n_524) );
NAND2x1_ASAP7_75t_L g183 ( .A(n_28), .B(n_148), .Y(n_183) );
INVx1_ASAP7_75t_L g544 ( .A(n_29), .Y(n_544) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_30), .A2(n_89), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g151 ( .A(n_30), .B(n_89), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_31), .B(n_470), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_32), .B(n_148), .Y(n_163) );
INVxp33_ASAP7_75t_L g822 ( .A(n_33), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_34), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_35), .B(n_148), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_36), .A2(n_139), .B(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g136 ( .A(n_37), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g140 ( .A(n_37), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g461 ( .A(n_37), .Y(n_461) );
OR2x6_ASAP7_75t_L g445 ( .A(n_38), .B(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_39), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_40), .B(n_130), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_41), .B(n_470), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_42), .A2(n_150), .B1(n_157), .B2(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_43), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_44), .B(n_131), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_45), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_46), .B(n_148), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_47), .A2(n_785), .B1(n_786), .B2(n_787), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_47), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_48), .B(n_125), .Y(n_514) );
XNOR2xp5_ASAP7_75t_SL g808 ( .A(n_48), .B(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_49), .B(n_131), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_50), .A2(n_139), .B(n_182), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_51), .Y(n_575) );
XOR2xp5_ASAP7_75t_L g787 ( .A(n_52), .B(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_53), .B(n_148), .Y(n_196) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_54), .A2(n_784), .B1(n_792), .B2(n_794), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_56), .B(n_131), .Y(n_536) );
INVx1_ASAP7_75t_L g133 ( .A(n_57), .Y(n_133) );
INVx1_ASAP7_75t_L g143 ( .A(n_57), .Y(n_143) );
AND2x2_ASAP7_75t_L g537 ( .A(n_58), .B(n_164), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_59), .A2(n_76), .B1(n_459), .B2(n_470), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_60), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_61), .B(n_146), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_62), .B(n_157), .Y(n_552) );
AOI21xp5_ASAP7_75t_SL g458 ( .A1(n_63), .A2(n_459), .B(n_464), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_64), .A2(n_139), .B(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g481 ( .A(n_65), .Y(n_481) );
AO21x1_ASAP7_75t_L g206 ( .A1(n_66), .A2(n_139), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_67), .B(n_130), .Y(n_159) );
INVx1_ASAP7_75t_L g535 ( .A(n_68), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_69), .B(n_130), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_70), .A2(n_459), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g219 ( .A(n_71), .B(n_165), .Y(n_219) );
INVx1_ASAP7_75t_L g135 ( .A(n_72), .Y(n_135) );
INVx1_ASAP7_75t_L g141 ( .A(n_72), .Y(n_141) );
AND2x2_ASAP7_75t_L g187 ( .A(n_73), .B(n_156), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_74), .B(n_470), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_75), .B(n_804), .Y(n_803) );
OAI22xp5_ASAP7_75t_SL g813 ( .A1(n_77), .A2(n_87), .B1(n_814), .B2(n_815), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_77), .Y(n_814) );
AND2x2_ASAP7_75t_L g497 ( .A(n_78), .B(n_156), .Y(n_497) );
INVx1_ASAP7_75t_L g482 ( .A(n_79), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_80), .A2(n_459), .B(n_494), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g576 ( .A1(n_81), .A2(n_459), .B(n_519), .C(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_82), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g447 ( .A(n_82), .Y(n_447) );
AND2x2_ASAP7_75t_L g155 ( .A(n_83), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_84), .B(n_130), .Y(n_175) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_85), .B(n_156), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_86), .A2(n_459), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g815 ( .A(n_87), .Y(n_815) );
AND2x2_ASAP7_75t_L g205 ( .A(n_88), .B(n_150), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_90), .B(n_148), .Y(n_174) );
AND2x2_ASAP7_75t_L g199 ( .A(n_91), .B(n_156), .Y(n_199) );
INVx1_ASAP7_75t_L g465 ( .A(n_92), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_93), .B(n_146), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_94), .A2(n_139), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_95), .B(n_148), .Y(n_227) );
AND2x2_ASAP7_75t_L g528 ( .A(n_96), .B(n_156), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_97), .A2(n_98), .B1(n_789), .B2(n_790), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_97), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_98), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_99), .B(n_146), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_100), .A2(n_542), .B(n_543), .C(n_545), .Y(n_541) );
BUFx2_ASAP7_75t_L g802 ( .A(n_101), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_102), .A2(n_139), .B(n_144), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_103), .B(n_131), .Y(n_468) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_114), .B(n_821), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_SL g823 ( .A(n_106), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_110), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_109), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OA22x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_798), .B1(n_802), .B2(n_807), .Y(n_114) );
OAI21xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_784), .B(n_791), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_440), .B1(n_448), .B2(n_782), .Y(n_117) );
INVx2_ASAP7_75t_L g793 ( .A(n_118), .Y(n_793) );
OAI22x1_ASAP7_75t_SL g809 ( .A1(n_118), .A2(n_810), .B1(n_811), .B2(n_812), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_118), .Y(n_810) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_361), .Y(n_118) );
NOR3xp33_ASAP7_75t_SL g119 ( .A(n_120), .B(n_273), .C(n_313), .Y(n_119) );
OAI221xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_188), .B1(n_237), .B2(n_252), .C(n_255), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_152), .Y(n_122) );
INVx2_ASAP7_75t_L g270 ( .A(n_123), .Y(n_270) );
AND2x2_ASAP7_75t_L g300 ( .A(n_123), .B(n_301), .Y(n_300) );
BUFx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g238 ( .A(n_124), .B(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g245 ( .A(n_124), .B(n_178), .Y(n_245) );
INVx2_ASAP7_75t_L g251 ( .A(n_124), .Y(n_251) );
AND2x2_ASAP7_75t_L g260 ( .A(n_124), .B(n_154), .Y(n_260) );
INVx1_ASAP7_75t_L g276 ( .A(n_124), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_124), .B(n_322), .Y(n_321) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_125), .A2(n_510), .B(n_514), .Y(n_509) );
INVx2_ASAP7_75t_SL g519 ( .A(n_125), .Y(n_519) );
BUFx4f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx3_ASAP7_75t_L g157 ( .A(n_126), .Y(n_157) );
AND2x4_ASAP7_75t_L g150 ( .A(n_127), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_127), .B(n_151), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_138), .B(n_150), .Y(n_128) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_136), .Y(n_130) );
INVx1_ASAP7_75t_L g483 ( .A(n_131), .Y(n_483) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
AND2x6_ASAP7_75t_L g148 ( .A(n_132), .B(n_141), .Y(n_148) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g146 ( .A(n_134), .B(n_143), .Y(n_146) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx5_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_136), .Y(n_545) );
AND2x2_ASAP7_75t_L g142 ( .A(n_137), .B(n_143), .Y(n_142) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_137), .Y(n_472) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
BUFx3_ASAP7_75t_L g473 ( .A(n_140), .Y(n_473) );
INVx2_ASAP7_75t_L g463 ( .A(n_141), .Y(n_463) );
AND2x4_ASAP7_75t_L g459 ( .A(n_142), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g467 ( .A(n_143), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_147), .B(n_149), .Y(n_144) );
INVxp67_ASAP7_75t_L g488 ( .A(n_146), .Y(n_488) );
INVxp67_ASAP7_75t_L g486 ( .A(n_148), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_149), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_149), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_149), .A2(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_149), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_149), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_149), .A2(n_216), .B(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_149), .A2(n_227), .B(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_149), .A2(n_465), .B(n_466), .C(n_468), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_149), .B(n_150), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g494 ( .A1(n_149), .A2(n_466), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_149), .A2(n_466), .B(n_512), .C(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g522 ( .A(n_149), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_149), .A2(n_466), .B(n_535), .C(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_149), .A2(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_SL g169 ( .A(n_150), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_150), .B(n_211), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_150), .A2(n_458), .B(n_469), .Y(n_457) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_166), .Y(n_152) );
INVx4_ASAP7_75t_L g241 ( .A(n_153), .Y(n_241) );
AND2x2_ASAP7_75t_L g272 ( .A(n_153), .B(n_179), .Y(n_272) );
AND2x2_ASAP7_75t_L g348 ( .A(n_153), .B(n_322), .Y(n_348) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_153), .B(n_178), .Y(n_390) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_154), .B(n_178), .Y(n_277) );
AND2x2_ASAP7_75t_L g301 ( .A(n_154), .B(n_179), .Y(n_301) );
BUFx2_ASAP7_75t_L g317 ( .A(n_154), .Y(n_317) );
NOR2x1_ASAP7_75t_SL g420 ( .A(n_154), .B(n_322), .Y(n_420) );
OR2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_158), .Y(n_154) );
INVx3_ASAP7_75t_L g198 ( .A(n_156), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_156), .A2(n_198), .B1(n_541), .B2(n_546), .Y(n_540) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_157), .B(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_164), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_164), .Y(n_186) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_164), .A2(n_225), .B(n_229), .Y(n_224) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_164), .A2(n_225), .B(n_229), .Y(n_287) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g297 ( .A(n_166), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_166), .A2(n_364), .B1(n_366), .B2(n_368), .C(n_373), .Y(n_363) );
AND2x2_ASAP7_75t_L g383 ( .A(n_166), .B(n_276), .Y(n_383) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_178), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g239 ( .A(n_168), .Y(n_239) );
INVx1_ASAP7_75t_L g292 ( .A(n_168), .Y(n_292) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_176), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_169), .B(n_177), .Y(n_176) );
AO21x2_ASAP7_75t_L g322 ( .A1(n_169), .A2(n_170), .B(n_176), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_175), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_178), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g261 ( .A(n_178), .B(n_249), .Y(n_261) );
INVx2_ASAP7_75t_L g303 ( .A(n_178), .Y(n_303) );
AND2x2_ASAP7_75t_L g436 ( .A(n_178), .B(n_251), .Y(n_436) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_179), .Y(n_293) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_186), .B(n_187), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_185), .Y(n_180) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_186), .A2(n_491), .B(n_497), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_220), .C(n_235), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_200), .Y(n_189) );
INVx2_ASAP7_75t_L g350 ( .A(n_190), .Y(n_350) );
AND2x2_ASAP7_75t_L g395 ( .A(n_190), .B(n_272), .Y(n_395) );
BUFx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g340 ( .A(n_191), .Y(n_340) );
AND2x4_ASAP7_75t_SL g355 ( .A(n_191), .B(n_267), .Y(n_355) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_198), .B(n_199), .Y(n_191) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_192), .A2(n_198), .B(n_199), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_197), .Y(n_192) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_198), .A2(n_213), .B(n_219), .Y(n_212) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_198), .A2(n_213), .B(n_219), .Y(n_232) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_198), .A2(n_531), .B(n_537), .Y(n_530) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_198), .A2(n_531), .B(n_537), .Y(n_560) );
INVx2_ASAP7_75t_L g309 ( .A(n_200), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_200), .B(n_339), .Y(n_365) );
AND2x4_ASAP7_75t_L g398 ( .A(n_200), .B(n_345), .Y(n_398) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_212), .Y(n_200) );
AND2x2_ASAP7_75t_L g236 ( .A(n_201), .B(n_231), .Y(n_236) );
OR2x2_ASAP7_75t_L g266 ( .A(n_201), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_SL g335 ( .A(n_201), .B(n_287), .Y(n_335) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx2_ASAP7_75t_L g280 ( .A(n_202), .Y(n_280) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g254 ( .A(n_203), .Y(n_254) );
OAI21x1_ASAP7_75t_SL g203 ( .A1(n_204), .A2(n_206), .B(n_210), .Y(n_203) );
INVx1_ASAP7_75t_L g211 ( .A(n_205), .Y(n_211) );
INVx2_ASAP7_75t_L g267 ( .A(n_212), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_214), .B(n_218), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_220), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_230), .Y(n_221) );
AND2x2_ASAP7_75t_L g235 ( .A(n_222), .B(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g308 ( .A(n_222), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g393 ( .A(n_222), .Y(n_393) );
BUFx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g253 ( .A(n_223), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g372 ( .A(n_223), .B(n_232), .Y(n_372) );
AND2x2_ASAP7_75t_L g376 ( .A(n_223), .B(n_242), .Y(n_376) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g345 ( .A(n_224), .Y(n_345) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_224), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_230), .B(n_253), .Y(n_329) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_231), .B(n_254), .Y(n_439) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g243 ( .A(n_232), .B(n_234), .Y(n_243) );
AND2x2_ASAP7_75t_L g325 ( .A(n_232), .B(n_287), .Y(n_325) );
AND2x2_ASAP7_75t_L g344 ( .A(n_232), .B(n_233), .Y(n_344) );
BUFx2_ASAP7_75t_L g265 ( .A(n_233), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_233), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
BUFx3_ASAP7_75t_L g242 ( .A(n_234), .Y(n_242) );
INVxp67_ASAP7_75t_L g285 ( .A(n_234), .Y(n_285) );
INVx1_ASAP7_75t_L g258 ( .A(n_236), .Y(n_258) );
AND2x2_ASAP7_75t_L g294 ( .A(n_236), .B(n_265), .Y(n_294) );
NAND2xp33_ASAP7_75t_L g375 ( .A(n_236), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g412 ( .A(n_236), .B(n_413), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_240), .B1(n_243), .B2(n_244), .C(n_246), .Y(n_237) );
AND2x2_ASAP7_75t_L g341 ( .A(n_238), .B(n_241), .Y(n_341) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_238), .B(n_301), .Y(n_360) );
AND2x2_ASAP7_75t_L g378 ( .A(n_238), .B(n_303), .Y(n_378) );
AND2x2_ASAP7_75t_L g433 ( .A(n_238), .B(n_272), .Y(n_433) );
INVx1_ASAP7_75t_L g249 ( .A(n_239), .Y(n_249) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_239), .Y(n_305) );
CKINVDCx16_ASAP7_75t_R g385 ( .A(n_240), .Y(n_385) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_241), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_241), .B(n_292), .Y(n_367) );
AND2x2_ASAP7_75t_L g334 ( .A(n_242), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g370 ( .A(n_242), .Y(n_370) );
AND2x2_ASAP7_75t_L g279 ( .A(n_243), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_243), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g421 ( .A(n_243), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_243), .B(n_345), .Y(n_431) );
AND2x4_ASAP7_75t_L g347 ( .A(n_244), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g418 ( .A(n_245), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
OR2x2_ASAP7_75t_L g289 ( .A(n_250), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g296 ( .A(n_251), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g327 ( .A(n_251), .B(n_301), .Y(n_327) );
AND2x2_ASAP7_75t_L g401 ( .A(n_251), .B(n_322), .Y(n_401) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g349 ( .A(n_253), .B(n_350), .Y(n_349) );
OAI32xp33_ASAP7_75t_L g414 ( .A1(n_253), .A2(n_415), .A3(n_417), .B1(n_418), .B2(n_421), .Y(n_414) );
AND2x4_ASAP7_75t_L g286 ( .A(n_254), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g384 ( .A(n_254), .B(n_287), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_259), .B1(n_262), .B2(n_268), .Y(n_255) );
INVxp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g373 ( .A1(n_257), .A2(n_271), .B(n_374), .C(n_375), .Y(n_373) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g357 ( .A(n_258), .B(n_285), .Y(n_357) );
INVx1_ASAP7_75t_SL g428 ( .A(n_259), .Y(n_428) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x4_ASAP7_75t_L g331 ( .A(n_261), .B(n_270), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_261), .A2(n_410), .B1(n_411), .B2(n_412), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_266), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_269), .A2(n_299), .B1(n_352), .B2(n_353), .Y(n_351) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
OAI211xp5_ASAP7_75t_SL g387 ( .A1(n_270), .A2(n_388), .B(n_396), .C(n_409), .Y(n_387) );
INVx2_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g307 ( .A(n_272), .B(n_276), .Y(n_307) );
OAI211xp5_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_278), .B(n_281), .C(n_310), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g304 ( .A(n_276), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g424 ( .A(n_276), .B(n_420), .Y(n_424) );
OAI32xp33_ASAP7_75t_L g381 ( .A1(n_277), .A2(n_382), .A3(n_384), .B1(n_385), .B2(n_386), .Y(n_381) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_280), .B(n_372), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_288), .B1(n_294), .B2(n_295), .C(n_298), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g438 ( .A(n_285), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_286), .B(n_350), .Y(n_352) );
A2O1A1O1Ixp25_ASAP7_75t_L g423 ( .A1(n_286), .A2(n_355), .B(n_371), .C(n_417), .D(n_424), .Y(n_423) );
AOI31xp33_ASAP7_75t_L g425 ( .A1(n_286), .A2(n_307), .A3(n_417), .B(n_424), .Y(n_425) );
AND2x2_ASAP7_75t_L g339 ( .A(n_287), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_289), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx2_ASAP7_75t_L g416 ( .A(n_291), .Y(n_416) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g411 ( .A(n_292), .B(n_303), .Y(n_411) );
INVx1_ASAP7_75t_L g326 ( .A(n_294), .Y(n_326) );
AND2x2_ASAP7_75t_L g311 ( .A(n_295), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AOI31xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .A3(n_306), .B(n_308), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_301), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g434 ( .A(n_301), .B(n_380), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g379 ( .A(n_303), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g405 ( .A(n_303), .Y(n_405) );
INVxp67_ASAP7_75t_L g374 ( .A(n_304), .Y(n_374) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g312 ( .A(n_308), .Y(n_312) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND3xp33_ASAP7_75t_SL g313 ( .A(n_314), .B(n_330), .C(n_346), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_323), .B1(n_327), .B2(n_328), .Y(n_314) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx2_ASAP7_75t_L g400 ( .A(n_317), .Y(n_400) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_321), .Y(n_380) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_321), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_321), .B(n_390), .Y(n_407) );
NAND2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g358 ( .A(n_325), .Y(n_358) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B1(n_341), .B2(n_342), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_333), .B(n_336), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_339), .A2(n_344), .B1(n_378), .B2(n_379), .C(n_381), .Y(n_377) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2x1_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g417 ( .A(n_344), .Y(n_417) );
AND2x2_ASAP7_75t_L g354 ( .A(n_345), .B(n_355), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_SL g402 ( .A1(n_345), .A2(n_403), .B(n_407), .C(n_408), .Y(n_402) );
AOI211xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B(n_351), .C(n_356), .Y(n_346) );
AND2x2_ASAP7_75t_L g397 ( .A(n_350), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g408 ( .A(n_355), .Y(n_408) );
AOI21xp33_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_358), .B(n_359), .Y(n_356) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
NOR3xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_387), .C(n_422), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_363), .B(n_377), .Y(n_362) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g386 ( .A(n_371), .Y(n_386) );
INVxp67_ASAP7_75t_L g410 ( .A(n_375), .Y(n_410) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g394 ( .A(n_384), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B1(n_394), .B2(n_395), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B(n_402), .Y(n_396) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g435 ( .A(n_420), .B(n_436), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_426), .B2(n_429), .C(n_432), .Y(n_422) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI31xp33_ASAP7_75t_SL g432 ( .A1(n_433), .A2(n_434), .A3(n_435), .B(n_437), .Y(n_432) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx4_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx3_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_442), .A2(n_449), .B1(n_782), .B2(n_793), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
AND2x6_ASAP7_75t_SL g443 ( .A(n_444), .B(n_445), .Y(n_443) );
OR2x6_ASAP7_75t_SL g782 ( .A(n_444), .B(n_783), .Y(n_782) );
OR2x2_ASAP7_75t_L g797 ( .A(n_444), .B(n_445), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_444), .B(n_783), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_445), .Y(n_783) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND3x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_669), .C(n_746), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_621), .Y(n_450) );
NOR2xp67_ASAP7_75t_L g451 ( .A(n_452), .B(n_561), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_498), .B1(n_505), .B2(n_554), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_474), .Y(n_453) );
NOR2xp67_ASAP7_75t_SL g604 ( .A(n_454), .B(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_L g619 ( .A(n_454), .B(n_620), .Y(n_619) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_454), .B(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_SL g676 ( .A(n_454), .B(n_677), .Y(n_676) );
INVx4_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_455), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_455), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g611 ( .A(n_455), .Y(n_611) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_455), .Y(n_616) );
AND2x2_ASAP7_75t_L g645 ( .A(n_455), .B(n_585), .Y(n_645) );
OR2x2_ASAP7_75t_L g649 ( .A(n_455), .B(n_490), .Y(n_649) );
AND2x4_ASAP7_75t_L g662 ( .A(n_455), .B(n_620), .Y(n_662) );
NOR2x1_ASAP7_75t_SL g664 ( .A(n_455), .B(n_477), .Y(n_664) );
AND2x2_ASAP7_75t_L g692 ( .A(n_455), .B(n_570), .Y(n_692) );
OR2x6_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVxp67_ASAP7_75t_L g551 ( .A(n_459), .Y(n_551) );
NOR2x1p5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g526 ( .A(n_462), .Y(n_526) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x6_ASAP7_75t_L g466 ( .A(n_463), .B(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_466), .A2(n_481), .B1(n_482), .B2(n_483), .Y(n_480) );
INVxp67_ASAP7_75t_L g542 ( .A(n_466), .Y(n_542) );
INVx2_ASAP7_75t_L g580 ( .A(n_466), .Y(n_580) );
AND2x2_ASAP7_75t_L g471 ( .A(n_467), .B(n_472), .Y(n_471) );
INVxp33_ASAP7_75t_L g525 ( .A(n_467), .Y(n_525) );
INVx1_ASAP7_75t_L g553 ( .A(n_470), .Y(n_553) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g573 ( .A(n_471), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_473), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_474), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_475), .A2(n_750), .B1(n_752), .B2(n_755), .Y(n_749) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_490), .Y(n_475) );
INVx1_ASAP7_75t_L g504 ( .A(n_476), .Y(n_504) );
AND2x2_ASAP7_75t_L g607 ( .A(n_476), .B(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g612 ( .A(n_476), .B(n_570), .Y(n_612) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g569 ( .A(n_477), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g585 ( .A(n_477), .Y(n_585) );
AND2x2_ASAP7_75t_L g618 ( .A(n_477), .B(n_490), .Y(n_618) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_484), .B(n_489), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_483), .B(n_544), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_484) );
INVx2_ASAP7_75t_L g502 ( .A(n_490), .Y(n_502) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_490), .Y(n_587) );
INVx1_ASAP7_75t_L g606 ( .A(n_490), .Y(n_606) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_490), .Y(n_675) );
INVx1_ASAP7_75t_L g687 ( .A(n_490), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI31xp33_ASAP7_75t_SL g741 ( .A1(n_499), .A2(n_742), .A3(n_743), .B(n_744), .Y(n_741) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_503), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g666 ( .A(n_501), .B(n_568), .Y(n_666) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g582 ( .A(n_502), .Y(n_582) );
AND2x4_ASAP7_75t_SL g702 ( .A(n_504), .B(n_606), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_505), .A2(n_623), .B(n_626), .Y(n_622) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
INVx2_ASAP7_75t_L g595 ( .A(n_506), .Y(n_595) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2x1p5_ASAP7_75t_L g722 ( .A(n_507), .B(n_630), .Y(n_722) );
BUFx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g632 ( .A(n_508), .B(n_538), .Y(n_632) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVxp67_ASAP7_75t_L g557 ( .A(n_509), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_509), .B(n_518), .Y(n_592) );
AND2x4_ASAP7_75t_L g602 ( .A(n_509), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g647 ( .A(n_509), .B(n_539), .Y(n_647) );
INVx2_ASAP7_75t_L g655 ( .A(n_509), .Y(n_655) );
INVx1_ASAP7_75t_L g754 ( .A(n_509), .Y(n_754) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_509), .Y(n_763) );
INVx1_ASAP7_75t_L g700 ( .A(n_515), .Y(n_700) );
NAND2x1p5_ASAP7_75t_L g515 ( .A(n_516), .B(n_529), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g556 ( .A(n_517), .B(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_L g695 ( .A(n_517), .B(n_630), .Y(n_695) );
AND2x2_ASAP7_75t_L g712 ( .A(n_517), .B(n_530), .Y(n_712) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_518), .B(n_560), .Y(n_735) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_528), .Y(n_518) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_519), .A2(n_520), .B(n_528), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_521), .B(n_527), .Y(n_520) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g658 ( .A(n_529), .B(n_556), .Y(n_658) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_538), .Y(n_529) );
INVx2_ASAP7_75t_L g564 ( .A(n_530), .Y(n_564) );
NOR2xp67_ASAP7_75t_L g745 ( .A(n_530), .B(n_538), .Y(n_745) );
NOR2x1_ASAP7_75t_L g753 ( .A(n_530), .B(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AND2x2_ASAP7_75t_L g661 ( .A(n_538), .B(n_565), .Y(n_661) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_539), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g590 ( .A(n_539), .Y(n_590) );
AND2x4_ASAP7_75t_L g654 ( .A(n_539), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g684 ( .A(n_539), .Y(n_684) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_547), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_551), .B1(n_552), .B2(n_553), .Y(n_547) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_555), .A2(n_568), .B1(n_706), .B2(n_707), .C(n_708), .Y(n_705) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
AND2x2_ASAP7_75t_L g682 ( .A(n_556), .B(n_683), .Y(n_682) );
BUFx2_ASAP7_75t_L g725 ( .A(n_556), .Y(n_725) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g668 ( .A(n_559), .B(n_592), .Y(n_668) );
INVx3_ASAP7_75t_L g630 ( .A(n_560), .Y(n_630) );
AND2x2_ASAP7_75t_L g762 ( .A(n_560), .B(n_763), .Y(n_762) );
NAND3xp33_ASAP7_75t_SL g561 ( .A(n_562), .B(n_593), .C(n_609), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_566), .B1(n_583), .B2(n_588), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_563), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g693 ( .A(n_563), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g704 ( .A(n_563), .B(n_599), .Y(n_704) );
AND2x2_ASAP7_75t_L g774 ( .A(n_563), .B(n_647), .Y(n_774) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g603 ( .A(n_565), .Y(n_603) );
INVx1_ASAP7_75t_L g652 ( .A(n_565), .Y(n_652) );
INVxp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI222xp33_ASAP7_75t_L g719 ( .A1(n_567), .A2(n_720), .B1(n_721), .B2(n_723), .C1(n_724), .C2(n_726), .Y(n_719) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_581), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_568), .B(n_595), .Y(n_594) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_568), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g686 ( .A(n_569), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g742 ( .A(n_569), .B(n_616), .Y(n_742) );
INVx2_ASAP7_75t_L g608 ( .A(n_570), .Y(n_608) );
INVx1_ASAP7_75t_L g620 ( .A(n_570), .Y(n_620) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_570), .Y(n_677) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_576), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .C(n_575), .Y(n_572) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_582), .Y(n_625) );
INVx3_ASAP7_75t_L g644 ( .A(n_582), .Y(n_644) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g710 ( .A(n_584), .Y(n_710) );
NAND2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g697 ( .A(n_586), .Y(n_697) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g698 ( .A(n_589), .Y(n_698) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g599 ( .A(n_590), .Y(n_599) );
AND2x2_ASAP7_75t_L g717 ( .A(n_590), .B(n_602), .Y(n_717) );
AND2x2_ASAP7_75t_L g780 ( .A(n_590), .B(n_712), .Y(n_780) );
AND2x2_ASAP7_75t_L g709 ( .A(n_591), .B(n_629), .Y(n_709) );
INVx1_ASAP7_75t_L g720 ( .A(n_591), .Y(n_720) );
AND2x2_ASAP7_75t_L g737 ( .A(n_591), .B(n_684), .Y(n_737) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_596), .B1(n_600), .B2(n_604), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_596), .A2(n_610), .B(n_613), .Y(n_609) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g641 ( .A(n_599), .B(n_602), .Y(n_641) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x4_ASAP7_75t_L g744 ( .A(n_602), .B(n_745), .Y(n_744) );
BUFx2_ASAP7_75t_L g707 ( .A(n_605), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_606), .Y(n_635) );
AND2x2_ASAP7_75t_SL g615 ( .A(n_607), .B(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g680 ( .A(n_607), .Y(n_680) );
AND2x2_ASAP7_75t_L g778 ( .A(n_607), .B(n_675), .Y(n_778) );
INVx1_ASAP7_75t_L g733 ( .A(n_608), .Y(n_733) );
INVx1_ASAP7_75t_L g639 ( .A(n_610), .Y(n_639) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g728 ( .A(n_611), .Y(n_728) );
INVx4_ASAP7_75t_L g637 ( .A(n_612), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI32xp33_ASAP7_75t_L g708 ( .A1(n_615), .A2(n_709), .A3(n_710), .B1(n_711), .B2(n_712), .Y(n_708) );
AND2x2_ASAP7_75t_L g703 ( .A(n_616), .B(n_618), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_SL g766 ( .A1(n_616), .A2(n_767), .B(n_768), .C(n_770), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_SL g731 ( .A(n_618), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g770 ( .A(n_618), .Y(n_770) );
AND2x2_ASAP7_75t_L g624 ( .A(n_619), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g751 ( .A(n_619), .Y(n_751) );
AND2x2_ASAP7_75t_L g757 ( .A(n_619), .B(n_644), .Y(n_757) );
NOR3x1_ASAP7_75t_L g621 ( .A(n_622), .B(n_638), .C(n_656), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_633), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
AND2x2_ASAP7_75t_L g646 ( .A(n_629), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g689 ( .A(n_629), .B(n_654), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_629), .B(n_675), .Y(n_716) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_637), .B(n_644), .Y(n_743) );
INVx2_ASAP7_75t_L g765 ( .A(n_637), .Y(n_765) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B(n_642), .Y(n_638) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_639), .A2(n_730), .B1(n_734), .B2(n_736), .C(n_741), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_640), .A2(n_760), .B1(n_761), .B2(n_764), .Y(n_759) );
INVx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B1(n_648), .B2(n_650), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
AND2x2_ASAP7_75t_L g688 ( .A(n_644), .B(n_664), .Y(n_688) );
INVx1_ASAP7_75t_L g694 ( .A(n_644), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_644), .B(n_662), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_647), .B(n_715), .Y(n_781) );
NAND2x1_ASAP7_75t_L g764 ( .A(n_648), .B(n_765), .Y(n_764) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
NOR2x1_ASAP7_75t_L g679 ( .A(n_649), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
NAND2x1_ASAP7_75t_SL g767 ( .A(n_652), .B(n_654), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_652), .B(n_752), .Y(n_773) );
OR2x2_ASAP7_75t_L g734 ( .A(n_653), .B(n_735), .Y(n_734) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g769 ( .A(n_654), .B(n_695), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_657), .B(n_663), .Y(n_656) );
OAI21xp33_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_659), .B(n_662), .Y(n_657) );
OR2x2_ASAP7_75t_L g721 ( .A(n_660), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g755 ( .A(n_661), .B(n_753), .Y(n_755) );
AND2x2_ASAP7_75t_SL g701 ( .A(n_662), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g711 ( .A(n_662), .Y(n_711) );
OAI21xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B(n_667), .Y(n_663) );
AND2x2_ASAP7_75t_L g696 ( .A(n_664), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_713), .Y(n_670) );
NOR3xp33_ASAP7_75t_SL g671 ( .A(n_672), .B(n_690), .C(n_705), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_678), .B(n_681), .C(n_685), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g739 ( .A(n_684), .Y(n_739) );
AND2x2_ASAP7_75t_L g752 ( .A(n_684), .B(n_753), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g760 ( .A(n_686), .Y(n_760) );
OAI21xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_698), .B(n_699), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_695), .B2(n_696), .Y(n_691) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_692), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_703), .B2(n_704), .Y(n_699) );
INVx1_ASAP7_75t_SL g706 ( .A(n_704), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_710), .B(n_751), .Y(n_750) );
OAI22xp33_ASAP7_75t_SL g776 ( .A1(n_711), .A2(n_777), .B1(n_779), .B2(n_781), .Y(n_776) );
AOI211x1_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_718), .B(n_719), .C(n_729), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_731), .A2(n_772), .B(n_774), .Y(n_771) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g740 ( .A(n_735), .Y(n_740) );
NOR2xp67_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_738), .B(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND4xp25_ASAP7_75t_L g747 ( .A(n_748), .B(n_758), .C(n_771), .D(n_775), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_756), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_766), .Y(n_758) );
INVxp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_803), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_803), .A2(n_808), .B(n_818), .Y(n_807) );
INVx1_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
BUFx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
BUFx2_ASAP7_75t_L g820 ( .A(n_806), .Y(n_820) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g817 ( .A(n_813), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
endmodule