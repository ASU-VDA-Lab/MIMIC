module fake_jpeg_19479_n_346 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_48),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_22),
.B(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_49),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_16),
.C(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_51),
.Y(n_74)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_68),
.B(n_24),
.Y(n_109)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_15),
.B1(n_25),
.B2(n_35),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_74),
.B(n_81),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_40),
.B1(n_39),
.B2(n_41),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_75),
.A2(n_101),
.B1(n_104),
.B2(n_32),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_44),
.C(n_16),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_42),
.B(n_48),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_77),
.B(n_111),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_80),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_50),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_83),
.B(n_93),
.Y(n_121)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_87),
.B1(n_91),
.B2(n_36),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_15),
.B1(n_25),
.B2(n_35),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_100),
.Y(n_123)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_102),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_31),
.B(n_29),
.C(n_32),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_39),
.B1(n_19),
.B2(n_24),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_57),
.A2(n_46),
.B1(n_47),
.B2(n_45),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_47),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_47),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_110),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_22),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_36),
.B1(n_38),
.B2(n_45),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_45),
.B1(n_38),
.B2(n_36),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_135),
.B1(n_89),
.B2(n_82),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_75),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_118),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_36),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_122),
.A2(n_86),
.B1(n_88),
.B2(n_33),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_134),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_44),
.C(n_30),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_141),
.B1(n_94),
.B2(n_84),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_96),
.A2(n_98),
.B1(n_100),
.B2(n_97),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_91),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_106),
.Y(n_150)
);

BUFx16f_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_160),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_152),
.B(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_112),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_163),
.B1(n_166),
.B2(n_169),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_121),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_168),
.Y(n_184)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_162),
.Y(n_178)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_127),
.A2(n_73),
.B1(n_84),
.B2(n_85),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_136),
.C(n_122),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_173),
.B1(n_113),
.B2(n_131),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_127),
.A2(n_85),
.B1(n_72),
.B2(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_167),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_95),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_77),
.B1(n_103),
.B2(n_44),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_170),
.A2(n_138),
.B1(n_141),
.B2(n_144),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_22),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_142),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_129),
.B(n_103),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_172),
.B(n_131),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_173)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_26),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_141),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_179),
.B(n_0),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_192),
.C(n_194),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_154),
.B1(n_161),
.B2(n_28),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_185),
.B(n_187),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_203),
.B1(n_13),
.B2(n_12),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_142),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_142),
.B1(n_141),
.B2(n_144),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_188),
.A2(n_202),
.B1(n_20),
.B2(n_1),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_150),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_199),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_131),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_130),
.C(n_78),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_167),
.B(n_92),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_197),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_153),
.B(n_78),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_157),
.C(n_155),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_124),
.B1(n_11),
.B2(n_13),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_169),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_145),
.B(n_143),
.C(n_30),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_30),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_148),
.B1(n_173),
.B2(n_149),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_211),
.B1(n_225),
.B2(n_227),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_162),
.B(n_160),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_209),
.A2(n_220),
.B(n_234),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_213),
.B(n_194),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_217),
.B1(n_233),
.B2(n_215),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_23),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_228),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_20),
.Y(n_223)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

NOR2x1_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_181),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_20),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_3),
.B(n_4),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_229),
.A2(n_193),
.B1(n_175),
.B2(n_176),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_199),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_191),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_232),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_5),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_235),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_180),
.A2(n_6),
.B(n_7),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_7),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_245),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_255),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_208),
.B(n_185),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_250),
.Y(n_268)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_178),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_186),
.C(n_181),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_208),
.C(n_219),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_210),
.B(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_206),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_226),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_253),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_220),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_207),
.B1(n_225),
.B2(n_220),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_213),
.Y(n_275)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_260),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_193),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_262),
.A2(n_264),
.B1(n_275),
.B2(n_236),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_247),
.A2(n_234),
.B1(n_228),
.B2(n_232),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_244),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_241),
.A2(n_216),
.B1(n_235),
.B2(n_227),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_276),
.B1(n_277),
.B2(n_239),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_219),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_272),
.B(n_254),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_241),
.A2(n_230),
.B1(n_205),
.B2(n_10),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_245),
.A2(n_205),
.B1(n_9),
.B2(n_10),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_8),
.Y(n_278)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_10),
.C(n_8),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_236),
.C(n_242),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_8),
.Y(n_282)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_288),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_251),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_287),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_261),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_290),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_292),
.B(n_277),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_259),
.C(n_237),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_281),
.C(n_272),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_254),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_297),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_295),
.A2(n_262),
.B1(n_279),
.B2(n_266),
.Y(n_312)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_300),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_243),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_263),
.A2(n_260),
.B1(n_240),
.B2(n_249),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_298),
.B(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_257),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_289),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_280),
.C(n_273),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_302),
.B(n_313),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_271),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_294),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_312),
.Y(n_320)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_315),
.B(n_301),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_285),
.Y(n_321)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_322),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_297),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_317),
.A2(n_283),
.B(n_295),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_327),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_318),
.B(n_302),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_307),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_329),
.B(n_314),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_333),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_330),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_315),
.B(n_307),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_336),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_334),
.A2(n_324),
.B(n_326),
.Y(n_337)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_337),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_339),
.B(n_338),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_303),
.B(n_320),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_342),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_303),
.B(n_325),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_344),
.B(n_325),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_276),
.B1(n_288),
.B2(n_319),
.Y(n_346)
);


endmodule