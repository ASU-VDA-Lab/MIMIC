module fake_jpeg_1050_n_685 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_685);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_685;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_19),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_61),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_63),
.Y(n_142)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_65),
.B(n_79),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_21),
.A2(n_35),
.B1(n_26),
.B2(n_58),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_66),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_68),
.Y(n_199)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_69),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_22),
.B(n_8),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_70),
.B(n_81),
.Y(n_143)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g210 ( 
.A(n_76),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_48),
.Y(n_78)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_78),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_27),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_80),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_28),
.B(n_9),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_9),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_85),
.B(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_22),
.B(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_24),
.B(n_9),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_87),
.B(n_101),
.Y(n_171)
);

BUFx4f_ASAP7_75t_SL g88 ( 
.A(n_37),
.Y(n_88)
);

CKINVDCx6p67_ASAP7_75t_R g181 ( 
.A(n_88),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_23),
.A2(n_7),
.B(n_17),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_89),
.B(n_39),
.C(n_29),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_90),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g213 ( 
.A(n_91),
.Y(n_213)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_92),
.Y(n_215)
);

BUFx4f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_93),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_94),
.B(n_105),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_97),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_100),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_11),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_103),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_49),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_106),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_24),
.B(n_6),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_107),
.B(n_113),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_49),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_108),
.B(n_109),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_49),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_51),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_112),
.B(n_123),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_18),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_18),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_114),
.B(n_117),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_116),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_43),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_40),
.B(n_6),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_118),
.B(n_12),
.Y(n_193)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_59),
.B(n_0),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_59),
.Y(n_135)
);

BUFx16f_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_122),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_58),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

BUFx2_ASAP7_75t_SL g203 ( 
.A(n_124),
.Y(n_203)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_126),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_127),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_58),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_128),
.B(n_35),
.Y(n_166)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_31),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_129),
.Y(n_216)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_26),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_42),
.Y(n_132)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_134),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_135),
.B(n_72),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_66),
.A2(n_26),
.B1(n_35),
.B2(n_52),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_136),
.A2(n_145),
.B1(n_146),
.B2(n_168),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_52),
.B1(n_26),
.B2(n_35),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_78),
.A2(n_53),
.B1(n_43),
.B2(n_40),
.Y(n_146)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_154),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_93),
.A2(n_52),
.B1(n_41),
.B2(n_44),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_157),
.A2(n_173),
.B1(n_201),
.B2(n_204),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_57),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_164),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_63),
.A2(n_53),
.B1(n_57),
.B2(n_56),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_165),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_166),
.B(n_3),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_89),
.A2(n_20),
.B1(n_50),
.B2(n_39),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_64),
.B(n_56),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_172),
.B(n_61),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_93),
.A2(n_41),
.B1(n_44),
.B2(n_50),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_175),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_95),
.A2(n_50),
.B1(n_20),
.B2(n_39),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_178),
.A2(n_185),
.B1(n_219),
.B2(n_220),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_L g303 ( 
.A1(n_179),
.A2(n_211),
.B(n_141),
.Y(n_303)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_98),
.A2(n_44),
.B1(n_41),
.B2(n_20),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_99),
.A2(n_30),
.B1(n_29),
.B2(n_33),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_186),
.A2(n_189),
.B1(n_190),
.B2(n_1),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_103),
.A2(n_30),
.B1(n_29),
.B2(n_33),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_104),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_190)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_193),
.B(n_221),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_97),
.B(n_38),
.C(n_37),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_194),
.B(n_91),
.C(n_77),
.Y(n_251)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_76),
.A2(n_32),
.B1(n_38),
.B2(n_37),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_69),
.Y(n_202)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_202),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_83),
.A2(n_32),
.B1(n_37),
.B2(n_12),
.Y(n_204)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_205),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_80),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_211),
.B1(n_222),
.B2(n_90),
.Y(n_236)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_115),
.Y(n_208)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_208),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_122),
.A2(n_84),
.B1(n_126),
.B2(n_116),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_120),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_88),
.B(n_5),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_92),
.A2(n_129),
.B1(n_119),
.B2(n_100),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_159),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_227),
.B(n_228),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_174),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_88),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_229),
.B(n_230),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_135),
.B(n_110),
.Y(n_230)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_232),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_168),
.B(n_110),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_233),
.B(n_254),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_234),
.B(n_241),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_236),
.Y(n_342)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_147),
.Y(n_239)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_240),
.B(n_251),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_187),
.Y(n_241)
);

BUFx4f_ASAP7_75t_SL g242 ( 
.A(n_223),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_242),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_243),
.B(n_262),
.Y(n_359)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_142),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_244),
.Y(n_351)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

INVx11_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

BUFx2_ASAP7_75t_SL g249 ( 
.A(n_181),
.Y(n_249)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_136),
.A2(n_127),
.B1(n_68),
.B2(n_91),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_250),
.A2(n_150),
.B1(n_151),
.B2(n_225),
.Y(n_308)
);

AND2x4_ASAP7_75t_SL g253 ( 
.A(n_158),
.B(n_124),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_253),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_183),
.B(n_0),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_203),
.A2(n_5),
.B1(n_15),
.B2(n_13),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_255),
.A2(n_258),
.B1(n_259),
.B2(n_271),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_256),
.A2(n_262),
.B1(n_244),
.B2(n_253),
.Y(n_358)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_133),
.Y(n_257)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_181),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_259)
);

OA22x2_ASAP7_75t_SL g260 ( 
.A1(n_181),
.A2(n_3),
.B1(n_4),
.B2(n_15),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_260),
.A2(n_188),
.B(n_195),
.C(n_198),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_143),
.B(n_3),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_261),
.B(n_295),
.Y(n_334)
);

INVx4_ASAP7_75t_SL g262 ( 
.A(n_223),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_263),
.B(n_267),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_137),
.B(n_17),
.C(n_4),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_264),
.B(n_288),
.C(n_207),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_149),
.B(n_4),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_155),
.Y(n_268)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_268),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_171),
.B(n_177),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_269),
.B(n_279),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_191),
.A2(n_172),
.B1(n_142),
.B2(n_170),
.Y(n_271)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_133),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_197),
.Y(n_273)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_163),
.Y(n_274)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

OR2x4_ASAP7_75t_L g275 ( 
.A(n_160),
.B(n_178),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_SL g326 ( 
.A(n_275),
.B(n_293),
.Y(n_326)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_277),
.Y(n_330)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_138),
.Y(n_278)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_160),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_192),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_280),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_144),
.B(n_140),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_281),
.B(n_289),
.Y(n_348)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_226),
.Y(n_282)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_282),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_190),
.A2(n_189),
.B1(n_186),
.B2(n_157),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_283),
.A2(n_304),
.B1(n_250),
.B2(n_301),
.Y(n_345)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_223),
.Y(n_284)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_284),
.Y(n_343)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_210),
.Y(n_285)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_199),
.Y(n_286)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_170),
.A2(n_163),
.B1(n_201),
.B2(n_216),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_287),
.A2(n_302),
.B1(n_225),
.B2(n_207),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_152),
.B(n_153),
.C(n_156),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_176),
.B(n_196),
.Y(n_289)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_291),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_292),
.Y(n_319)
);

OR2x4_ASAP7_75t_L g293 ( 
.A(n_206),
.B(n_204),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_224),
.B(n_180),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_294),
.B(n_299),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_184),
.B(n_162),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_162),
.Y(n_296)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_218),
.Y(n_297)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_214),
.A2(n_217),
.B1(n_215),
.B2(n_213),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_188),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_214),
.B(n_213),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_217),
.Y(n_300)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_300),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_134),
.B(n_208),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_212),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_173),
.A2(n_222),
.B1(n_161),
.B2(n_167),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_303),
.B(n_305),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_154),
.A2(n_205),
.B1(n_182),
.B2(n_148),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_138),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_141),
.B(n_148),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_307),
.B(n_257),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_308),
.A2(n_331),
.B1(n_313),
.B2(n_336),
.Y(n_415)
);

AOI211xp5_ASAP7_75t_SL g317 ( 
.A1(n_275),
.A2(n_161),
.B(n_151),
.C(n_150),
.Y(n_317)
);

AO21x1_ASAP7_75t_L g373 ( 
.A1(n_317),
.A2(n_321),
.B(n_358),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_233),
.A2(n_237),
.B1(n_258),
.B2(n_283),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_318),
.A2(n_337),
.B1(n_362),
.B2(n_238),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_321),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_323),
.B(n_338),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_303),
.A2(n_195),
.B(n_198),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_324),
.A2(n_272),
.B(n_278),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_260),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_325),
.B(n_332),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_260),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_333),
.A2(n_357),
.B1(n_245),
.B2(n_284),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_335),
.B(n_353),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_237),
.A2(n_212),
.B1(n_231),
.B2(n_293),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_254),
.B(n_246),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_355),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_345),
.A2(n_349),
.B1(n_265),
.B2(n_290),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_231),
.A2(n_235),
.B1(n_251),
.B2(n_229),
.Y(n_349)
);

A2O1A1Ixp33_ASAP7_75t_L g353 ( 
.A1(n_230),
.A2(n_248),
.B(n_240),
.C(n_261),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_295),
.B(n_243),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_240),
.A2(n_304),
.B1(n_253),
.B2(n_252),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_270),
.Y(n_391)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_298),
.A2(n_306),
.B1(n_238),
.B2(n_273),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_360),
.A2(n_308),
.B1(n_364),
.B2(n_317),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_288),
.A2(n_232),
.B1(n_305),
.B2(n_306),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_264),
.B(n_239),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_286),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_368),
.B(n_247),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_326),
.A2(n_276),
.B(n_266),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_370),
.A2(n_375),
.B(n_376),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_371),
.A2(n_381),
.B1(n_406),
.B2(n_408),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_373),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_326),
.A2(n_277),
.B(n_296),
.Y(n_375)
);

NOR2x1_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_282),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_368),
.Y(n_378)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_378),
.Y(n_420)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_379),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_380),
.A2(n_391),
.B(n_401),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_345),
.A2(n_311),
.B1(n_349),
.B2(n_332),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_312),
.B(n_268),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_384),
.B(n_389),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_385),
.A2(n_395),
.B1(n_411),
.B2(n_415),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_386),
.B(n_418),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_320),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_387),
.B(n_390),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_334),
.B(n_265),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_320),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_344),
.Y(n_392)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_392),
.Y(n_433)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_393),
.Y(n_453)
);

INVx8_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_394),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_311),
.A2(n_290),
.B1(n_247),
.B2(n_291),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_396),
.B(n_399),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_274),
.C(n_270),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_413),
.C(n_404),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_398),
.A2(n_405),
.B1(n_409),
.B2(n_416),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_312),
.B(n_242),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_334),
.B(n_242),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_400),
.B(n_402),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_355),
.B(n_341),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_363),
.B(n_245),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_403),
.B(n_404),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_367),
.B(n_335),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_325),
.A2(n_324),
.B1(n_347),
.B2(n_350),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_353),
.A2(n_350),
.B(n_316),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_407),
.A2(n_362),
.B(n_319),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_347),
.A2(n_350),
.B1(n_342),
.B2(n_321),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_339),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_340),
.Y(n_410)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_410),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_338),
.A2(n_310),
.B1(n_323),
.B2(n_356),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_359),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_412),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_310),
.B(n_356),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_359),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_414),
.Y(n_421)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_339),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_369),
.B(n_327),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_417),
.A2(n_390),
.B(n_387),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_348),
.B(n_363),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_422),
.B(n_425),
.Y(n_484)
);

XNOR2x1_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_348),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_408),
.A2(n_369),
.B1(n_327),
.B2(n_322),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_430),
.A2(n_434),
.B(n_445),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_384),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_431),
.B(n_436),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_388),
.B(n_413),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_449),
.C(n_452),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_399),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_456),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_385),
.A2(n_331),
.B1(n_336),
.B2(n_319),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_443),
.A2(n_415),
.B1(n_395),
.B2(n_392),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_382),
.A2(n_322),
.B(n_313),
.Y(n_445)
);

MAJx2_ASAP7_75t_L g449 ( 
.A(n_388),
.B(n_365),
.C(n_346),
.Y(n_449)
);

AOI22x1_ASAP7_75t_SL g450 ( 
.A1(n_381),
.A2(n_346),
.B1(n_343),
.B2(n_329),
.Y(n_450)
);

OAI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_450),
.A2(n_373),
.B1(n_401),
.B2(n_376),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_407),
.A2(n_375),
.B(n_370),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_383),
.B(n_365),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_377),
.A2(n_336),
.B1(n_315),
.B2(n_330),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_454),
.A2(n_458),
.B1(n_405),
.B2(n_379),
.Y(n_468)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_382),
.A2(n_352),
.B(n_315),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_455),
.B(n_398),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_386),
.B(n_354),
.C(n_330),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_383),
.B(n_354),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_457),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_377),
.A2(n_352),
.B1(n_309),
.B2(n_314),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_402),
.B(n_343),
.C(n_314),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_459),
.B(n_393),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_423),
.A2(n_406),
.B1(n_372),
.B2(n_412),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_460),
.A2(n_472),
.B(n_485),
.Y(n_501)
);

A2O1A1Ixp33_ASAP7_75t_SL g521 ( 
.A1(n_461),
.A2(n_480),
.B(n_439),
.C(n_444),
.Y(n_521)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_428),
.Y(n_462)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_463),
.B(n_422),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_419),
.A2(n_414),
.B1(n_371),
.B2(n_411),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_465),
.A2(n_469),
.B1(n_477),
.B2(n_482),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_438),
.A2(n_378),
.B1(n_380),
.B2(n_389),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_466),
.A2(n_424),
.B1(n_454),
.B2(n_420),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_468),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_424),
.A2(n_391),
.B1(n_396),
.B2(n_400),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_428),
.Y(n_470)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_470),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_419),
.B(n_397),
.Y(n_471)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_471),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_426),
.A2(n_391),
.B(n_373),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_421),
.B(n_397),
.Y(n_473)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_473),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_421),
.B(n_417),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_474),
.B(n_478),
.Y(n_509)
);

INVx6_ASAP7_75t_L g475 ( 
.A(n_448),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_475),
.Y(n_507)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_433),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_476),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g480 ( 
.A1(n_429),
.A2(n_376),
.B(n_416),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_431),
.B(n_418),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_481),
.B(n_486),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_438),
.A2(n_403),
.B1(n_409),
.B2(n_394),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_423),
.A2(n_410),
.B1(n_374),
.B2(n_329),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_433),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_445),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_488),
.B(n_489),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_455),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_437),
.B(n_374),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_490),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_455),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_491),
.Y(n_529)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_453),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_493),
.Y(n_506)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_453),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_420),
.A2(n_394),
.B1(n_410),
.B2(n_328),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_494),
.A2(n_446),
.B1(n_448),
.B2(n_328),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_432),
.B(n_309),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_496),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_455),
.Y(n_496)
);

AO21x1_ASAP7_75t_L g537 ( 
.A1(n_499),
.A2(n_502),
.B(n_508),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_479),
.A2(n_429),
.B(n_451),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_467),
.B(n_440),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g540 ( 
.A(n_503),
.B(n_505),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_489),
.A2(n_427),
.B1(n_432),
.B2(n_447),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_504),
.A2(n_526),
.B1(n_480),
.B2(n_466),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_472),
.A2(n_434),
.B(n_426),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g510 ( 
.A1(n_461),
.A2(n_436),
.B(n_439),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_510),
.B(n_480),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_464),
.A2(n_447),
.B1(n_458),
.B2(n_443),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_511),
.A2(n_525),
.B1(n_469),
.B2(n_468),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_484),
.B(n_449),
.C(n_457),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_512),
.B(n_514),
.C(n_531),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_484),
.B(n_467),
.C(n_483),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_483),
.B(n_425),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g552 ( 
.A(n_515),
.B(n_480),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_441),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_516),
.B(n_520),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_459),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_521),
.A2(n_527),
.B(n_485),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_471),
.B(n_435),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_524),
.B(n_532),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_464),
.A2(n_444),
.B1(n_452),
.B2(n_450),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_491),
.A2(n_430),
.B1(n_435),
.B2(n_456),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_497),
.A2(n_442),
.B(n_351),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_473),
.B(n_442),
.C(n_351),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_481),
.B(n_463),
.Y(n_532)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_534),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_505),
.B(n_474),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_536),
.B(n_547),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_519),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_538),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_541),
.A2(n_555),
.B(n_521),
.Y(n_585)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_506),
.Y(n_542)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_542),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_495),
.Y(n_543)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_543),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_533),
.Y(n_545)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_545),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_546),
.A2(n_548),
.B1(n_554),
.B2(n_558),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_523),
.B(n_488),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_519),
.Y(n_548)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_509),
.Y(n_549)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_549),
.Y(n_579)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_513),
.Y(n_550)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_550),
.Y(n_593)
);

A2O1A1O1Ixp25_ASAP7_75t_L g551 ( 
.A1(n_502),
.A2(n_496),
.B(n_497),
.C(n_461),
.D(n_460),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_551),
.A2(n_560),
.B(n_566),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_552),
.B(n_521),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_553),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_518),
.A2(n_482),
.B1(n_477),
.B2(n_490),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_525),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_556),
.B(n_510),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_514),
.B(n_493),
.C(n_492),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_557),
.B(n_512),
.C(n_531),
.Y(n_571)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_533),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_530),
.A2(n_470),
.B(n_486),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_500),
.A2(n_462),
.B1(n_476),
.B2(n_494),
.Y(n_561)
);

OAI22xp33_ASAP7_75t_L g573 ( 
.A1(n_561),
.A2(n_562),
.B1(n_507),
.B2(n_522),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_500),
.A2(n_446),
.B1(n_475),
.B2(n_351),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_532),
.B(n_475),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_563),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_523),
.B(n_361),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_564),
.B(n_504),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_499),
.A2(n_511),
.B1(n_509),
.B2(n_528),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_565),
.B(n_567),
.Y(n_575)
);

AOI21x1_ASAP7_75t_L g566 ( 
.A1(n_530),
.A2(n_361),
.B(n_527),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_522),
.B(n_528),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_571),
.B(n_577),
.Y(n_613)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_573),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_574),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_557),
.B(n_503),
.C(n_524),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_578),
.B(n_542),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_535),
.B(n_526),
.C(n_515),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_580),
.B(n_583),
.C(n_589),
.Y(n_601)
);

BUFx12_ASAP7_75t_L g581 ( 
.A(n_544),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_581),
.Y(n_611)
);

AO221x1_ASAP7_75t_L g582 ( 
.A1(n_554),
.A2(n_507),
.B1(n_521),
.B2(n_510),
.C(n_498),
.Y(n_582)
);

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_582),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_535),
.B(n_501),
.C(n_508),
.Y(n_583)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_585),
.A2(n_567),
.B(n_543),
.Y(n_612)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_559),
.Y(n_588)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_588),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_544),
.B(n_501),
.C(n_517),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_SL g605 ( 
.A(n_591),
.B(n_537),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_541),
.A2(n_521),
.B(n_498),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_592),
.A2(n_566),
.B(n_555),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_545),
.B(n_517),
.Y(n_594)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_594),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_597),
.B(n_612),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_584),
.A2(n_565),
.B1(n_553),
.B2(n_550),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_600),
.A2(n_576),
.B1(n_592),
.B2(n_575),
.Y(n_627)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_602),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_571),
.B(n_540),
.C(n_563),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_604),
.B(n_606),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_605),
.B(n_614),
.Y(n_630)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_594),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_588),
.B(n_546),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_607),
.B(n_608),
.Y(n_629)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_594),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_583),
.B(n_540),
.C(n_558),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_609),
.B(n_616),
.Y(n_622)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_575),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_610),
.B(n_615),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_570),
.B(n_538),
.Y(n_614)
);

XNOR2x1_ASAP7_75t_L g615 ( 
.A(n_589),
.B(n_552),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_568),
.B(n_537),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_570),
.B(n_548),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_617),
.B(n_614),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_613),
.B(n_601),
.C(n_604),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_620),
.B(n_621),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_601),
.B(n_577),
.C(n_584),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_580),
.C(n_586),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_624),
.B(n_626),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_603),
.A2(n_593),
.B1(n_568),
.B2(n_576),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_625),
.A2(n_627),
.B1(n_632),
.B2(n_595),
.Y(n_643)
);

BUFx24_ASAP7_75t_SL g626 ( 
.A(n_598),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_600),
.B(n_590),
.C(n_573),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_628),
.B(n_633),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_603),
.A2(n_569),
.B1(n_575),
.B2(n_579),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_598),
.B(n_593),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_634),
.B(n_579),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_597),
.B(n_572),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_635),
.B(n_636),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_595),
.B(n_585),
.C(n_587),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_622),
.A2(n_612),
.B(n_587),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_637),
.B(n_643),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_619),
.B(n_611),
.Y(n_641)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_641),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_620),
.B(n_596),
.C(n_606),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_644),
.B(n_645),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_621),
.B(n_596),
.C(n_608),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_623),
.A2(n_631),
.B(n_618),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_646),
.A2(n_648),
.B(n_632),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_624),
.B(n_611),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_647),
.B(n_650),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_623),
.A2(n_617),
.B(n_551),
.Y(n_648)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_649),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_636),
.B(n_599),
.C(n_610),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_628),
.B(n_599),
.C(n_615),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_651),
.B(n_627),
.Y(n_657)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_630),
.B(n_605),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_652),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_639),
.B(n_629),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_653),
.B(n_657),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_640),
.B(n_630),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_654),
.B(n_660),
.Y(n_666)
);

AO21x1_ASAP7_75t_L g672 ( 
.A1(n_655),
.A2(n_648),
.B(n_569),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_641),
.B(n_539),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_642),
.B(n_539),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_663),
.B(n_652),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_659),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_665),
.B(n_667),
.Y(n_674)
);

XOR2xp5_ASAP7_75t_L g668 ( 
.A(n_659),
.B(n_651),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_668),
.B(n_671),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_661),
.A2(n_638),
.B(n_649),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_670),
.A2(n_672),
.B(n_673),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g671 ( 
.A(n_658),
.B(n_645),
.C(n_644),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_664),
.A2(n_650),
.B(n_602),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_669),
.A2(n_656),
.B(n_662),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_675),
.A2(n_562),
.B(n_591),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_666),
.B(n_656),
.C(n_560),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_676),
.B(n_561),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_678),
.A2(n_665),
.B(n_672),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_679),
.A2(n_681),
.B(n_677),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_SL g682 ( 
.A(n_680),
.B(n_674),
.Y(n_682)
);

XNOR2xp5_ASAP7_75t_L g684 ( 
.A(n_682),
.B(n_683),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_684),
.A2(n_581),
.B(n_683),
.Y(n_685)
);


endmodule