module fake_jpeg_5140_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_17),
.B1(n_19),
.B2(n_15),
.Y(n_43)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_1),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_1),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_16),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_40),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_17),
.B1(n_27),
.B2(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_44),
.B1(n_29),
.B2(n_34),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_18),
.B1(n_15),
.B2(n_25),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_22),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_61),
.B1(n_63),
.B2(n_41),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_26),
.C(n_23),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_56),
.B(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_54),
.Y(n_82)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_30),
.B(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_13),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_64),
.Y(n_68)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_13),
.B1(n_23),
.B2(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_81),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_58),
.B1(n_54),
.B2(n_67),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_83),
.Y(n_86)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_55),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_94),
.C(n_84),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_39),
.B1(n_32),
.B2(n_31),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_92),
.B1(n_77),
.B2(n_25),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_39),
.B1(n_31),
.B2(n_25),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_83),
.B(n_84),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_93),
.A2(n_84),
.B(n_75),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_1),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_71),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_101),
.C(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_105),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_85),
.Y(n_114)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_77),
.B(n_25),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_106),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_113),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_89),
.C(n_93),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_114),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_116),
.A2(n_104),
.B1(n_103),
.B2(n_108),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_90),
.C(n_94),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_122),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_105),
.B1(n_99),
.B2(n_109),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_115),
.C(n_68),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_123),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_126),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_119),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_6),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_7),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_129),
.A2(n_131),
.B(n_132),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_7),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_124),
.C(n_9),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_133),
.B(n_135),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_9),
.C(n_10),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_134),
.B(n_10),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_136),
.B(n_11),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_12),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_2),
.Y(n_140)
);


endmodule