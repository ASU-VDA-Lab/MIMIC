module fake_jpeg_17581_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_69),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_54),
.B1(n_53),
.B2(n_49),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_52),
.B1(n_45),
.B2(n_50),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_77),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_79),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_54),
.B1(n_61),
.B2(n_44),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_62),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_8),
.B(n_9),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_97),
.B1(n_12),
.B2(n_13),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_91),
.B1(n_100),
.B2(n_104),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_47),
.B1(n_56),
.B2(n_4),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_101),
.Y(n_113)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_7),
.Y(n_106)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

BUFx2_ASAP7_75t_SL g107 ( 
.A(n_98),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

BUFx4f_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_102),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_57),
.B1(n_7),
.B2(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_109),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_11),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_14),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_114),
.B(n_88),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_102),
.B1(n_103),
.B2(n_89),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_95),
.B1(n_107),
.B2(n_99),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_106),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_107),
.B(n_19),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_94),
.C(n_113),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_115),
.C(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_124),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_126),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_18),
.C(n_20),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_127),
.B(n_26),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_133),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_132),
.B1(n_30),
.B2(n_31),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

OAI21x1_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_25),
.B(n_32),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_33),
.B(n_35),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_37),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_41),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_42),
.C(n_43),
.Y(n_144)
);


endmodule