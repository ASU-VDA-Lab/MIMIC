module fake_jpeg_221_n_199 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_199);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_77),
.Y(n_88)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_1),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_79),
.Y(n_90)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_72),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_84),
.Y(n_99)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_53),
.Y(n_98)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_53),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_51),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_97),
.Y(n_103)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_98),
.B(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_108),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_71),
.Y(n_125)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_54),
.B1(n_71),
.B2(n_68),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_70),
.B1(n_56),
.B2(n_58),
.Y(n_126)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_64),
.B(n_55),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_68),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_2),
.C(n_3),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_61),
.B(n_73),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_117),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_54),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_121),
.B(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_2),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_66),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_118),
.C(n_121),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_66),
.B1(n_58),
.B2(n_4),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_158)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_133),
.Y(n_142)
);

AO22x2_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_22),
.B1(n_47),
.B2(n_46),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_3),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_99),
.B(n_6),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_6),
.B(n_7),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_160),
.B(n_26),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_38),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_48),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_45),
.C(n_19),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_151),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_150),
.B(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_162),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_10),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_168)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

AO22x1_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_27),
.B1(n_14),
.B2(n_16),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_11),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_37),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_170),
.B(n_173),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_28),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_171),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_34),
.C(n_35),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_175),
.B(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_176),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_177),
.A2(n_161),
.B1(n_152),
.B2(n_142),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_167),
.B1(n_165),
.B2(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_183),
.A2(n_172),
.B1(n_166),
.B2(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_187),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_173),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_194),
.B1(n_181),
.B2(n_192),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_187),
.B1(n_188),
.B2(n_170),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_184),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_141),
.C(n_155),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_150),
.C(n_164),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_40),
.Y(n_199)
);


endmodule