module real_jpeg_12466_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_1),
.A2(n_59),
.B1(n_63),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_1),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_1),
.A2(n_45),
.B1(n_47),
.B2(n_77),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_1),
.A2(n_34),
.B1(n_40),
.B2(n_77),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_2),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_2),
.A2(n_59),
.B1(n_63),
.B2(n_125),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_2),
.A2(n_45),
.B1(n_47),
.B2(n_125),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_2),
.A2(n_34),
.B1(n_40),
.B2(n_125),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_4),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_4),
.A2(n_59),
.B1(n_63),
.B2(n_161),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_4),
.A2(n_45),
.B1(n_47),
.B2(n_161),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_4),
.A2(n_34),
.B1(n_40),
.B2(n_161),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_5),
.A2(n_59),
.B1(n_63),
.B2(n_69),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_5),
.A2(n_45),
.B1(n_47),
.B2(n_69),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_5),
.A2(n_34),
.B1(n_40),
.B2(n_69),
.Y(n_231)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_7),
.A2(n_44),
.B1(n_59),
.B2(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_7),
.A2(n_44),
.B1(n_65),
.B2(n_66),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_7),
.A2(n_34),
.B1(n_40),
.B2(n_44),
.Y(n_152)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_9),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_9),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_9),
.A2(n_39),
.B1(n_59),
.B2(n_63),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_9),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_10),
.A2(n_59),
.B1(n_63),
.B2(n_71),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_10),
.A2(n_45),
.B1(n_47),
.B2(n_71),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_10),
.A2(n_34),
.B1(n_40),
.B2(n_71),
.Y(n_200)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_11),
.Y(n_341)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_16),
.A2(n_65),
.B1(n_66),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_16),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_16),
.A2(n_59),
.B1(n_63),
.B2(n_176),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_16),
.A2(n_45),
.B1(n_47),
.B2(n_176),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_16),
.A2(n_34),
.B1(n_40),
.B2(n_176),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_21),
.B(n_340),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_17),
.B(n_341),
.Y(n_340)
);

AOI21xp33_ASAP7_75t_L g171 ( 
.A1(n_18),
.A2(n_65),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_18),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_18),
.B(n_198),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_18),
.A2(n_45),
.B1(n_47),
.B2(n_174),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_18),
.A2(n_47),
.B(n_50),
.C(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_18),
.B(n_84),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_18),
.B(n_37),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_18),
.B(n_55),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_18),
.A2(n_63),
.B(n_78),
.C(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_19),
.A2(n_45),
.B1(n_47),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_19),
.A2(n_54),
.B1(n_59),
.B2(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_19),
.A2(n_34),
.B1(n_40),
.B2(n_54),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_19),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_322)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_335),
.B(n_338),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_327),
.B(n_331),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_314),
.B(n_326),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_139),
.B(n_311),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_126),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_101),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_27),
.B(n_101),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_72),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_28),
.B(n_87),
.C(n_99),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_56),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_29),
.A2(n_30),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_41),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_31),
.A2(n_32),
.B1(n_56),
.B2(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_31),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_37),
.B(n_38),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_33),
.A2(n_37),
.B1(n_38),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_33),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_33),
.A2(n_37),
.B1(n_152),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_33),
.A2(n_37),
.B1(n_188),
.B2(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_33),
.A2(n_37),
.B1(n_200),
.B2(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_33),
.A2(n_37),
.B1(n_231),
.B2(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_33),
.A2(n_37),
.B1(n_174),
.B2(n_264),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_33),
.A2(n_37),
.B1(n_257),
.B2(n_264),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_40),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_34),
.B(n_266),
.Y(n_265)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_36),
.A2(n_115),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_36),
.A2(n_150),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_40),
.A2(n_51),
.B(n_174),
.Y(n_245)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_48),
.B1(n_53),
.B2(n_55),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_43),
.A2(n_48),
.B1(n_55),
.B2(n_118),
.Y(n_117)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_47),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

OAI32xp33_ASAP7_75t_L g227 ( 
.A1(n_45),
.A2(n_63),
.A3(n_80),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_47),
.B(n_81),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_53),
.B1(n_55),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_55),
.B(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_48),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_48),
.A2(n_55),
.B1(n_155),
.B2(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_48),
.A2(n_55),
.B1(n_182),
.B2(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_48),
.A2(n_55),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_48),
.A2(n_55),
.B1(n_243),
.B2(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_52),
.A2(n_119),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_52),
.A2(n_156),
.B1(n_223),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_68),
.B2(n_70),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_58),
.B1(n_70),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_57),
.A2(n_58),
.B1(n_68),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_57),
.A2(n_58),
.B1(n_90),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_57),
.A2(n_58),
.B1(n_124),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_57),
.A2(n_58),
.B1(n_171),
.B2(n_175),
.Y(n_170)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_57),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_64),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_58),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_63),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_59),
.A2(n_62),
.A3(n_65),
.B1(n_173),
.B2(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_59),
.B(n_174),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_61),
.B(n_63),
.Y(n_191)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_66),
.B(n_174),
.Y(n_173)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_87),
.B1(n_99),
.B2(n_100),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_74),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_85),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_82),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_83),
.B1(n_84),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_78),
.A2(n_84),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_78),
.A2(n_84),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_78),
.A2(n_84),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_82),
.A2(n_97),
.B1(n_121),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_82),
.A2(n_121),
.B1(n_122),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_82),
.A2(n_121),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_82),
.A2(n_195),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_89),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_93),
.C(n_95),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_89),
.B(n_129),
.C(n_132),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_98),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_93),
.B(n_135),
.C(n_137),
.Y(n_325)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.C(n_109),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_120),
.C(n_123),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_111),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_297)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_123),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_126),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_127),
.B(n_128),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_136),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_138),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_164),
.B(n_310),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_162),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_141),
.B(n_162),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_146),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_142),
.B(n_145),
.Y(n_308)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_146),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_157),
.C(n_159),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_147),
.A2(n_148),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_153),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_157),
.B(n_159),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_305),
.B(n_309),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_215),
.B(n_293),
.C(n_304),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_201),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_167),
.B(n_201),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_185),
.C(n_192),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_168),
.A2(n_169),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_178),
.C(n_184),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_177)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_185),
.B(n_192),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_186),
.B(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.C(n_199),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_193),
.B(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_199),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_198),
.A2(n_212),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_198),
.A2(n_212),
.B1(n_322),
.B2(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_198),
.A2(n_212),
.B(n_329),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_203),
.B(n_204),
.C(n_205),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_214),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_207),
.B(n_210),
.C(n_214),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_292),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_235),
.B(n_291),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_232),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_218),
.B(n_232),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.C(n_224),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_219),
.B(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_221),
.A2(n_224),
.B1(n_225),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_221),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_226),
.A2(n_227),
.B1(n_230),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_228),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_230),
.Y(n_283)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_285),
.B(n_290),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_273),
.B(n_284),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_253),
.B(n_272),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_246),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_239),
.B(n_246),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_241),
.B1(n_244),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_249),
.C(n_251),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_252),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_261),
.B(n_271),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_255),
.B(n_259),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_267),
.B(n_270),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_274),
.B(n_275),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_282),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_280),
.C(n_282),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_295),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_303),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_302),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_302),
.C(n_303),
.Y(n_306)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_316),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_325),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_320),
.B1(n_323),
.B2(n_324),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_323),
.C(n_325),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_328),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_336),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_337),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);


endmodule