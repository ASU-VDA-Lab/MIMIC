module fake_jpeg_7855_n_297 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_34),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_42),
.Y(n_67)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_18),
.B(n_28),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_24),
.B1(n_18),
.B2(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_26),
.B1(n_19),
.B2(n_17),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_18),
.B1(n_21),
.B2(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_29),
.B1(n_19),
.B2(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_61),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_28),
.B(n_20),
.C(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_65),
.Y(n_89)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_35),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_30),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_20),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_68),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_71),
.B(n_87),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_27),
.B(n_22),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_76),
.B(n_88),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_29),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_21),
.B1(n_37),
.B2(n_40),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_90),
.B1(n_95),
.B2(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_81),
.B(n_9),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_23),
.B1(n_19),
.B2(n_26),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_85),
.B1(n_35),
.B2(n_22),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_19),
.B1(n_26),
.B2(n_17),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_29),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_45),
.A2(n_26),
.B1(n_17),
.B2(n_35),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_94),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_0),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_11),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_49),
.A2(n_37),
.B1(n_35),
.B2(n_27),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_49),
.B1(n_59),
.B2(n_46),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_105),
.A2(n_112),
.B1(n_119),
.B2(n_129),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_62),
.B(n_59),
.C(n_64),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_109),
.A2(n_124),
.B(n_101),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_67),
.C(n_52),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_126),
.C(n_72),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_59),
.B1(n_46),
.B2(n_67),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_47),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_125),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_47),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_53),
.B1(n_35),
.B2(n_27),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_22),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_121),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_22),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_0),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_91),
.B(n_86),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_1),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_72),
.B(n_1),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_22),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_127),
.B(n_10),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_1),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_127),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_9),
.B1(n_15),
.B2(n_4),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_132),
.B(n_133),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_80),
.B1(n_99),
.B2(n_92),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_151),
.B1(n_109),
.B2(n_129),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_135),
.B(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_146),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_141),
.B(n_143),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_91),
.B(n_86),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_142),
.A2(n_150),
.B(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_84),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_76),
.C(n_101),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_154),
.C(n_159),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_76),
.B(n_88),
.C(n_71),
.D(n_100),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_152),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_103),
.B(n_100),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_97),
.B1(n_94),
.B2(n_96),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_78),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_153),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_75),
.C(n_70),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_156),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_106),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_158),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_93),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_124),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_171),
.B1(n_134),
.B2(n_147),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_107),
.C(n_119),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_175),
.C(n_182),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_169),
.A2(n_188),
.B(n_143),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_112),
.B1(n_107),
.B2(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_173),
.B(n_176),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_120),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_136),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_124),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_180),
.B(n_187),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_121),
.C(n_124),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_184),
.B(n_186),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_154),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_141),
.B(n_158),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_104),
.B(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_208),
.B1(n_169),
.B2(n_190),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_152),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_116),
.B(n_130),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_142),
.C(n_156),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_199),
.Y(n_221)
);

NAND2x1_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_150),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_198),
.C(n_207),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_148),
.B1(n_157),
.B2(n_160),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_200),
.B1(n_210),
.B2(n_177),
.Y(n_219)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_137),
.B1(n_150),
.B2(n_155),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_146),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_162),
.C(n_170),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_131),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_131),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_97),
.Y(n_206)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_164),
.B1(n_167),
.B2(n_187),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_198),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_141),
.B1(n_105),
.B2(n_116),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_130),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_213),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_178),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_236),
.B1(n_226),
.B2(n_210),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_195),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_163),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_227),
.C(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_188),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_226),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_163),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_172),
.A3(n_175),
.B1(n_168),
.B2(n_182),
.C1(n_162),
.C2(n_165),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_200),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_170),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_231),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_116),
.B(n_8),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_202),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_239),
.B1(n_216),
.B2(n_218),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_193),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_238),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_224),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_248),
.B(n_250),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_251),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_207),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_247),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_208),
.B1(n_197),
.B2(n_201),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_250),
.B1(n_237),
.B2(n_201),
.Y(n_270)
);

NOR2x1_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_223),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_204),
.B(n_230),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_225),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_258),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_227),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_229),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_261),
.B(n_240),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_221),
.C(n_231),
.Y(n_262)
);

NAND4xp25_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_263),
.C(n_6),
.D(n_7),
.Y(n_276)
);

NAND4xp25_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_236),
.C(n_232),
.D(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_232),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_5),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_241),
.A2(n_202),
.B(n_235),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_216),
.B(n_251),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_261),
.C(n_11),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_252),
.B1(n_248),
.B2(n_249),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_271),
.B1(n_258),
.B2(n_256),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_274),
.B(n_253),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_275),
.B(n_276),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_7),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_257),
.B(n_5),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_8),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_5),
.B(n_6),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_6),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_259),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_257),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_266),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_283),
.B1(n_275),
.B2(n_280),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_284),
.C(n_8),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_288),
.C(n_289),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_12),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_266),
.B1(n_12),
.B2(n_13),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_290),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_16),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_292),
.A2(n_293),
.B(n_14),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_16),
.B(n_13),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_291),
.C(n_14),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_294),
.Y(n_297)
);


endmodule