module fake_aes_9758_n_29 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_29);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx2_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
CKINVDCx16_ASAP7_75t_R g9 ( .A(n_5), .Y(n_9) );
NOR2x1p5_ASAP7_75t_L g10 ( .A(n_6), .B(n_3), .Y(n_10) );
OAI22xp5_ASAP7_75t_L g11 ( .A1(n_7), .A2(n_1), .B1(n_6), .B2(n_0), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_2), .B(n_1), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_9), .B(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_12), .B(n_0), .Y(n_15) );
OAI21x1_ASAP7_75t_L g16 ( .A1(n_8), .A2(n_1), .B(n_2), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_12), .B(n_2), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_14), .B(n_8), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_15), .B(n_13), .Y(n_20) );
OAI22xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_11), .B1(n_17), .B2(n_10), .Y(n_21) );
INVxp67_ASAP7_75t_SL g22 ( .A(n_19), .Y(n_22) );
A2O1A1Ixp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_19), .B(n_18), .C(n_10), .Y(n_23) );
OAI21xp33_ASAP7_75t_SL g24 ( .A1(n_22), .A2(n_3), .B(n_4), .Y(n_24) );
NAND3xp33_ASAP7_75t_L g25 ( .A(n_23), .B(n_21), .C(n_4), .Y(n_25) );
NAND2xp5_ASAP7_75t_SL g26 ( .A(n_24), .B(n_14), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_28), .B(n_27), .Y(n_29) );
endmodule