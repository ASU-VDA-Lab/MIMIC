module fake_jpeg_8205_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_55),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_18),
.B1(n_27),
.B2(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_35),
.B1(n_26),
.B2(n_34),
.Y(n_86)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_18),
.B1(n_24),
.B2(n_22),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_40),
.B1(n_21),
.B2(n_26),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_31),
.Y(n_75)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_32),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_30),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_29),
.Y(n_122)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_75),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_82),
.B1(n_86),
.B2(n_89),
.Y(n_109)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_78),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_40),
.B1(n_18),
.B2(n_44),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_62),
.B1(n_68),
.B2(n_20),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_85),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_21),
.B1(n_26),
.B2(n_34),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_35),
.B1(n_31),
.B2(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_49),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_92)
);

OAI22x1_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_15),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_16),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_59),
.B1(n_66),
.B2(n_65),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_108),
.B1(n_115),
.B2(n_78),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_119),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_39),
.B1(n_48),
.B2(n_37),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_113),
.A2(n_51),
.B1(n_67),
.B2(n_54),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_48),
.B1(n_19),
.B2(n_33),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_121),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

NAND2xp67_ASAP7_75t_SL g120 ( 
.A(n_70),
.B(n_36),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_124),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_76),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_128),
.B(n_77),
.Y(n_130)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_127),
.Y(n_148)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_132),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_130),
.A2(n_111),
.B1(n_25),
.B2(n_23),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_77),
.B(n_73),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_151),
.B(n_105),
.Y(n_173)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_72),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_136),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_139),
.B1(n_154),
.B2(n_155),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_72),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_82),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_138),
.C(n_113),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_30),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_85),
.B1(n_96),
.B2(n_80),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_140),
.B(n_144),
.Y(n_163)
);

CKINVDCx12_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_75),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_149),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_0),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_30),
.B(n_32),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_81),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_110),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_32),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_125),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_109),
.A2(n_96),
.B1(n_80),
.B2(n_88),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_99),
.A2(n_88),
.B1(n_33),
.B2(n_28),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_112),
.B1(n_103),
.B2(n_117),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_114),
.B(n_118),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_157),
.A2(n_147),
.B(n_143),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_106),
.B1(n_128),
.B2(n_114),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_158),
.A2(n_170),
.B1(n_185),
.B2(n_142),
.Y(n_193)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_160),
.B(n_167),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_124),
.B(n_118),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_173),
.B(n_177),
.Y(n_199)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_171),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_115),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_181),
.C(n_187),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_174),
.B1(n_183),
.B2(n_132),
.Y(n_210)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_138),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_101),
.B1(n_113),
.B2(n_103),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_110),
.B1(n_105),
.B2(n_127),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_179),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_25),
.A3(n_23),
.B1(n_148),
.B2(n_134),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_83),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_111),
.Y(n_182)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_144),
.A2(n_33),
.B1(n_30),
.B2(n_98),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_156),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_98),
.B1(n_25),
.B2(n_23),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_0),
.Y(n_186)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_98),
.C(n_30),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_194),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_191),
.C(n_196),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_130),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_158),
.B1(n_170),
.B2(n_180),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_159),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_154),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_203),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_161),
.A2(n_147),
.B(n_146),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_205),
.B(n_207),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_152),
.B(n_147),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_213),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_210),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_171),
.B(n_140),
.Y(n_211)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_212),
.B(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_139),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_134),
.C(n_16),
.Y(n_238)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_0),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_177),
.B1(n_162),
.B2(n_148),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_218),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_231),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_165),
.B1(n_166),
.B2(n_163),
.Y(n_225)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_165),
.B1(n_185),
.B2(n_160),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_227),
.B1(n_230),
.B2(n_234),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_186),
.B(n_167),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_200),
.B1(n_192),
.B2(n_195),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_187),
.B1(n_172),
.B2(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_242),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_236),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_244),
.C(n_196),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_189),
.B(n_206),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_243),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_16),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_14),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_245),
.B(n_266),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_215),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_253),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_199),
.C(n_201),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_254),
.C(n_260),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_190),
.Y(n_252)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_199),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_238),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

XOR2x2_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_232),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_257),
.B(n_227),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_193),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_261),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_192),
.C(n_195),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_230),
.C(n_221),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_11),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_264),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_231),
.B(n_10),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_268),
.A2(n_263),
.B1(n_256),
.B2(n_253),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_265),
.A2(n_225),
.B1(n_229),
.B2(n_226),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_263),
.B1(n_245),
.B2(n_258),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_277),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_279),
.C(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_233),
.C(n_237),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_248),
.A2(n_233),
.B1(n_228),
.B2(n_237),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_281),
.B(n_282),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_257),
.A2(n_219),
.B1(n_220),
.B2(n_217),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_239),
.B(n_10),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_9),
.B(n_8),
.Y(n_292)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_288),
.C(n_291),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_249),
.Y(n_288)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_251),
.C(n_254),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_298),
.B(n_284),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_251),
.C(n_263),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_299),
.C(n_273),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_8),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_296),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_7),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_1),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_283),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_1),
.B(n_2),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_1),
.C(n_2),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_301),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_288),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_303),
.B(n_305),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_281),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_310),
.C(n_299),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_275),
.B1(n_282),
.B2(n_268),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_269),
.C(n_277),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_287),
.A2(n_278),
.B(n_270),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_312),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_285),
.A2(n_267),
.B1(n_3),
.B2(n_4),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_293),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_315),
.C(n_317),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_291),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_322),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_302),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_267),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_3),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_308),
.Y(n_323)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_323),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_307),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_328),
.B(n_329),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_304),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_325),
.A2(n_321),
.B(n_314),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_332),
.C(n_327),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_315),
.C(n_4),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_333),
.A2(n_323),
.B(n_326),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_335),
.B(n_331),
.C(n_6),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_3),
.C(n_5),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_5),
.B(n_7),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_5),
.Y(n_340)
);


endmodule