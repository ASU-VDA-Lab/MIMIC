module fake_aes_11586_n_562 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_562);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_562;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_73;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g70 ( .A(n_48), .Y(n_70) );
INVx2_ASAP7_75t_L g71 ( .A(n_58), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_64), .Y(n_72) );
INVxp33_ASAP7_75t_SL g73 ( .A(n_53), .Y(n_73) );
BUFx2_ASAP7_75t_L g74 ( .A(n_27), .Y(n_74) );
CKINVDCx5p33_ASAP7_75t_R g75 ( .A(n_29), .Y(n_75) );
INVxp67_ASAP7_75t_SL g76 ( .A(n_6), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_33), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_38), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_43), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_67), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_26), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_5), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_3), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_60), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_49), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_68), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_65), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_36), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_5), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_3), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_59), .Y(n_91) );
CKINVDCx14_ASAP7_75t_R g92 ( .A(n_56), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_20), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_31), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_52), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_69), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_19), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_57), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_22), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_55), .Y(n_100) );
HB1xp67_ASAP7_75t_L g101 ( .A(n_8), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_7), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_21), .B(n_46), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_32), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_25), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_12), .Y(n_106) );
NOR2xp67_ASAP7_75t_L g107 ( .A(n_34), .B(n_37), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_12), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_63), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_16), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_50), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_74), .B(n_0), .Y(n_114) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_72), .A2(n_23), .B(n_62), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_93), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_91), .Y(n_117) );
INVx3_ASAP7_75t_L g118 ( .A(n_91), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_91), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_105), .B(n_0), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_80), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_93), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_84), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_79), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_105), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_87), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_82), .B(n_1), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_101), .Y(n_133) );
INVx5_ASAP7_75t_L g134 ( .A(n_96), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_89), .B(n_1), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_88), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_96), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_94), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_94), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_95), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_79), .B(n_2), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_90), .B(n_102), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_70), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_70), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_116), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_132), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_119), .B(n_92), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_128), .B(n_108), .Y(n_153) );
INVx2_ASAP7_75t_SL g154 ( .A(n_119), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_138), .B(n_99), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_138), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_117), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_138), .B(n_99), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_129), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_117), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_147), .B(n_90), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_138), .Y(n_163) );
NAND2x1p5_ASAP7_75t_L g164 ( .A(n_114), .B(n_112), .Y(n_164) );
AND3x4_ASAP7_75t_L g165 ( .A(n_147), .B(n_127), .C(n_107), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_147), .Y(n_166) );
NAND3xp33_ASAP7_75t_L g167 ( .A(n_128), .B(n_102), .C(n_111), .Y(n_167) );
BUFx4f_ASAP7_75t_L g168 ( .A(n_147), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_133), .B(n_75), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_123), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
INVx5_ASAP7_75t_L g172 ( .A(n_117), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_114), .B(n_111), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_133), .B(n_85), .Y(n_174) );
INVx4_ASAP7_75t_SL g175 ( .A(n_117), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_129), .Y(n_176) );
NAND2x1p5_ASAP7_75t_L g177 ( .A(n_114), .B(n_112), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_123), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_123), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_137), .B(n_109), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_145), .Y(n_181) );
NAND3x1_ASAP7_75t_L g182 ( .A(n_146), .B(n_106), .C(n_109), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_135), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_118), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_117), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
NAND3xp33_ASAP7_75t_L g187 ( .A(n_135), .B(n_106), .C(n_95), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_118), .Y(n_190) );
INVxp67_ASAP7_75t_SL g191 ( .A(n_137), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_113), .B(n_110), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_113), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_132), .Y(n_194) );
INVx2_ASAP7_75t_SL g195 ( .A(n_134), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_132), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_118), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_122), .B(n_86), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_117), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_122), .B(n_110), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_155), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_183), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_155), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_168), .B(n_124), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_156), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_155), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_168), .B(n_124), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_191), .B(n_126), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_183), .B(n_126), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_173), .B(n_146), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_173), .B(n_146), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_168), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_169), .B(n_125), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_190), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_166), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_180), .B(n_141), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_162), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_180), .B(n_141), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_162), .Y(n_219) );
BUFx8_ASAP7_75t_L g220 ( .A(n_160), .Y(n_220) );
OR2x2_ASAP7_75t_L g221 ( .A(n_160), .B(n_131), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_176), .Y(n_222) );
BUFx8_ASAP7_75t_L g223 ( .A(n_154), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_176), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_156), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_162), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_164), .B(n_140), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_190), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_164), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_164), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_156), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_174), .B(n_125), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_154), .B(n_131), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_190), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_177), .Y(n_235) );
INVx5_ASAP7_75t_L g236 ( .A(n_156), .Y(n_236) );
AND2x6_ASAP7_75t_L g237 ( .A(n_157), .B(n_97), .Y(n_237) );
OAI221xp5_ASAP7_75t_L g238 ( .A1(n_177), .A2(n_136), .B1(n_130), .B2(n_144), .C(n_143), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_156), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_177), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_170), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_153), .A2(n_121), .B(n_130), .C(n_144), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_152), .A2(n_77), .B1(n_143), .B2(n_140), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_152), .B(n_136), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_163), .B(n_134), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_173), .B(n_123), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_192), .B(n_134), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_192), .B(n_134), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_198), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_170), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_192), .B(n_134), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_170), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_184), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_229), .B(n_200), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_215), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_249), .B(n_200), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_221), .B(n_167), .Y(n_257) );
INVx5_ASAP7_75t_L g258 ( .A(n_205), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_209), .B(n_200), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_230), .A2(n_182), .B1(n_165), .B2(n_187), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_209), .B(n_156), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_240), .B(n_178), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_235), .B(n_159), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_201), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_201), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_203), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_220), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_204), .A2(n_186), .B(n_188), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_204), .A2(n_181), .B(n_189), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_203), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_206), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
OAI22xp33_ASAP7_75t_L g273 ( .A1(n_224), .A2(n_179), .B1(n_178), .B2(n_193), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_214), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_207), .A2(n_195), .B(n_197), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_214), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_225), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
AO22x1_ASAP7_75t_L g279 ( .A1(n_223), .A2(n_165), .B1(n_159), .B2(n_73), .Y(n_279) );
BUFx4_ASAP7_75t_SL g280 ( .A(n_222), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_228), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_220), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_234), .Y(n_283) );
AOI21xp33_ASAP7_75t_L g284 ( .A1(n_233), .A2(n_182), .B(n_197), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_238), .A2(n_184), .B1(n_178), .B2(n_179), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_205), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_210), .B(n_179), .Y(n_287) );
BUFx2_ASAP7_75t_SL g288 ( .A(n_225), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_205), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_210), .B(n_150), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_211), .B(n_159), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_234), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_213), .A2(n_150), .B(n_139), .C(n_116), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_255), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_280), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_264), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_256), .B(n_211), .Y(n_297) );
INVx4_ASAP7_75t_L g298 ( .A(n_258), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_293), .B(n_223), .C(n_243), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_255), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_260), .A2(n_222), .B1(n_202), .B2(n_159), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_265), .Y(n_302) );
OAI211xp5_ASAP7_75t_L g303 ( .A1(n_284), .A2(n_242), .B(n_232), .C(n_213), .Y(n_303) );
OAI22xp33_ASAP7_75t_L g304 ( .A1(n_267), .A2(n_227), .B1(n_216), .B2(n_218), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_SL g305 ( .A1(n_261), .A2(n_247), .B(n_248), .C(n_251), .Y(n_305) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_267), .A2(n_231), .B1(n_205), .B2(n_239), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_257), .B(n_244), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_257), .B(n_212), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_282), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_290), .B(n_208), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_254), .A2(n_159), .B1(n_237), .B2(n_217), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_259), .A2(n_219), .B1(n_226), .B2(n_239), .Y(n_313) );
CKINVDCx8_ASAP7_75t_R g314 ( .A(n_288), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_290), .B(n_246), .Y(n_315) );
OR2x6_ASAP7_75t_L g316 ( .A(n_288), .B(n_231), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_258), .Y(n_317) );
NOR2xp67_ASAP7_75t_L g318 ( .A(n_258), .B(n_236), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_254), .A2(n_159), .B1(n_237), .B2(n_212), .Y(n_319) );
OAI22xp5_ASAP7_75t_SL g320 ( .A1(n_295), .A2(n_279), .B1(n_291), .B2(n_76), .Y(n_320) );
AOI22xp33_ASAP7_75t_SL g321 ( .A1(n_299), .A2(n_254), .B1(n_237), .B2(n_279), .Y(n_321) );
OAI22xp33_ASAP7_75t_L g322 ( .A1(n_304), .A2(n_273), .B1(n_239), .B2(n_231), .Y(n_322) );
CKINVDCx16_ASAP7_75t_R g323 ( .A(n_309), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_301), .A2(n_237), .B1(n_232), .B2(n_287), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_307), .B(n_208), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_305), .A2(n_269), .B(n_268), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_294), .B(n_263), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_307), .A2(n_237), .B1(n_148), .B2(n_274), .Y(n_328) );
AOI222xp33_ASAP7_75t_L g329 ( .A1(n_310), .A2(n_262), .B1(n_207), .B2(n_251), .C1(n_285), .C2(n_272), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_311), .B(n_287), .Y(n_330) );
NAND2x1_ASAP7_75t_L g331 ( .A(n_298), .B(n_286), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_315), .B(n_262), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_308), .A2(n_263), .B1(n_241), .B2(n_252), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_297), .A2(n_292), .B1(n_266), .B2(n_281), .C(n_265), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_303), .A2(n_292), .B1(n_281), .B2(n_266), .C(n_272), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_294), .Y(n_336) );
AOI21xp33_ASAP7_75t_SL g337 ( .A1(n_300), .A2(n_115), .B(n_4), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_300), .B(n_263), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_314), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_315), .A2(n_274), .B1(n_148), .B2(n_250), .C(n_116), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_302), .B(n_264), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_302), .A2(n_148), .B1(n_142), .B2(n_139), .C(n_245), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_296), .B(n_270), .Y(n_343) );
AOI31xp33_ASAP7_75t_SL g344 ( .A1(n_329), .A2(n_103), .A3(n_78), .B(n_81), .Y(n_344) );
CKINVDCx14_ASAP7_75t_R g345 ( .A(n_339), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_320), .A2(n_313), .B1(n_312), .B2(n_319), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_324), .A2(n_275), .B(n_306), .Y(n_347) );
OAI222xp33_ASAP7_75t_L g348 ( .A1(n_321), .A2(n_314), .B1(n_316), .B2(n_298), .C1(n_97), .C2(n_104), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_325), .B(n_296), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_336), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_341), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_321), .A2(n_317), .B1(n_298), .B2(n_316), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g353 ( .A1(n_328), .A2(n_142), .B1(n_139), .B2(n_107), .C(n_104), .Y(n_353) );
OAI221xp5_ASAP7_75t_L g354 ( .A1(n_328), .A2(n_142), .B1(n_98), .B2(n_100), .C(n_245), .Y(n_354) );
OAI221xp5_ASAP7_75t_L g355 ( .A1(n_330), .A2(n_100), .B1(n_98), .B2(n_317), .C(n_316), .Y(n_355) );
OR2x6_ASAP7_75t_L g356 ( .A(n_331), .B(n_316), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_332), .B(n_323), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_343), .Y(n_358) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_322), .A2(n_81), .B1(n_78), .B2(n_71), .C1(n_134), .C2(n_132), .Y(n_359) );
OAI31xp33_ASAP7_75t_L g360 ( .A1(n_322), .A2(n_71), .A3(n_276), .B(n_270), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_327), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_333), .A2(n_271), .B1(n_283), .B2(n_278), .C(n_276), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_327), .B(n_271), .Y(n_363) );
OA21x2_ASAP7_75t_L g364 ( .A1(n_326), .A2(n_199), .B(n_158), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_338), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_338), .B(n_278), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_334), .B(n_115), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_335), .Y(n_368) );
OAI211xp5_ASAP7_75t_SL g369 ( .A1(n_342), .A2(n_158), .B(n_161), .C(n_185), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_337), .B(n_283), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_340), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_336), .Y(n_372) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_321), .B(n_149), .C(n_132), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_336), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_336), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_356), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_363), .Y(n_377) );
NAND2xp67_ASAP7_75t_L g378 ( .A(n_372), .B(n_2), .Y(n_378) );
NOR3xp33_ASAP7_75t_L g379 ( .A(n_355), .B(n_199), .C(n_185), .Y(n_379) );
AOI322xp5_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_132), .A3(n_149), .B1(n_134), .B2(n_8), .C1(n_9), .C2(n_10), .Y(n_380) );
AOI211xp5_ASAP7_75t_L g381 ( .A1(n_344), .A2(n_149), .B(n_117), .C(n_120), .Y(n_381) );
AOI33xp33_ASAP7_75t_L g382 ( .A1(n_374), .A2(n_4), .A3(n_6), .B1(n_7), .B2(n_9), .B3(n_10), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_351), .B(n_149), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_350), .B(n_115), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_350), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_372), .B(n_115), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_351), .B(n_149), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_370), .A2(n_318), .B(n_115), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_375), .B(n_149), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_375), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_358), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_353), .A2(n_149), .B1(n_120), .B2(n_151), .C(n_171), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_358), .Y(n_393) );
AO22x1_ASAP7_75t_L g394 ( .A1(n_365), .A2(n_258), .B1(n_277), .B2(n_289), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_359), .B(n_120), .C(n_151), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_356), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_361), .B(n_11), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_357), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_360), .A2(n_286), .B(n_231), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_368), .A2(n_120), .B1(n_318), .B2(n_286), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_357), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_349), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_364), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_373), .A2(n_286), .B(n_239), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_364), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_371), .A2(n_258), .B1(n_289), .B2(n_286), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_368), .A2(n_346), .B1(n_345), .B2(n_352), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_370), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_356), .B(n_47), .Y(n_411) );
AND2x2_ASAP7_75t_SL g412 ( .A(n_348), .B(n_277), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_366), .B(n_11), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_366), .B(n_13), .Y(n_414) );
NOR3xp33_ASAP7_75t_L g415 ( .A(n_354), .B(n_161), .C(n_277), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_356), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_367), .A2(n_120), .B1(n_196), .B2(n_151), .C(n_194), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_367), .A2(n_120), .B1(n_236), .B2(n_195), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_362), .Y(n_419) );
OAI31xp33_ASAP7_75t_SL g420 ( .A1(n_347), .A2(n_13), .A3(n_14), .B(n_15), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_369), .A2(n_120), .B1(n_196), .B2(n_194), .C(n_171), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_390), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_385), .Y(n_423) );
AND2x2_ASAP7_75t_SL g424 ( .A(n_376), .B(n_15), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_402), .B(n_16), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_390), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_385), .B(n_17), .Y(n_427) );
NAND5xp2_ASAP7_75t_L g428 ( .A(n_420), .B(n_17), .C(n_18), .D(n_24), .E(n_28), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_391), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_405), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_411), .B(n_236), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_405), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_410), .B(n_196), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_393), .Y(n_434) );
OAI31xp33_ASAP7_75t_L g435 ( .A1(n_409), .A2(n_253), .A3(n_35), .B(n_39), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_398), .B(n_196), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_404), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_401), .B(n_196), .Y(n_438) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_411), .B(n_236), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_403), .B(n_30), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_416), .B(n_194), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_377), .B(n_194), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_416), .B(n_40), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_404), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_396), .B(n_171), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_378), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_407), .B(n_151), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_411), .B(n_41), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_413), .B(n_151), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_397), .B(n_172), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_383), .B(n_42), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_384), .B(n_44), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_384), .B(n_45), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_389), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_387), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_386), .B(n_51), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_386), .B(n_54), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_412), .A2(n_253), .B1(n_172), .B2(n_175), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_388), .B(n_61), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_397), .B(n_419), .Y(n_461) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_414), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_395), .B(n_66), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_382), .B(n_172), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_382), .B(n_172), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_412), .A2(n_172), .B1(n_175), .B2(n_381), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_417), .B(n_175), .Y(n_467) );
NAND4xp25_ASAP7_75t_L g468 ( .A(n_380), .B(n_175), .C(n_379), .D(n_400), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_394), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_461), .B(n_394), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_423), .B(n_378), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_462), .B(n_461), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_429), .B(n_408), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_449), .B(n_399), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_434), .B(n_418), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_422), .B(n_406), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_437), .B(n_392), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_437), .B(n_421), .Y(n_478) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_424), .B(n_415), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_426), .B(n_438), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_424), .B(n_469), .Y(n_481) );
NAND4xp25_ASAP7_75t_L g482 ( .A(n_428), .B(n_435), .C(n_468), .D(n_446), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_444), .B(n_447), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_426), .B(n_438), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_447), .B(n_455), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_455), .B(n_456), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_433), .B(n_427), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_456), .B(n_433), .Y(n_488) );
INVx3_ASAP7_75t_SL g489 ( .A(n_449), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_427), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_430), .B(n_432), .Y(n_491) );
NOR2xp67_ASAP7_75t_SL g492 ( .A(n_431), .B(n_453), .Y(n_492) );
XOR2x2_ASAP7_75t_L g493 ( .A(n_439), .B(n_449), .Y(n_493) );
XNOR2xp5_ASAP7_75t_L g494 ( .A(n_439), .B(n_425), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_436), .Y(n_495) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_442), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_445), .B(n_443), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_448), .B(n_445), .Y(n_498) );
NAND4xp25_ASAP7_75t_SL g499 ( .A(n_466), .B(n_459), .C(n_465), .D(n_464), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_453), .B(n_454), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_439), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_441), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_472), .B(n_458), .Y(n_503) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_481), .A2(n_441), .B(n_450), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_479), .A2(n_482), .B1(n_499), .B2(n_470), .Y(n_505) );
NOR3xp33_ASAP7_75t_L g506 ( .A(n_471), .B(n_465), .C(n_440), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_489), .B(n_463), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_492), .A2(n_463), .B1(n_460), .B2(n_451), .Y(n_508) );
XNOR2xp5_ASAP7_75t_L g509 ( .A(n_493), .B(n_457), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_485), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_487), .B(n_460), .Y(n_511) );
XNOR2x2_ASAP7_75t_L g512 ( .A(n_494), .B(n_452), .Y(n_512) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_501), .B(n_463), .Y(n_513) );
XOR2x2_ASAP7_75t_L g514 ( .A(n_500), .B(n_460), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_485), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_486), .B(n_452), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_486), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_471), .A2(n_467), .B(n_496), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_477), .B(n_475), .C(n_478), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_478), .A2(n_477), .B(n_475), .Y(n_520) );
OAI21xp5_ASAP7_75t_SL g521 ( .A1(n_500), .A2(n_497), .B(n_474), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_498), .A2(n_474), .B1(n_488), .B2(n_502), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_480), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_491), .A2(n_495), .B(n_484), .Y(n_524) );
XNOR2xp5_ASAP7_75t_L g525 ( .A(n_473), .B(n_491), .Y(n_525) );
XOR2x2_ASAP7_75t_L g526 ( .A(n_476), .B(n_424), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_489), .Y(n_527) );
AOI21xp33_ASAP7_75t_SL g528 ( .A1(n_489), .A2(n_481), .B(n_479), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_483), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_472), .B(n_490), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_489), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_479), .A2(n_424), .B(n_481), .C(n_492), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_483), .Y(n_533) );
OAI21xp33_ASAP7_75t_SL g534 ( .A1(n_481), .A2(n_469), .B(n_472), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_515), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_529), .Y(n_536) );
BUFx2_ASAP7_75t_R g537 ( .A(n_509), .Y(n_537) );
OAI211xp5_ASAP7_75t_L g538 ( .A1(n_505), .A2(n_528), .B(n_532), .C(n_534), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_531), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_510), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_533), .Y(n_541) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_532), .A2(n_519), .B(n_520), .C(n_527), .Y(n_542) );
OAI321xp33_ASAP7_75t_L g543 ( .A1(n_507), .A2(n_513), .A3(n_518), .B1(n_512), .B2(n_508), .C(n_516), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g544 ( .A1(n_519), .A2(n_521), .B1(n_522), .B2(n_526), .C(n_506), .Y(n_544) );
INVxp33_ASAP7_75t_SL g545 ( .A(n_506), .Y(n_545) );
XNOR2x1_ASAP7_75t_L g546 ( .A(n_539), .B(n_526), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_535), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_540), .Y(n_548) );
AOI211xp5_ASAP7_75t_SL g549 ( .A1(n_538), .A2(n_516), .B(n_524), .C(n_503), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_544), .A2(n_522), .B1(n_525), .B2(n_507), .Y(n_550) );
NAND4xp75_ASAP7_75t_L g551 ( .A(n_537), .B(n_504), .C(n_511), .D(n_530), .Y(n_551) );
AOI211x1_ASAP7_75t_L g552 ( .A1(n_550), .A2(n_542), .B(n_545), .C(n_543), .Y(n_552) );
OAI222xp33_ASAP7_75t_L g553 ( .A1(n_549), .A2(n_545), .B1(n_513), .B2(n_523), .C1(n_541), .C2(n_536), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_546), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_554), .A2(n_551), .B1(n_548), .B2(n_547), .Y(n_555) );
XNOR2x1_ASAP7_75t_L g556 ( .A(n_552), .B(n_549), .Y(n_556) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_555), .A2(n_553), .B(n_536), .Y(n_557) );
OR2x2_ASAP7_75t_SL g558 ( .A(n_556), .B(n_504), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_558), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_559), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_560), .A2(n_557), .B(n_514), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_561), .A2(n_557), .B(n_517), .Y(n_562) );
endmodule