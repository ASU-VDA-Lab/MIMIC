module fake_netlist_1_7944_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_4), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_2), .Y(n_15) );
O2A1O1Ixp33_ASAP7_75t_L g16 ( .A1(n_14), .A2(n_0), .B(n_1), .C(n_2), .Y(n_16) );
OAI22xp5_ASAP7_75t_L g17 ( .A1(n_14), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_11), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_11), .A2(n_5), .B(n_6), .Y(n_19) );
NAND2x1_ASAP7_75t_L g20 ( .A(n_11), .B(n_13), .Y(n_20) );
NOR3xp33_ASAP7_75t_SL g21 ( .A(n_17), .B(n_15), .C(n_12), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_18), .A2(n_13), .B1(n_15), .B2(n_10), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_20), .Y(n_24) );
INVx3_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_23), .B(n_19), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
AOI321xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_16), .A3(n_24), .B1(n_26), .B2(n_21), .C(n_25), .Y(n_28) );
BUFx6f_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
INVx1_ASAP7_75t_SL g30 ( .A(n_28), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
AOI22xp33_ASAP7_75t_R g33 ( .A1(n_31), .A2(n_7), .B1(n_8), .B2(n_32), .Y(n_33) );
endmodule