module fake_jpeg_1266_n_187 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_1),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_13),
.B(n_9),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_31),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_31),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_32),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_68),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_78),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_33),
.A2(n_21),
.B1(n_19),
.B2(n_26),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_21),
.B1(n_25),
.B2(n_17),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_30),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_34),
.B(n_13),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_16),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_37),
.C(n_38),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_63),
.C(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_44),
.B1(n_43),
.B2(n_48),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_68),
.B1(n_57),
.B2(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_53),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_82),
.Y(n_124)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_103),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_84),
.B1(n_85),
.B2(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_106),
.Y(n_114)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_60),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_70),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_9),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_7),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_111),
.B1(n_121),
.B2(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_77),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_125),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_93),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_61),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_102),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_54),
.B1(n_69),
.B2(n_71),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_82),
.B1(n_72),
.B2(n_5),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_3),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_3),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_100),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_4),
.C(n_5),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_93),
.C(n_89),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_137),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_103),
.B(n_109),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_139),
.B(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_87),
.B1(n_95),
.B2(n_90),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_123),
.B1(n_128),
.B2(n_127),
.Y(n_150)
);

HAxp5_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_109),
.CON(n_136),
.SN(n_136)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_94),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_144),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_99),
.B(n_101),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_92),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_143),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_111),
.B1(n_110),
.B2(n_121),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_150),
.B1(n_145),
.B2(n_140),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_117),
.B(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_153),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_128),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_129),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_132),
.B1(n_142),
.B2(n_136),
.Y(n_162)
);

AOI321xp33_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_132),
.A3(n_130),
.B1(n_143),
.B2(n_138),
.C(n_133),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_164),
.B(n_165),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_151),
.B1(n_153),
.B2(n_148),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_168),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_147),
.B(n_130),
.C(n_152),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_152),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_161),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_164),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_175),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_160),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_174),
.A2(n_6),
.B1(n_86),
.B2(n_176),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_171),
.B(n_128),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_177),
.A2(n_171),
.B(n_112),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_179),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_176),
.A2(n_107),
.B1(n_98),
.B2(n_6),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_86),
.C(n_174),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_179),
.B(n_117),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_183),
.A2(n_181),
.B(n_180),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_186),
.B(n_185),
.CI(n_167),
.CON(n_187),
.SN(n_187)
);


endmodule