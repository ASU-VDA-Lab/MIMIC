module real_jpeg_31379_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_710, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_710;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_704;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_707;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_703;
wire n_110;
wire n_195;
wire n_533;
wire n_592;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_431;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_699;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_708;
wire n_196;
wire n_375;
wire n_667;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_702;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_706;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_705;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_641;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_0),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_0),
.Y(n_227)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_0),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_0),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_0),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_1),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_1),
.A2(n_75),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_1),
.A2(n_75),
.B1(n_238),
.B2(n_242),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_1),
.A2(n_75),
.B1(n_341),
.B2(n_345),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_2),
.A2(n_359),
.B1(n_360),
.B2(n_361),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_2),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_2),
.A2(n_47),
.B1(n_359),
.B2(n_462),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_2),
.A2(n_359),
.B1(n_561),
.B2(n_562),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_2),
.A2(n_359),
.B1(n_641),
.B2(n_645),
.Y(n_640)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_3),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_3),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_4),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_4),
.A2(n_51),
.B1(n_193),
.B2(n_199),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_4),
.A2(n_51),
.B1(n_149),
.B2(n_238),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_4),
.A2(n_51),
.B1(n_293),
.B2(n_296),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_5),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_5),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_5),
.A2(n_121),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_5),
.A2(n_121),
.B1(n_348),
.B2(n_351),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_5),
.A2(n_121),
.B1(n_478),
.B2(n_480),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_6),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_6),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_6),
.A2(n_158),
.B1(n_170),
.B2(n_175),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_6),
.A2(n_158),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_6),
.A2(n_158),
.B1(n_695),
.B2(n_698),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_7),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_7),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_7),
.A2(n_252),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_7),
.A2(n_252),
.B1(n_446),
.B2(n_450),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_7),
.A2(n_252),
.B1(n_540),
.B2(n_543),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_8),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_8),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_8),
.A2(n_311),
.B1(n_386),
.B2(n_389),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g506 ( 
.A1(n_8),
.A2(n_311),
.B1(n_507),
.B2(n_511),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_8),
.A2(n_311),
.B1(n_604),
.B2(n_618),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_84),
.B1(n_89),
.B2(n_90),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_9),
.A2(n_89),
.B1(n_262),
.B2(n_267),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_9),
.A2(n_89),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_9),
.A2(n_89),
.B1(n_420),
.B2(n_422),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_10),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_13),
.Y(n_137)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_13),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_13),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_13),
.Y(n_298)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_14),
.Y(n_142)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_14),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_15),
.B(n_703),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_15),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_16),
.B(n_92),
.Y(n_406)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_16),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_16),
.B(n_97),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_16),
.B(n_532),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_16),
.A2(n_457),
.B1(n_569),
.B2(n_574),
.Y(n_568)
);

OAI21xp33_ASAP7_75t_L g658 ( 
.A1(n_16),
.A2(n_219),
.B(n_621),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_17),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_17),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_18),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_18),
.Y(n_266)
);

OAI311xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_687),
.A3(n_702),
.B1(n_704),
.C1(n_707),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_20),
.B(n_708),
.Y(n_707)
);

OAI21x1_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_203),
.B(n_685),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_185),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_23),
.B(n_185),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_163),
.C(n_164),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_25),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_25),
.B(n_208),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_81),
.C(n_127),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_27),
.A2(n_127),
.B1(n_167),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_27),
.Y(n_214)
);

AO22x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_45),
.B1(n_60),
.B2(n_72),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_28),
.A2(n_45),
.B1(n_60),
.B2(n_169),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_SL g189 ( 
.A1(n_28),
.A2(n_60),
.B(n_169),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_28),
.A2(n_72),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_28),
.A2(n_60),
.B1(n_261),
.B2(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_28),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_28),
.B(n_368),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_28),
.A2(n_60),
.B1(n_460),
.B2(n_461),
.Y(n_459)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_61),
.Y(n_60)
);

AOI22x1_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_34),
.B1(n_37),
.B2(n_41),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_30),
.A2(n_146),
.B1(n_149),
.B2(n_152),
.Y(n_145)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_32),
.Y(n_350)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_33),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_33),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_33),
.Y(n_587)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_39),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_40),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_40),
.Y(n_354)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_44),
.Y(n_529)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_48),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_49),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_49),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_50),
.Y(n_174)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_50),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_50),
.Y(n_577)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_58),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_59),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_60),
.Y(n_260)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_60),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_60),
.B(n_368),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_63),
.Y(n_525)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_80),
.Y(n_369)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_81),
.B(n_165),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_82),
.B(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_96),
.B1(n_108),
.B2(n_120),
.Y(n_82)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_83),
.Y(n_178)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_111),
.B1(n_114),
.B2(n_116),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_95),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_95),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_95),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_95),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_95),
.Y(n_697)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_96),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_96),
.A2(n_108),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g693 ( 
.A1(n_96),
.A2(n_108),
.B1(n_192),
.B2(n_694),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_97),
.B(n_120),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_97),
.B(n_250),
.Y(n_316)
);

AO22x1_ASAP7_75t_SL g357 ( 
.A1(n_97),
.A2(n_109),
.B1(n_310),
.B2(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_97),
.B(n_358),
.Y(n_395)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_104),
.B2(n_106),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_103),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g391 ( 
.A(n_105),
.Y(n_391)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_109),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_109),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_109),
.B(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_113),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_113),
.Y(n_413)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_126),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_167),
.B1(n_168),
.B2(n_176),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_143),
.B(n_155),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_128),
.A2(n_143),
.B1(n_155),
.B2(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_128),
.A2(n_143),
.B1(n_445),
.B2(n_453),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_128),
.B(n_445),
.Y(n_514)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_144),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_129),
.Y(n_628)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_130),
.B(n_145),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_135),
.B1(n_138),
.B2(n_140),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_131),
.A2(n_135),
.B1(n_138),
.B2(n_140),
.Y(n_247)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g592 ( 
.A(n_133),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_136),
.Y(n_295)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_136),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_137),
.Y(n_421)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_137),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_137),
.Y(n_547)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_139),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_141),
.Y(n_611)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_143),
.B(n_614),
.Y(n_613)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_143),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_151),
.Y(n_565)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_156),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx5_ASAP7_75t_L g452 ( 
.A(n_157),
.Y(n_452)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_157),
.Y(n_513)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_162),
.Y(n_449)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_162),
.Y(n_602)
);

INVxp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_177),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_176),
.C(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_170),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_174),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_184),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g691 ( 
.A(n_186),
.B(n_190),
.C(n_201),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_201),
.B2(n_202),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_193),
.A2(n_457),
.B(n_458),
.Y(n_456)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_198),
.Y(n_401)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21x1_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_321),
.B(n_679),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_268),
.Y(n_205)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_206),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_209),
.B(n_210),
.Y(n_206)
);

NOR3xp33_ASAP7_75t_L g684 ( 
.A(n_207),
.B(n_209),
.C(n_210),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.C(n_256),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_212),
.A2(n_256),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_212),
.Y(n_319)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_216),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_248),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_SL g332 ( 
.A1(n_217),
.A2(n_218),
.B(n_234),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_234),
.Y(n_217)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

AOI21x1_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_225),
.B(n_228),
.Y(n_218)
);

OAI22x1_ASAP7_75t_SL g291 ( 
.A1(n_219),
.A2(n_228),
.B1(n_292),
.B2(n_299),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_219),
.A2(n_419),
.B1(n_477),
.B2(n_483),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_219),
.A2(n_617),
.B(n_621),
.Y(n_616)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_220),
.B(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_220),
.A2(n_340),
.B1(n_415),
.B2(n_418),
.Y(n_414)
);

AO22x1_ASAP7_75t_SL g538 ( 
.A1(n_220),
.A2(n_539),
.B1(n_548),
.B2(n_549),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_220),
.A2(n_636),
.B1(n_638),
.B2(n_639),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_R g656 ( 
.A(n_220),
.B(n_539),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_222),
.Y(n_338)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx4f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_231),
.Y(n_620)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_233),
.Y(n_344)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_233),
.Y(n_479)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_233),
.Y(n_597)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_233),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_245),
.B2(n_246),
.Y(n_235)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_236),
.A2(n_237),
.B1(n_246),
.B2(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_236),
.A2(n_246),
.B1(n_286),
.B2(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_236),
.A2(n_246),
.B1(n_506),
.B2(n_560),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_237),
.Y(n_274)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_241),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_258),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_255),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_249),
.B(n_395),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_251),
.Y(n_360)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_259),
.Y(n_280)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_317),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_L g681 ( 
.A(n_269),
.B(n_317),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_279),
.C(n_281),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_271),
.B(n_280),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_278),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_276),
.B(n_277),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_275),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_282),
.B(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_302),
.C(n_307),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_291),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_285),
.B(n_291),
.Y(n_424)
);

BUFx4f_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_292),
.A2(n_337),
.B(n_339),
.Y(n_336)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_298),
.Y(n_542)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_298),
.Y(n_609)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_299),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_301),
.Y(n_655)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_308),
.Y(n_330)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_304),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

INVx11_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx12f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_316),
.B(n_455),
.Y(n_454)
);

NAND2x1_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_494),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_433),
.B(n_490),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_324),
.B(n_676),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_376),
.B(n_379),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_325),
.B(n_376),
.Y(n_493)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_326),
.B(n_377),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.C(n_333),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_328),
.A2(n_329),
.B1(n_332),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_332),
.Y(n_432)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_334),
.B(n_431),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_355),
.B(n_375),
.Y(n_334)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_346),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_336),
.B(n_346),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_338),
.Y(n_622)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_347),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_354),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_364),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_364),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_356),
.A2(n_357),
.B1(n_365),
.B2(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

OAI22x1_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_373),
.B2(n_374),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_366),
.A2(n_385),
.B(n_392),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_366),
.A2(n_392),
.B(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_374),
.A2(n_474),
.B(n_475),
.Y(n_473)
);

NOR2x1_ASAP7_75t_R g624 ( 
.A(n_374),
.B(n_457),
.Y(n_624)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_430),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_380),
.B(n_430),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_424),
.C(n_425),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_381),
.B(n_436),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_393),
.C(n_396),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_383),
.A2(n_384),
.B1(n_393),
.B2(n_394),
.Y(n_442)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_385),
.Y(n_460)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_442),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_414),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_398),
.B(n_414),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_402),
.B1(n_406),
.B2(n_407),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_406),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_417),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_417),
.Y(n_664)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_424),
.A2(n_426),
.B1(n_437),
.B2(n_438),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_424),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_426),
.Y(n_437)
);

XNOR2x1_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_439),
.C(n_466),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_435),
.A2(n_677),
.B(n_678),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_439),
.Y(n_677)
);

MAJx2_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_443),
.C(n_464),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_440),
.A2(n_441),
.B1(n_488),
.B2(n_489),
.Y(n_487)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_L g488 ( 
.A(n_443),
.B(n_465),
.Y(n_488)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_454),
.C(n_459),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_459),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_445),
.Y(n_627)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_449),
.Y(n_561)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_469),
.Y(n_468)
);

OAI211xp5_ASAP7_75t_L g517 ( 
.A1(n_457),
.A2(n_518),
.B(n_522),
.C(n_526),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_457),
.B(n_600),
.Y(n_599)
);

OAI21xp33_ASAP7_75t_SL g614 ( 
.A1(n_457),
.A2(n_508),
.B(n_599),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_457),
.B(n_628),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_457),
.B(n_661),
.Y(n_660)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_461),
.Y(n_474)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_487),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_467),
.B(n_487),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_470),
.C(n_471),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g550 ( 
.A(n_468),
.B(n_551),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_470),
.A2(n_471),
.B1(n_472),
.B2(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_470),
.Y(n_552)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_476),
.C(n_485),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_473),
.B(n_501),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_476),
.A2(n_485),
.B1(n_486),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_476),
.Y(n_502)
);

INVxp33_ASAP7_75t_SL g548 ( 
.A(n_477),
.Y(n_548)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_482),
.Y(n_647)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_488),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_492),
.B(n_493),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_675),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_496),
.A2(n_553),
.B(n_673),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_550),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_498),
.B(n_674),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_503),
.C(n_515),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_500),
.B(n_556),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_503),
.A2(n_504),
.B1(n_515),
.B2(n_557),
.Y(n_556)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_505),
.A2(n_506),
.B(n_514),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_512),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_514),
.B(n_613),
.Y(n_612)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_538),
.Y(n_515)
);

XOR2x1_ASAP7_75t_L g578 ( 
.A(n_516),
.B(n_538),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_530),
.Y(n_516)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_533),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_534),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_SL g621 ( 
.A(n_539),
.B(n_622),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_541),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g674 ( 
.A(n_550),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g553 ( 
.A1(n_554),
.A2(n_579),
.B(n_672),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_555),
.B(n_558),
.Y(n_554)
);

NOR2x1_ASAP7_75t_L g672 ( 
.A(n_555),
.B(n_558),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_SL g558 ( 
.A(n_559),
.B(n_566),
.C(n_578),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_559),
.B(n_567),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_560),
.A2(n_626),
.B1(n_627),
.B2(n_628),
.Y(n_625)
);

BUFx4f_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

BUFx2_ASAP7_75t_SL g570 ( 
.A(n_571),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_578),
.B(n_632),
.Y(n_631)
);

OAI321xp33_ASAP7_75t_L g579 ( 
.A1(n_580),
.A2(n_629),
.A3(n_633),
.B1(n_670),
.B2(n_671),
.C(n_710),
.Y(n_579)
);

NOR2xp67_ASAP7_75t_L g580 ( 
.A(n_581),
.B(n_615),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_581),
.B(n_615),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_582),
.B(n_612),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_582),
.B(n_612),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_583),
.A2(n_593),
.B1(n_598),
.B2(n_603),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_588),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_604),
.B(n_610),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_611),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_616),
.B(n_623),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_616),
.B(n_624),
.C(n_625),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_617),
.Y(n_638)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

BUFx2_ASAP7_75t_SL g619 ( 
.A(n_620),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_624),
.B(n_625),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_630),
.B(n_631),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_630),
.B(n_631),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_634),
.A2(n_649),
.B(n_669),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_635),
.B(n_648),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_635),
.B(n_648),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_640),
.A2(n_653),
.B(n_656),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_642),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

BUFx2_ASAP7_75t_SL g643 ( 
.A(n_644),
.Y(n_643)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_647),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_SL g649 ( 
.A1(n_650),
.A2(n_657),
.B(n_668),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_651),
.B(n_652),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_651),
.B(n_652),
.Y(n_668)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_654),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_655),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_658),
.B(n_659),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_SL g659 ( 
.A(n_660),
.B(n_665),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_662),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_663),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_666),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_667),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_680),
.A2(n_682),
.B(n_683),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_681),
.Y(n_680)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_684),
.Y(n_683)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_686),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_688),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_SL g708 ( 
.A(n_688),
.B(n_702),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_689),
.B(n_700),
.Y(n_688)
);

NAND2x1_ASAP7_75t_L g689 ( 
.A(n_690),
.B(n_692),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_691),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_691),
.B(n_693),
.Y(n_701)
);

CKINVDCx16_ASAP7_75t_R g692 ( 
.A(n_693),
.Y(n_692)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_696),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_697),
.Y(n_696)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_699),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_701),
.Y(n_700)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_702),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_705),
.B(n_706),
.Y(n_704)
);


endmodule