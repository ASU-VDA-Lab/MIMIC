module fake_jpeg_31883_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_5),
.B(n_21),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_43),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_38),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_44),
.B1(n_45),
.B2(n_41),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_0),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_70)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_62),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_54),
.B1(n_42),
.B2(n_9),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_66),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_7),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_3),
.B(n_4),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_10),
.B(n_13),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_39),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_46),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_78),
.B1(n_82),
.B2(n_67),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_23),
.B(n_35),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_78),
.B(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_77),
.Y(n_90)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_37),
.B1(n_18),
.B2(n_11),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_84),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_15),
.B(n_17),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_85),
.B(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_14),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_27),
.C(n_28),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_77),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_97),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_89),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_72),
.A3(n_86),
.B1(n_71),
.B2(n_89),
.C1(n_33),
.C2(n_30),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_99),
.C(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_105),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_104),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_106),
.B(n_96),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_29),
.B(n_31),
.Y(n_111)
);

AOI221xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_32),
.B1(n_76),
.B2(n_74),
.C(n_63),
.Y(n_112)
);


endmodule