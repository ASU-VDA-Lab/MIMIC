module real_aes_252_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_847, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_847;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g571 ( .A(n_0), .B(n_140), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_1), .A2(n_106), .B1(n_834), .B2(n_843), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_2), .B(n_842), .Y(n_841) );
OAI22xp5_ASAP7_75t_SL g828 ( .A1(n_3), .A2(n_12), .B1(n_829), .B2(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g830 ( .A(n_3), .Y(n_830) );
INVx1_ASAP7_75t_L g147 ( .A(n_4), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_5), .B(n_505), .Y(n_531) );
NAND2xp33_ASAP7_75t_SL g590 ( .A(n_6), .B(n_146), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g118 ( .A(n_7), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g583 ( .A(n_8), .Y(n_583) );
INVx1_ASAP7_75t_L g196 ( .A(n_9), .Y(n_196) );
CKINVDCx16_ASAP7_75t_R g842 ( .A(n_10), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_11), .Y(n_187) );
AND2x2_ASAP7_75t_L g529 ( .A(n_12), .B(n_174), .Y(n_529) );
INVxp67_ASAP7_75t_L g829 ( .A(n_12), .Y(n_829) );
INVx2_ASAP7_75t_L g121 ( .A(n_13), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_14), .Y(n_491) );
AND3x1_ASAP7_75t_L g839 ( .A(n_14), .B(n_38), .C(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g141 ( .A(n_15), .Y(n_141) );
AOI221x1_ASAP7_75t_L g586 ( .A1(n_16), .A2(n_153), .B1(n_507), .B2(n_587), .C(n_589), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_17), .B(n_505), .Y(n_552) );
INVx1_ASAP7_75t_L g807 ( .A(n_18), .Y(n_807) );
INVx1_ASAP7_75t_L g494 ( .A(n_19), .Y(n_494) );
INVx1_ASAP7_75t_L g138 ( .A(n_20), .Y(n_138) );
INVx1_ASAP7_75t_SL g257 ( .A(n_21), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_22), .B(n_132), .Y(n_230) );
AOI33xp33_ASAP7_75t_L g206 ( .A1(n_23), .A2(n_54), .A3(n_126), .B1(n_167), .B2(n_207), .B3(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_24), .A2(n_507), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_25), .B(n_140), .Y(n_534) );
AOI221xp5_ASAP7_75t_SL g561 ( .A1(n_26), .A2(n_43), .B1(n_505), .B2(n_507), .C(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g181 ( .A(n_27), .Y(n_181) );
OAI22x1_ASAP7_75t_R g798 ( .A1(n_28), .A2(n_52), .B1(n_799), .B2(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_28), .Y(n_800) );
OR2x2_ASAP7_75t_L g120 ( .A(n_29), .B(n_93), .Y(n_120) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_29), .A2(n_93), .B(n_121), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_30), .B(n_143), .Y(n_556) );
INVxp67_ASAP7_75t_L g585 ( .A(n_31), .Y(n_585) );
AND2x2_ASAP7_75t_L g526 ( .A(n_32), .B(n_173), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_33), .B(n_158), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_34), .A2(n_507), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_35), .B(n_143), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_36), .A2(n_53), .B1(n_343), .B2(n_825), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_36), .Y(n_825) );
AND2x2_ASAP7_75t_L g146 ( .A(n_37), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g162 ( .A(n_37), .B(n_129), .Y(n_162) );
INVx1_ASAP7_75t_L g166 ( .A(n_37), .Y(n_166) );
OR2x6_ASAP7_75t_L g492 ( .A(n_38), .B(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_39), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_40), .B(n_158), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_41), .A2(n_119), .B1(n_154), .B2(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_42), .B(n_232), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_44), .A2(n_85), .B1(n_164), .B2(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_45), .B(n_132), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_46), .B(n_140), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_47), .B(n_193), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_48), .B(n_132), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_49), .Y(n_227) );
AND2x2_ASAP7_75t_L g574 ( .A(n_50), .B(n_173), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_51), .B(n_173), .Y(n_565) );
INVx1_ASAP7_75t_L g799 ( .A(n_52), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_53), .Y(n_343) );
HB1xp67_ASAP7_75t_SL g414 ( .A(n_53), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_55), .B(n_132), .Y(n_171) );
OAI22x1_ASAP7_75t_R g823 ( .A1(n_56), .A2(n_824), .B1(n_826), .B2(n_827), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_56), .Y(n_827) );
INVx1_ASAP7_75t_L g127 ( .A(n_57), .Y(n_127) );
INVx1_ASAP7_75t_L g134 ( .A(n_57), .Y(n_134) );
AND2x2_ASAP7_75t_L g172 ( .A(n_58), .B(n_173), .Y(n_172) );
AOI221xp5_ASAP7_75t_L g194 ( .A1(n_59), .A2(n_78), .B1(n_158), .B2(n_164), .C(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_60), .B(n_158), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_61), .B(n_505), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_62), .B(n_154), .Y(n_189) );
XNOR2xp5_ASAP7_75t_L g794 ( .A(n_63), .B(n_795), .Y(n_794) );
AOI21xp5_ASAP7_75t_SL g216 ( .A1(n_64), .A2(n_164), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g517 ( .A(n_65), .B(n_173), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_66), .B(n_143), .Y(n_572) );
INVx1_ASAP7_75t_L g124 ( .A(n_67), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_68), .B(n_140), .Y(n_515) );
AND2x2_ASAP7_75t_SL g557 ( .A(n_69), .B(n_174), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_70), .A2(n_507), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g170 ( .A(n_71), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_72), .B(n_143), .Y(n_535) );
AND2x2_ASAP7_75t_SL g508 ( .A(n_73), .B(n_193), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_74), .A2(n_164), .B(n_169), .Y(n_163) );
INVx1_ASAP7_75t_L g129 ( .A(n_75), .Y(n_129) );
INVx1_ASAP7_75t_L g136 ( .A(n_75), .Y(n_136) );
AOI22x1_ASAP7_75t_L g795 ( .A1(n_76), .A2(n_796), .B1(n_797), .B2(n_798), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_76), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_77), .B(n_158), .Y(n_209) );
AND2x2_ASAP7_75t_L g259 ( .A(n_79), .B(n_153), .Y(n_259) );
INVx1_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_81), .A2(n_164), .B(n_256), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_82), .A2(n_164), .B(n_201), .C(n_229), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_83), .A2(n_88), .B1(n_158), .B2(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_84), .B(n_505), .Y(n_516) );
INVx1_ASAP7_75t_L g495 ( .A(n_86), .Y(n_495) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_87), .B(n_153), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_89), .A2(n_164), .B1(n_204), .B2(n_205), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_90), .B(n_140), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_91), .B(n_140), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_92), .A2(n_507), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g218 ( .A(n_94), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_95), .B(n_143), .Y(n_514) );
AND2x2_ASAP7_75t_L g210 ( .A(n_96), .B(n_153), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_97), .A2(n_179), .B(n_180), .C(n_182), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_98), .B(n_505), .Y(n_573) );
INVxp67_ASAP7_75t_L g588 ( .A(n_99), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_100), .B(n_143), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_101), .A2(n_507), .B(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g813 ( .A(n_102), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_103), .B(n_132), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_104), .B(n_815), .Y(n_814) );
OA22x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_810), .B1(n_813), .B2(n_818), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_801), .Y(n_107) );
NAND2xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_793), .Y(n_108) );
OAI22xp5_ASAP7_75t_SL g109 ( .A1(n_110), .A2(n_487), .B1(n_496), .B2(n_789), .Y(n_109) );
INVx1_ASAP7_75t_L g804 ( .A(n_110), .Y(n_804) );
AOI211x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_343), .B(n_344), .C(n_484), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND4x1_ASAP7_75t_L g484 ( .A(n_112), .B(n_345), .C(n_485), .D(n_486), .Y(n_484) );
NAND3x1_ASAP7_75t_L g821 ( .A(n_112), .B(n_345), .C(n_822), .Y(n_821) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_311), .Y(n_112) );
AOI211xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_233), .B(n_245), .C(n_287), .Y(n_113) );
OAI21xp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_148), .B(n_211), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_SL g233 ( .A1(n_116), .A2(n_234), .B(n_239), .C(n_244), .Y(n_233) );
NAND2x1_ASAP7_75t_L g364 ( .A(n_116), .B(n_365), .Y(n_364) );
NOR2x1_ASAP7_75t_L g455 ( .A(n_116), .B(n_384), .Y(n_455) );
AND2x2_ASAP7_75t_L g474 ( .A(n_116), .B(n_213), .Y(n_474) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx3_ASAP7_75t_L g250 ( .A(n_117), .Y(n_250) );
AND2x2_ASAP7_75t_L g322 ( .A(n_117), .B(n_251), .Y(n_322) );
AND2x2_ASAP7_75t_L g327 ( .A(n_117), .B(n_222), .Y(n_327) );
NOR2x1_ASAP7_75t_SL g443 ( .A(n_117), .B(n_213), .Y(n_443) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_119), .B(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_119), .A2(n_216), .B(n_220), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_119), .A2(n_531), .B(n_532), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_119), .B(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_119), .B(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_119), .B(n_588), .Y(n_587) );
NOR3xp33_ASAP7_75t_L g589 ( .A(n_119), .B(n_131), .C(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_120), .B(n_121), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_137), .B(n_144), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_130), .B2(n_131), .Y(n_123) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_125), .A2(n_145), .B(n_170), .C(n_171), .Y(n_169) );
INVxp67_ASAP7_75t_L g179 ( .A(n_125), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_SL g195 ( .A1(n_125), .A2(n_145), .B(n_196), .C(n_197), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_125), .A2(n_145), .B(n_218), .C(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g232 ( .A(n_125), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g256 ( .A1(n_125), .A2(n_145), .B(n_257), .C(n_258), .Y(n_256) );
OR2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
AND2x2_ASAP7_75t_L g159 ( .A(n_126), .B(n_160), .Y(n_159) );
INVxp33_ASAP7_75t_L g207 ( .A(n_126), .Y(n_207) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g143 ( .A(n_127), .B(n_135), .Y(n_143) );
AND2x2_ASAP7_75t_L g168 ( .A(n_127), .B(n_147), .Y(n_168) );
INVx3_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x6_ASAP7_75t_L g140 ( .A(n_129), .B(n_133), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_131), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g505 ( .A(n_132), .B(n_146), .Y(n_505) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B1(n_141), .B2(n_142), .Y(n_137) );
INVxp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVxp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_145), .A2(n_230), .B(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_145), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_145), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_145), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_145), .A2(n_555), .B(n_556), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_145), .A2(n_563), .B(n_564), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_145), .A2(n_571), .B(n_572), .Y(n_570) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_147), .Y(n_160) );
INVx1_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_191), .Y(n_149) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_150), .B(n_292), .Y(n_358) );
AND2x2_ASAP7_75t_L g475 ( .A(n_150), .B(n_316), .Y(n_475) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_175), .Y(n_150) );
NOR2x1_ASAP7_75t_L g242 ( .A(n_151), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g264 ( .A(n_151), .Y(n_264) );
AND2x2_ASAP7_75t_L g272 ( .A(n_151), .B(n_273), .Y(n_272) );
NOR2xp67_ASAP7_75t_L g410 ( .A(n_151), .B(n_175), .Y(n_410) );
AO21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_156), .B(n_172), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_152), .A2(n_153), .B1(n_178), .B2(n_183), .Y(n_177) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_152), .A2(n_156), .B(n_172), .Y(n_295) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_154), .B(n_186), .Y(n_185) );
AOI21x1_ASAP7_75t_L g567 ( .A1(n_154), .A2(n_568), .B(n_574), .Y(n_567) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx4f_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_163), .Y(n_156) );
INVx1_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_158), .A2(n_164), .B1(n_582), .B2(n_584), .Y(n_581) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_161), .Y(n_158) );
INVx1_ASAP7_75t_L g225 ( .A(n_159), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_161), .Y(n_226) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x6_ASAP7_75t_L g507 ( .A(n_162), .B(n_168), .Y(n_507) );
INVxp67_ASAP7_75t_L g188 ( .A(n_164), .Y(n_188) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_168), .Y(n_164) );
NOR2x1p5_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx1_ASAP7_75t_L g208 ( .A(n_167), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_173), .Y(n_252) );
OA21x2_ASAP7_75t_L g560 ( .A1(n_173), .A2(n_561), .B(n_565), .Y(n_560) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g362 ( .A(n_175), .B(n_200), .Y(n_362) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x4_ASAP7_75t_L g237 ( .A(n_176), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g241 ( .A(n_176), .Y(n_241) );
INVx1_ASAP7_75t_L g262 ( .A(n_176), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_176), .B(n_295), .Y(n_319) );
AND2x2_ASAP7_75t_L g368 ( .A(n_176), .B(n_192), .Y(n_368) );
OR2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_184), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_188), .B1(n_189), .B2(n_190), .Y(n_184) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g323 ( .A(n_191), .B(n_318), .Y(n_323) );
AND2x2_ASAP7_75t_L g379 ( .A(n_191), .B(n_262), .Y(n_379) );
AND2x2_ASAP7_75t_L g394 ( .A(n_191), .B(n_308), .Y(n_394) );
AND2x2_ASAP7_75t_L g431 ( .A(n_191), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g447 ( .A(n_191), .Y(n_447) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_199), .Y(n_191) );
INVx2_ASAP7_75t_L g238 ( .A(n_192), .Y(n_238) );
INVx1_ASAP7_75t_L g243 ( .A(n_192), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_192), .B(n_274), .Y(n_277) );
INVx1_ASAP7_75t_L g291 ( .A(n_192), .Y(n_291) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_192), .Y(n_301) );
INVxp67_ASAP7_75t_L g317 ( .A(n_192), .Y(n_317) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_198), .Y(n_192) );
INVx2_ASAP7_75t_SL g201 ( .A(n_193), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_193), .A2(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g235 ( .A(n_200), .Y(n_235) );
AND2x4_ASAP7_75t_L g263 ( .A(n_200), .B(n_264), .Y(n_263) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_210), .Y(n_200) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_201), .A2(n_202), .B(n_210), .Y(n_274) );
AOI21x1_ASAP7_75t_L g502 ( .A1(n_201), .A2(n_503), .B(n_508), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_203), .B(n_209), .Y(n_202) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g244 ( .A(n_211), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_211), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_SL g266 ( .A(n_212), .B(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_212), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_212), .B(n_280), .Y(n_423) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_212), .Y(n_461) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_221), .Y(n_212) );
INVx2_ASAP7_75t_L g286 ( .A(n_213), .Y(n_286) );
AND2x2_ASAP7_75t_L g297 ( .A(n_213), .B(n_222), .Y(n_297) );
INVx4_ASAP7_75t_L g305 ( .A(n_213), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_213), .B(n_281), .Y(n_341) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_213), .Y(n_354) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AND2x4_ASAP7_75t_L g332 ( .A(n_221), .B(n_305), .Y(n_332) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x4_ASAP7_75t_L g283 ( .A(n_222), .B(n_250), .Y(n_283) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_222), .Y(n_304) );
INVx2_ASAP7_75t_L g353 ( .A(n_222), .Y(n_353) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_228), .Y(n_222) );
NOR3xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .C(n_227), .Y(n_224) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_235), .B(n_240), .Y(n_342) );
NAND2x1_ASAP7_75t_SL g456 ( .A(n_235), .B(n_237), .Y(n_456) );
OR2x2_ASAP7_75t_L g335 ( .A(n_236), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g438 ( .A(n_236), .Y(n_438) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g328 ( .A(n_237), .B(n_263), .Y(n_328) );
AND2x2_ASAP7_75t_L g444 ( .A(n_237), .B(n_437), .Y(n_444) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_239), .A2(n_453), .B1(n_456), .B2(n_457), .C(n_459), .Y(n_452) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_240), .A2(n_397), .B1(n_399), .B2(n_401), .Y(n_396) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_241), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g310 ( .A(n_241), .Y(n_310) );
BUFx2_ASAP7_75t_L g391 ( .A(n_241), .Y(n_391) );
AND2x2_ASAP7_75t_L g361 ( .A(n_242), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_246), .B(n_265), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_260), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_SL g334 ( .A(n_249), .Y(n_334) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_249), .B(n_460), .C(n_461), .D(n_462), .Y(n_459) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g269 ( .A(n_250), .Y(n_269) );
AND2x2_ASAP7_75t_L g352 ( .A(n_250), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g268 ( .A(n_251), .Y(n_268) );
INVx2_ASAP7_75t_L g282 ( .A(n_251), .Y(n_282) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_251), .Y(n_309) );
INVx1_ASAP7_75t_L g326 ( .A(n_251), .Y(n_326) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_251), .Y(n_366) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B(n_259), .Y(n_251) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_252), .A2(n_511), .B(n_517), .Y(n_510) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_252), .A2(n_520), .B(n_526), .Y(n_519) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_252), .A2(n_520), .B(n_526), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g473 ( .A(n_261), .Y(n_473) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g271 ( .A(n_262), .Y(n_271) );
AND2x2_ASAP7_75t_L g367 ( .A(n_263), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g467 ( .A(n_263), .B(n_468), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_270), .B1(n_275), .B2(n_278), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_267), .B(n_332), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_267), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g448 ( .A(n_267), .B(n_426), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_267), .A2(n_303), .B(n_425), .Y(n_478) );
AND2x4_ASAP7_75t_SL g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_268), .B(n_352), .Y(n_389) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_268), .Y(n_405) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AND2x2_ASAP7_75t_L g275 ( .A(n_271), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g292 ( .A(n_273), .Y(n_292) );
AND2x2_ASAP7_75t_L g316 ( .A(n_273), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g437 ( .A(n_273), .B(n_294), .Y(n_437) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_274), .B(n_295), .Y(n_336) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g412 ( .A(n_277), .B(n_319), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_284), .Y(n_278) );
INVx1_ASAP7_75t_L g393 ( .A(n_279), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
NOR3xp33_ASAP7_75t_L g288 ( .A(n_280), .B(n_289), .C(n_293), .Y(n_288) );
AND2x2_ASAP7_75t_L g331 ( .A(n_280), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g360 ( .A(n_280), .B(n_303), .Y(n_360) );
AND2x2_ASAP7_75t_L g442 ( .A(n_280), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g468 ( .A(n_280), .Y(n_468) );
INVx1_ASAP7_75t_L g482 ( .A(n_280), .Y(n_482) );
INVx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g285 ( .A(n_283), .B(n_286), .Y(n_285) );
INVx4_ASAP7_75t_L g441 ( .A(n_283), .Y(n_441) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g481 ( .A(n_285), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g384 ( .A(n_286), .Y(n_384) );
AO22x1_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_296), .B1(n_298), .B2(n_306), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_290), .B(n_294), .Y(n_374) );
INVx3_ASAP7_75t_L g408 ( .A(n_290), .Y(n_408) );
BUFx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g308 ( .A(n_294), .Y(n_308) );
INVx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g386 ( .A(n_295), .B(n_301), .Y(n_386) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_295), .Y(n_433) );
AOI31xp33_ASAP7_75t_L g337 ( .A1(n_296), .A2(n_338), .A3(n_340), .B(n_342), .Y(n_337) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI22xp33_ASAP7_75t_SL g313 ( .A1(n_297), .A2(n_314), .B1(n_320), .B2(n_323), .Y(n_313) );
AND2x2_ASAP7_75t_L g397 ( .A(n_297), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g404 ( .A(n_297), .B(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_303), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_SL g303 ( .A(n_304), .B(n_305), .Y(n_303) );
OR2x2_ASAP7_75t_L g333 ( .A(n_305), .B(n_334), .Y(n_333) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_305), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_310), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x2_ASAP7_75t_L g428 ( .A(n_308), .B(n_368), .Y(n_428) );
INVx1_ASAP7_75t_L g463 ( .A(n_308), .Y(n_463) );
AND2x2_ASAP7_75t_L g413 ( .A(n_309), .B(n_352), .Y(n_413) );
BUFx2_ASAP7_75t_L g458 ( .A(n_309), .Y(n_458) );
AND2x2_ASAP7_75t_L g401 ( .A(n_310), .B(n_402), .Y(n_401) );
NOR3xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_329), .C(n_337), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_313), .B(n_324), .Y(n_312) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
AND2x2_ASAP7_75t_L g390 ( .A(n_316), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_322), .B(n_332), .Y(n_355) );
AND2x2_ASAP7_75t_L g377 ( .A(n_322), .B(n_354), .Y(n_377) );
AND2x2_ASAP7_75t_SL g425 ( .A(n_322), .B(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
AND2x2_ASAP7_75t_L g480 ( .A(n_325), .B(n_354), .Y(n_480) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g454 ( .A(n_326), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g371 ( .A(n_327), .Y(n_371) );
AND2x2_ASAP7_75t_L g471 ( .A(n_327), .B(n_354), .Y(n_471) );
AOI21xp33_ASAP7_75t_R g329 ( .A1(n_330), .A2(n_333), .B(n_335), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_331), .B(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_332), .Y(n_339) );
INVx1_ASAP7_75t_L g402 ( .A(n_336), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_338), .A2(n_356), .B1(n_370), .B2(n_372), .Y(n_369) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g370 ( .A(n_341), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_343), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_343), .B(n_450), .Y(n_449) );
NOR2xp67_ASAP7_75t_SL g485 ( .A(n_343), .B(n_416), .Y(n_485) );
OAI211xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_414), .B(n_415), .C(n_449), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_380), .Y(n_345) );
NOR3xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_369), .C(n_375), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_356), .B(n_359), .Y(n_347) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_355), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_351), .A2(n_390), .B1(n_393), .B2(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_SL g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g427 ( .A(n_353), .Y(n_427) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g419 ( .A(n_358), .B(n_408), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_363), .B2(n_367), .Y(n_359) );
INVx1_ASAP7_75t_L g373 ( .A(n_362), .Y(n_373) );
AND2x4_ASAP7_75t_L g385 ( .A(n_362), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g421 ( .A(n_364), .Y(n_421) );
INVx1_ASAP7_75t_L g398 ( .A(n_365), .Y(n_398) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_367), .A2(n_377), .B1(n_425), .B2(n_428), .Y(n_424) );
INVxp67_ASAP7_75t_L g469 ( .A(n_368), .Y(n_469) );
NOR2x1_ASAP7_75t_L g383 ( .A(n_371), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVxp33_ASAP7_75t_L g483 ( .A(n_374), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_395), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_382), .B(n_392), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B1(n_387), .B2(n_390), .Y(n_382) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_396), .B(n_403), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B1(n_411), .B2(n_413), .Y(n_403) );
NOR2xp33_ASAP7_75t_SL g406 ( .A(n_407), .B(n_409), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g460 ( .A(n_408), .Y(n_460) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g822 ( .A(n_417), .B(n_451), .Y(n_822) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_418), .B(n_429), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_424), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND4xp25_ASAP7_75t_SL g429 ( .A(n_430), .B(n_434), .C(n_439), .D(n_445), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g472 ( .A(n_437), .B(n_473), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .B(n_444), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g486 ( .A(n_450), .Y(n_486) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR3x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_464), .C(n_476), .Y(n_451) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_469), .B(n_470), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_474), .B2(n_475), .Y(n_470) );
INVx1_ASAP7_75t_L g477 ( .A(n_475), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_479), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_483), .Y(n_479) );
CKINVDCx6p67_ASAP7_75t_R g487 ( .A(n_488), .Y(n_487) );
CKINVDCx11_ASAP7_75t_R g805 ( .A(n_488), .Y(n_805) );
INVx3_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_490), .Y(n_489) );
AND2x6_ASAP7_75t_SL g490 ( .A(n_491), .B(n_492), .Y(n_490) );
OR2x6_ASAP7_75t_SL g791 ( .A(n_491), .B(n_792), .Y(n_791) );
OR2x2_ASAP7_75t_L g809 ( .A(n_491), .B(n_492), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_491), .B(n_792), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_492), .Y(n_792) );
INVx1_ASAP7_75t_L g838 ( .A(n_493), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g803 ( .A(n_496), .Y(n_803) );
AND3x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_660), .C(n_734), .Y(n_496) );
NOR3xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_602), .C(n_633), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_538), .B(n_547), .C(n_575), .Y(n_498) );
AOI21x1_ASAP7_75t_SL g499 ( .A1(n_500), .A2(n_518), .B(n_536), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_500), .A2(n_636), .B1(n_642), .B2(n_645), .Y(n_635) );
AND2x2_ASAP7_75t_L g769 ( .A(n_500), .B(n_540), .Y(n_769) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_509), .Y(n_500) );
BUFx2_ASAP7_75t_L g543 ( .A(n_501), .Y(n_543) );
AND2x2_ASAP7_75t_L g628 ( .A(n_501), .B(n_510), .Y(n_628) );
AND2x2_ASAP7_75t_L g699 ( .A(n_501), .B(n_546), .Y(n_699) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_502), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
AND2x4_ASAP7_75t_L g592 ( .A(n_509), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g537 ( .A(n_510), .B(n_528), .Y(n_537) );
OR2x2_ASAP7_75t_L g545 ( .A(n_510), .B(n_546), .Y(n_545) );
AND2x4_ASAP7_75t_L g597 ( .A(n_510), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g644 ( .A(n_510), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_510), .B(n_546), .Y(n_652) );
AND2x2_ASAP7_75t_L g689 ( .A(n_510), .B(n_593), .Y(n_689) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_510), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_510), .B(n_527), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_516), .Y(n_511) );
INVx2_ASAP7_75t_L g631 ( .A(n_518), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_518), .B(n_592), .Y(n_687) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_518), .Y(n_788) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_527), .Y(n_518) );
AND2x2_ASAP7_75t_L g536 ( .A(n_519), .B(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g613 ( .A(n_519), .B(n_528), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_519), .B(n_644), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
AND2x2_ASAP7_75t_L g680 ( .A(n_527), .B(n_597), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_527), .B(n_592), .Y(n_736) );
INVx5_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g541 ( .A(n_528), .Y(n_541) );
AND2x2_ASAP7_75t_L g607 ( .A(n_528), .B(n_598), .Y(n_607) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_528), .Y(n_627) );
AND2x4_ASAP7_75t_L g634 ( .A(n_528), .B(n_546), .Y(n_634) );
AND2x2_ASAP7_75t_SL g781 ( .A(n_528), .B(n_593), .Y(n_781) );
OR2x6_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g760 ( .A(n_536), .Y(n_760) );
INVx1_ASAP7_75t_L g702 ( .A(n_537), .Y(n_702) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g624 ( .A(n_541), .B(n_545), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_541), .B(n_593), .Y(n_717) );
AND2x2_ASAP7_75t_L g719 ( .A(n_541), .B(n_544), .Y(n_719) );
AOI32xp33_ASAP7_75t_L g785 ( .A1(n_541), .A2(n_601), .A3(n_756), .B1(n_786), .B2(n_788), .Y(n_785) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
AND2x2_ASAP7_75t_L g611 ( .A(n_543), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g729 ( .A(n_543), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g752 ( .A(n_543), .B(n_613), .Y(n_752) );
AND2x2_ASAP7_75t_L g779 ( .A(n_543), .B(n_680), .Y(n_779) );
AND2x2_ASAP7_75t_L g705 ( .A(n_544), .B(n_593), .Y(n_705) );
AND2x2_ASAP7_75t_L g780 ( .A(n_544), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g598 ( .A(n_546), .Y(n_598) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_558), .Y(n_548) );
NOR2x1p5_ASAP7_75t_L g638 ( .A(n_549), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g656 ( .A(n_549), .Y(n_656) );
OR2x2_ASAP7_75t_L g684 ( .A(n_549), .B(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_SL g601 ( .A(n_550), .B(n_580), .Y(n_601) );
AND2x4_ASAP7_75t_L g617 ( .A(n_550), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g620 ( .A(n_550), .B(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g648 ( .A(n_550), .B(n_560), .Y(n_648) );
OR2x2_ASAP7_75t_L g673 ( .A(n_550), .B(n_622), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_550), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_550), .B(n_560), .Y(n_708) );
INVx2_ASAP7_75t_L g724 ( .A(n_550), .Y(n_724) );
AND2x2_ASAP7_75t_L g739 ( .A(n_550), .B(n_579), .Y(n_739) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_550), .Y(n_763) );
INVx1_ASAP7_75t_L g768 ( .A(n_550), .Y(n_768) );
OR2x6_ASAP7_75t_L g550 ( .A(n_551), .B(n_557), .Y(n_550) );
AND2x2_ASAP7_75t_L g632 ( .A(n_558), .B(n_617), .Y(n_632) );
AND2x2_ASAP7_75t_L g653 ( .A(n_558), .B(n_601), .Y(n_653) );
INVx1_ASAP7_75t_L g685 ( .A(n_558), .Y(n_685) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_566), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g578 ( .A(n_560), .Y(n_578) );
INVx2_ASAP7_75t_L g622 ( .A(n_560), .Y(n_622) );
BUFx3_ASAP7_75t_L g639 ( .A(n_560), .Y(n_639) );
AND2x2_ASAP7_75t_L g678 ( .A(n_560), .B(n_566), .Y(n_678) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_560), .Y(n_776) );
INVx2_ASAP7_75t_L g591 ( .A(n_566), .Y(n_591) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_566), .Y(n_600) );
INVx1_ASAP7_75t_L g616 ( .A(n_566), .Y(n_616) );
OR2x2_ASAP7_75t_L g621 ( .A(n_566), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g641 ( .A(n_566), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_566), .B(n_618), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_566), .B(n_724), .Y(n_723) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_573), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_592), .B(n_594), .Y(n_575) );
AND2x2_ASAP7_75t_SL g576 ( .A(n_577), .B(n_579), .Y(n_576) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_577), .Y(n_784) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_578), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_578), .B(n_616), .Y(n_658) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_578), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_579), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g663 ( .A(n_579), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g714 ( .A(n_579), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_579), .A2(n_719), .B1(n_720), .B2(n_725), .C(n_728), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_579), .B(n_768), .Y(n_767) );
AND2x4_ASAP7_75t_L g579 ( .A(n_580), .B(n_591), .Y(n_579) );
INVx3_ASAP7_75t_L g618 ( .A(n_580), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_580), .B(n_622), .Y(n_722) );
AND2x2_ASAP7_75t_L g751 ( .A(n_580), .B(n_724), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_580), .B(n_783), .Y(n_782) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_586), .Y(n_580) );
AND2x2_ASAP7_75t_L g659 ( .A(n_592), .B(n_634), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_592), .A2(n_612), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g596 ( .A(n_593), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g605 ( .A(n_593), .Y(n_605) );
OR2x2_ASAP7_75t_L g651 ( .A(n_593), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_593), .B(n_634), .Y(n_743) );
OR2x2_ASAP7_75t_L g775 ( .A(n_593), .B(n_776), .Y(n_775) );
OR2x2_ASAP7_75t_L g787 ( .A(n_593), .B(n_693), .Y(n_787) );
INVxp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
INVx2_ASAP7_75t_L g665 ( .A(n_596), .Y(n_665) );
INVx3_ASAP7_75t_SL g731 ( .A(n_597), .Y(n_731) );
INVxp67_ASAP7_75t_L g681 ( .A(n_599), .Y(n_681) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AOI322xp5_ASAP7_75t_L g603 ( .A1(n_601), .A2(n_604), .A3(n_608), .B1(n_611), .B2(n_614), .C1(n_619), .C2(n_623), .Y(n_603) );
INVx1_ASAP7_75t_SL g692 ( .A(n_601), .Y(n_692) );
AND2x4_ASAP7_75t_L g777 ( .A(n_601), .B(n_664), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_625), .Y(n_602) );
NOR2x1_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
OR2x2_ASAP7_75t_L g630 ( .A(n_605), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g726 ( .A(n_605), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g754 ( .A(n_605), .B(n_607), .Y(n_754) );
AOI32xp33_ASAP7_75t_L g755 ( .A1(n_605), .A2(n_606), .A3(n_756), .B1(n_758), .B2(n_761), .Y(n_755) );
OR2x2_ASAP7_75t_L g759 ( .A(n_605), .B(n_652), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g715 ( .A(n_606), .B(n_631), .C(n_716), .Y(n_715) );
OAI22xp33_ASAP7_75t_SL g735 ( .A1(n_606), .A2(n_672), .B1(n_736), .B2(n_737), .Y(n_735) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVxp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g738 ( .A(n_609), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_613), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
OAI322xp33_ASAP7_75t_L g661 ( .A1(n_617), .A2(n_621), .A3(n_630), .B1(n_662), .B2(n_665), .C1(n_666), .C2(n_667), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_617), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_617), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g640 ( .A(n_618), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g672 ( .A(n_618), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_618), .B(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g733 ( .A(n_621), .Y(n_733) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_622), .Y(n_664) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_629), .B(n_632), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_628), .B(n_676), .Y(n_675) );
AOI322xp5_ASAP7_75t_SL g770 ( .A1(n_628), .A2(n_634), .A3(n_751), .B1(n_769), .B2(n_771), .C1(n_774), .C2(n_777), .Y(n_770) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI21xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B(n_649), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_634), .B(n_644), .Y(n_666) );
INVx2_ASAP7_75t_SL g676 ( .A(n_634), .Y(n_676) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_SL g701 ( .A(n_640), .Y(n_701) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_641), .Y(n_671) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g746 ( .A(n_647), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g700 ( .A(n_648), .B(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B1(n_654), .B2(n_659), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR4xp75_ASAP7_75t_L g660 ( .A(n_661), .B(n_674), .C(n_694), .D(n_710), .Y(n_660) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_669), .B(n_672), .Y(n_668) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_672), .A2(n_749), .B1(n_752), .B2(n_753), .Y(n_748) );
OR2x2_ASAP7_75t_L g713 ( .A(n_673), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g757 ( .A(n_673), .Y(n_757) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B1(n_679), .B2(n_681), .C(n_682), .Y(n_674) );
INVx2_ASAP7_75t_L g693 ( .A(n_678), .Y(n_693) );
AND2x2_ASAP7_75t_L g750 ( .A(n_678), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_686), .B1(n_688), .B2(n_690), .Y(n_682) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g745 ( .A(n_689), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_690), .A2(n_696), .B1(n_712), .B2(n_715), .Y(n_711) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_700), .B1(n_702), .B2(n_703), .C(n_847), .Y(n_694) );
AND2x2_ASAP7_75t_SL g696 ( .A(n_697), .B(n_699), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g762 ( .A(n_701), .B(n_763), .Y(n_762) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g747 ( .A(n_709), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_718), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
AOI21xp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B(n_732), .Y(n_728) );
NOR3xp33_ASAP7_75t_SL g734 ( .A(n_735), .B(n_740), .C(n_764), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_755), .Y(n_740) );
O2A1O1Ixp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_744), .B(n_746), .C(n_748), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND2x4_ASAP7_75t_L g756 ( .A(n_747), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
NAND4xp25_ASAP7_75t_SL g764 ( .A(n_765), .B(n_770), .C(n_778), .D(n_785), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_769), .Y(n_765) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
OAI21xp5_ASAP7_75t_SL g778 ( .A1(n_779), .A2(n_780), .B(n_782), .Y(n_778) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx3_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
CKINVDCx11_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
OAI22x1_ASAP7_75t_L g802 ( .A1(n_791), .A2(n_803), .B1(n_804), .B2(n_805), .Y(n_802) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
AOI21xp33_ASAP7_75t_L g801 ( .A1(n_794), .A2(n_802), .B(n_806), .Y(n_801) );
CKINVDCx16_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
BUFx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_814), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_812), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_813), .Y(n_812) );
OAI21xp5_ASAP7_75t_L g818 ( .A1(n_814), .A2(n_819), .B(n_833), .Y(n_818) );
INVx1_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g833 ( .A(n_816), .Y(n_833) );
BUFx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_828), .B1(n_831), .B2(n_832), .Y(n_819) );
INVx2_ASAP7_75t_L g832 ( .A(n_820), .Y(n_832) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_821), .B(n_823), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_824), .Y(n_826) );
INVx1_ASAP7_75t_L g831 ( .A(n_828), .Y(n_831) );
BUFx4f_ASAP7_75t_SL g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_SL g845 ( .A(n_836), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_837), .Y(n_836) );
AND2x2_ASAP7_75t_SL g837 ( .A(n_838), .B(n_839), .Y(n_837) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx4_ASAP7_75t_SL g843 ( .A(n_844), .Y(n_843) );
BUFx4f_ASAP7_75t_SL g844 ( .A(n_845), .Y(n_844) );
endmodule