module real_aes_827_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_0), .B(n_149), .Y(n_172) );
AOI22xp5_ASAP7_75t_SL g125 ( .A1(n_1), .A2(n_126), .B1(n_129), .B2(n_130), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_1), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_2), .A2(n_143), .B(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_3), .B(n_796), .Y(n_795) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_4), .B(n_160), .Y(n_188) );
INVx1_ASAP7_75t_L g148 ( .A(n_5), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_6), .B(n_160), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_7), .B(n_184), .Y(n_568) );
INVx1_ASAP7_75t_L g485 ( .A(n_8), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g796 ( .A(n_9), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_10), .Y(n_501) );
NAND2xp33_ASAP7_75t_L g260 ( .A(n_11), .B(n_158), .Y(n_260) );
INVx2_ASAP7_75t_L g140 ( .A(n_12), .Y(n_140) );
AOI221x1_ASAP7_75t_L g142 ( .A1(n_13), .A2(n_25), .B1(n_143), .B2(n_149), .C(n_156), .Y(n_142) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_14), .Y(n_117) );
AND3x1_ASAP7_75t_L g793 ( .A(n_14), .B(n_38), .C(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_15), .B(n_149), .Y(n_256) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_16), .A2(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g576 ( .A(n_17), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_18), .B(n_138), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_19), .B(n_160), .Y(n_242) );
AO21x1_ASAP7_75t_L g182 ( .A1(n_20), .A2(n_149), .B(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g121 ( .A(n_21), .Y(n_121) );
INVx1_ASAP7_75t_L g574 ( .A(n_22), .Y(n_574) );
INVx1_ASAP7_75t_SL g539 ( .A(n_23), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_24), .B(n_150), .Y(n_560) );
NAND2x1_ASAP7_75t_L g170 ( .A(n_26), .B(n_160), .Y(n_170) );
AOI33xp33_ASAP7_75t_L g513 ( .A1(n_27), .A2(n_54), .A3(n_467), .B1(n_472), .B2(n_514), .B3(n_515), .Y(n_513) );
NAND2x1_ASAP7_75t_L g216 ( .A(n_28), .B(n_158), .Y(n_216) );
INVx1_ASAP7_75t_L g494 ( .A(n_29), .Y(n_494) );
OR2x2_ASAP7_75t_L g141 ( .A(n_30), .B(n_90), .Y(n_141) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_30), .A2(n_90), .B(n_140), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_31), .B(n_475), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_32), .B(n_158), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_33), .A2(n_95), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_33), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_34), .B(n_160), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_35), .B(n_158), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_36), .A2(n_143), .B(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g144 ( .A(n_37), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g155 ( .A(n_37), .B(n_148), .Y(n_155) );
INVx1_ASAP7_75t_L g466 ( .A(n_37), .Y(n_466) );
OR2x6_ASAP7_75t_L g119 ( .A(n_38), .B(n_120), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_39), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_40), .A2(n_51), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_40), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_41), .B(n_149), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_42), .B(n_475), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_43), .A2(n_175), .B1(n_184), .B2(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_44), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_45), .B(n_150), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_46), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_47), .B(n_158), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_48), .B(n_254), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_49), .B(n_150), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_50), .A2(n_143), .B(n_215), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_51), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_52), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_53), .B(n_158), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_55), .B(n_150), .Y(n_525) );
INVx1_ASAP7_75t_L g147 ( .A(n_56), .Y(n_147) );
INVx1_ASAP7_75t_L g152 ( .A(n_56), .Y(n_152) );
AND2x2_ASAP7_75t_L g526 ( .A(n_57), .B(n_138), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_58), .A2(n_76), .B1(n_464), .B2(n_475), .C(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_59), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_60), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_61), .B(n_175), .Y(n_503) );
AOI21xp5_ASAP7_75t_SL g463 ( .A1(n_62), .A2(n_464), .B(n_469), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_63), .A2(n_143), .B(n_169), .Y(n_168) );
XNOR2xp5_ASAP7_75t_L g447 ( .A(n_64), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g571 ( .A(n_65), .Y(n_571) );
AO21x1_ASAP7_75t_L g185 ( .A1(n_66), .A2(n_143), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_67), .B(n_149), .Y(n_206) );
INVx1_ASAP7_75t_L g524 ( .A(n_68), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_69), .B(n_149), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_70), .A2(n_464), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g199 ( .A(n_71), .B(n_139), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_72), .A2(n_447), .B1(n_452), .B2(n_779), .Y(n_446) );
INVx1_ASAP7_75t_L g145 ( .A(n_73), .Y(n_145) );
INVx1_ASAP7_75t_L g154 ( .A(n_73), .Y(n_154) );
AND2x2_ASAP7_75t_L g220 ( .A(n_74), .B(n_174), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_75), .B(n_475), .Y(n_516) );
AND2x2_ASAP7_75t_L g541 ( .A(n_77), .B(n_174), .Y(n_541) );
INVx1_ASAP7_75t_L g572 ( .A(n_78), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_79), .A2(n_464), .B(n_538), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_80), .A2(n_464), .B(n_508), .C(n_559), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_81), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_82), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g122 ( .A(n_83), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_83), .B(n_121), .Y(n_792) );
AND2x2_ASAP7_75t_L g204 ( .A(n_84), .B(n_174), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_85), .B(n_149), .Y(n_244) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_86), .B(n_174), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_87), .A2(n_464), .B1(n_511), .B2(n_512), .Y(n_510) );
XNOR2xp5_ASAP7_75t_L g448 ( .A(n_88), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g183 ( .A(n_89), .B(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g177 ( .A(n_91), .B(n_174), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_92), .B(n_158), .Y(n_243) );
INVx1_ASAP7_75t_L g470 ( .A(n_93), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_94), .B(n_160), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_95), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_96), .B(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_97), .A2(n_143), .B(n_241), .Y(n_240) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_98), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g517 ( .A(n_98), .B(n_174), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_99), .B(n_160), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_100), .A2(n_492), .B(n_493), .C(n_496), .Y(n_491) );
BUFx2_ASAP7_75t_L g111 ( .A(n_101), .Y(n_111) );
BUFx2_ASAP7_75t_SL g444 ( .A(n_101), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_102), .A2(n_143), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_103), .B(n_150), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_789), .B(n_797), .Y(n_104) );
OA22x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_112), .B1(n_441), .B2(n_445), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI21x1_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_123), .B(n_438), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g440 ( .A(n_116), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
OR2x6_ASAP7_75t_SL g774 ( .A(n_117), .B(n_118), .Y(n_774) );
AND2x6_ASAP7_75t_SL g778 ( .A(n_117), .B(n_119), .Y(n_778) );
OR2x2_ASAP7_75t_L g781 ( .A(n_117), .B(n_119), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
XNOR2x2_ASAP7_75t_SL g124 ( .A(n_125), .B(n_131), .Y(n_124) );
INVx1_ASAP7_75t_L g129 ( .A(n_126), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_131), .A2(n_453), .B1(n_772), .B2(n_775), .Y(n_452) );
INVx3_ASAP7_75t_L g786 ( .A(n_131), .Y(n_786) );
NAND4xp75_ASAP7_75t_L g131 ( .A(n_132), .B(n_348), .C(n_388), .D(n_417), .Y(n_131) );
NOR2x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_310), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_267), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_200), .B(n_221), .Y(n_134) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_136), .B(n_163), .Y(n_135) );
AND2x4_ASAP7_75t_L g266 ( .A(n_136), .B(n_226), .Y(n_266) );
INVx1_ASAP7_75t_SL g319 ( .A(n_136), .Y(n_319) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_136), .A2(n_355), .B(n_358), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_SL g358 ( .A1(n_136), .A2(n_359), .B(n_360), .C(n_361), .Y(n_358) );
NAND2x1_ASAP7_75t_L g399 ( .A(n_136), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_136), .B(n_360), .Y(n_421) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g224 ( .A(n_137), .Y(n_224) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_137), .Y(n_298) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_142), .B(n_162), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_138), .A2(n_206), .B(n_207), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_138), .Y(n_219) );
OA21x2_ASAP7_75t_L g308 ( .A1(n_138), .A2(n_142), .B(n_162), .Y(n_308) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x4_ASAP7_75t_L g184 ( .A(n_140), .B(n_141), .Y(n_184) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
BUFx3_ASAP7_75t_L g478 ( .A(n_144), .Y(n_478) );
AND2x6_ASAP7_75t_L g158 ( .A(n_145), .B(n_151), .Y(n_158) );
INVx2_ASAP7_75t_L g468 ( .A(n_145), .Y(n_468) );
AND2x4_ASAP7_75t_L g464 ( .A(n_146), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x4_ASAP7_75t_L g160 ( .A(n_147), .B(n_153), .Y(n_160) );
INVx2_ASAP7_75t_L g472 ( .A(n_147), .Y(n_472) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_148), .Y(n_477) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_155), .Y(n_149) );
INVx1_ASAP7_75t_L g495 ( .A(n_150), .Y(n_495) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx5_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_155), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_161), .Y(n_156) );
INVxp67_ASAP7_75t_L g575 ( .A(n_158), .Y(n_575) );
INVxp67_ASAP7_75t_L g577 ( .A(n_160), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_161), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_161), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_161), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_161), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_161), .A2(n_216), .B(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_161), .A2(n_242), .B(n_243), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_161), .A2(n_259), .B(n_260), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_161), .A2(n_470), .B(n_471), .C(n_473), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_161), .A2(n_471), .B(n_485), .C(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g511 ( .A(n_161), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_161), .A2(n_471), .B(n_524), .C(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_SL g538 ( .A1(n_161), .A2(n_471), .B(n_539), .C(n_540), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_161), .A2(n_560), .B(n_561), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_161), .B(n_184), .Y(n_578) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_178), .Y(n_163) );
AND2x2_ASAP7_75t_L g290 ( .A(n_164), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g371 ( .A(n_164), .B(n_226), .Y(n_371) );
INVx1_ASAP7_75t_L g431 ( .A(n_164), .Y(n_431) );
BUFx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g275 ( .A(n_165), .B(n_191), .Y(n_275) );
AND2x2_ASAP7_75t_L g400 ( .A(n_165), .B(n_192), .Y(n_400) );
AND2x2_ASAP7_75t_L g405 ( .A(n_165), .B(n_365), .Y(n_405) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVxp67_ASAP7_75t_L g281 ( .A(n_166), .Y(n_281) );
BUFx3_ASAP7_75t_L g314 ( .A(n_166), .Y(n_314) );
AND2x2_ASAP7_75t_L g360 ( .A(n_166), .B(n_192), .Y(n_360) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_173), .B(n_177), .Y(n_166) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_167), .A2(n_173), .B(n_177), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_172), .Y(n_167) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_173), .A2(n_193), .B(n_199), .Y(n_192) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_173), .A2(n_193), .B(n_199), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_173), .A2(n_174), .B1(n_491), .B2(n_497), .Y(n_490) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_173), .A2(n_520), .B(n_526), .Y(n_519) );
AO21x2_ASAP7_75t_L g584 ( .A1(n_173), .A2(n_520), .B(n_526), .Y(n_584) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_175), .B(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx4f_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
AND2x2_ASAP7_75t_L g345 ( .A(n_178), .B(n_223), .Y(n_345) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_191), .Y(n_178) );
AND2x4_ASAP7_75t_L g226 ( .A(n_179), .B(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g337 ( .A(n_179), .B(n_321), .Y(n_337) );
AND2x2_ASAP7_75t_SL g380 ( .A(n_179), .B(n_308), .Y(n_380) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx2_ASAP7_75t_L g316 ( .A(n_180), .Y(n_316) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g277 ( .A(n_181), .Y(n_277) );
OAI21x1_ASAP7_75t_SL g181 ( .A1(n_182), .A2(n_185), .B(n_189), .Y(n_181) );
INVx1_ASAP7_75t_L g190 ( .A(n_183), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_184), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_SL g238 ( .A(n_184), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_184), .A2(n_256), .B(n_257), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_184), .A2(n_463), .B(n_474), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_191), .B(n_277), .Y(n_280) );
AND2x2_ASAP7_75t_L g365 ( .A(n_191), .B(n_308), .Y(n_365) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g362 ( .A(n_192), .B(n_224), .Y(n_362) );
AND2x2_ASAP7_75t_L g382 ( .A(n_192), .B(n_308), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_194), .B(n_198), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_200), .B(n_271), .Y(n_300) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_200), .A2(n_394), .B1(n_395), .B2(n_396), .C(n_398), .Y(n_393) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OAI332xp33_ASAP7_75t_L g427 ( .A1(n_201), .A2(n_287), .A3(n_294), .B1(n_353), .B2(n_428), .B3(n_429), .C1(n_430), .C2(n_432), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g201 ( .A(n_202), .B(n_211), .Y(n_201) );
AND2x2_ASAP7_75t_L g232 ( .A(n_202), .B(n_212), .Y(n_232) );
AND2x2_ASAP7_75t_L g249 ( .A(n_202), .B(n_250), .Y(n_249) );
INVx4_ASAP7_75t_L g262 ( .A(n_202), .Y(n_262) );
AND2x2_ASAP7_75t_SL g322 ( .A(n_202), .B(n_263), .Y(n_322) );
INVx5_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2x1_ASAP7_75t_SL g284 ( .A(n_203), .B(n_250), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_203), .B(n_211), .Y(n_288) );
AND2x2_ASAP7_75t_L g295 ( .A(n_203), .B(n_212), .Y(n_295) );
BUFx2_ASAP7_75t_L g330 ( .A(n_203), .Y(n_330) );
AND2x2_ASAP7_75t_L g385 ( .A(n_203), .B(n_253), .Y(n_385) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
OR2x2_ASAP7_75t_L g252 ( .A(n_211), .B(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g263 ( .A(n_211), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g303 ( .A(n_211), .Y(n_303) );
AND2x2_ASAP7_75t_L g373 ( .A(n_211), .B(n_272), .Y(n_373) );
AND2x2_ASAP7_75t_L g386 ( .A(n_211), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_211), .B(n_387), .Y(n_404) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_212), .Y(n_270) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_219), .B(n_220), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_218), .Y(n_213) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_219), .A2(n_535), .B(n_541), .Y(n_534) );
OAI32xp33_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_228), .A3(n_233), .B1(n_247), .B2(n_265), .Y(n_221) );
INVx2_ASAP7_75t_L g331 ( .A(n_222), .Y(n_331) );
OR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_225), .Y(n_222) );
INVx1_ASAP7_75t_L g342 ( .A(n_223), .Y(n_342) );
BUFx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x4_ASAP7_75t_L g276 ( .A(n_224), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g409 ( .A(n_224), .B(n_314), .Y(n_409) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g321 ( .A(n_227), .Y(n_321) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
INVx2_ASAP7_75t_L g309 ( .A(n_230), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_230), .B(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x4_ASAP7_75t_SL g320 ( .A(n_231), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g397 ( .A(n_231), .Y(n_397) );
AND2x2_ASAP7_75t_L g415 ( .A(n_231), .B(n_277), .Y(n_415) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NOR2xp67_ASAP7_75t_SL g359 ( .A(n_234), .B(n_288), .Y(n_359) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_235), .B(n_270), .Y(n_357) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g433 ( .A(n_236), .B(n_303), .Y(n_433) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g264 ( .A(n_237), .Y(n_264) );
INVx2_ASAP7_75t_L g305 ( .A(n_237), .Y(n_305) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_245), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_238), .B(n_246), .Y(n_245) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_238), .A2(n_239), .B(n_245), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_244), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_248), .B(n_261), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_248), .B(n_307), .Y(n_392) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
AND3x2_ASAP7_75t_L g347 ( .A(n_249), .B(n_294), .C(n_303), .Y(n_347) );
AND2x2_ASAP7_75t_L g271 ( .A(n_250), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_250), .B(n_253), .Y(n_328) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g282 ( .A(n_252), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g272 ( .A(n_253), .Y(n_272) );
INVx1_ASAP7_75t_L g287 ( .A(n_253), .Y(n_287) );
BUFx3_ASAP7_75t_L g294 ( .A(n_253), .Y(n_294) );
AND2x2_ASAP7_75t_L g304 ( .A(n_253), .B(n_305), .Y(n_304) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_254), .A2(n_483), .B(n_487), .Y(n_482) );
INVx2_ASAP7_75t_SL g508 ( .A(n_254), .Y(n_508) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AND2x4_ASAP7_75t_L g313 ( .A(n_262), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_262), .B(n_272), .Y(n_356) );
AND2x2_ASAP7_75t_L g312 ( .A(n_263), .B(n_287), .Y(n_312) );
INVx2_ASAP7_75t_L g339 ( .A(n_263), .Y(n_339) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
AOI211xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_273), .B(n_278), .C(n_299), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g419 ( .A1(n_268), .A2(n_395), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_271), .B(n_330), .Y(n_329) );
AOI211xp5_ASAP7_75t_SL g349 ( .A1(n_271), .A2(n_350), .B(n_354), .C(n_363), .Y(n_349) );
AND2x2_ASAP7_75t_L g335 ( .A(n_272), .B(n_295), .Y(n_335) );
OR2x2_ASAP7_75t_L g338 ( .A(n_272), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_275), .B(n_380), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_276), .B(n_321), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_276), .A2(n_302), .B1(n_382), .B2(n_385), .C(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g307 ( .A(n_277), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g353 ( .A(n_277), .B(n_308), .Y(n_353) );
OAI221xp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_282), .B1(n_285), .B2(n_289), .C(n_292), .Y(n_278) );
AND2x2_ASAP7_75t_L g424 ( .A(n_279), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g291 ( .A(n_280), .Y(n_291) );
INVx1_ASAP7_75t_L g377 ( .A(n_281), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_282), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g296 ( .A(n_284), .B(n_287), .Y(n_296) );
AND2x2_ASAP7_75t_L g372 ( .A(n_284), .B(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g297 ( .A(n_291), .B(n_298), .Y(n_297) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_296), .B(n_297), .Y(n_292) );
INVx1_ASAP7_75t_L g416 ( .A(n_293), .Y(n_416) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g395 ( .A(n_294), .B(n_322), .Y(n_395) );
AND2x2_ASAP7_75t_SL g368 ( .A(n_295), .B(n_304), .Y(n_368) );
AOI21xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B(n_306), .Y(n_299) );
OAI22xp33_ASAP7_75t_L g336 ( .A1(n_300), .A2(n_334), .B1(n_337), .B2(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g406 ( .A(n_300), .Y(n_406) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g326 ( .A(n_303), .Y(n_326) );
INVx1_ASAP7_75t_L g387 ( .A(n_305), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_307), .B(n_309), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_307), .B(n_377), .Y(n_428) );
AND2x2_ASAP7_75t_L g396 ( .A(n_308), .B(n_397), .Y(n_396) );
OAI211xp5_ASAP7_75t_L g389 ( .A1(n_309), .A2(n_390), .B(n_393), .C(n_401), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_332), .Y(n_310) );
AOI322xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .A3(n_315), .B1(n_317), .B2(n_322), .C1(n_323), .C2(n_331), .Y(n_311) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_313), .Y(n_429) );
AND2x2_ASAP7_75t_L g379 ( .A(n_314), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g413 ( .A(n_314), .Y(n_413) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_SL g364 ( .A(n_316), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_SL g370 ( .A(n_316), .B(n_362), .Y(n_370) );
AND2x2_ASAP7_75t_L g394 ( .A(n_316), .B(n_360), .Y(n_394) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g366 ( .A(n_320), .Y(n_366) );
NAND2xp33_ASAP7_75t_SL g323 ( .A(n_324), .B(n_329), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI221xp5_ASAP7_75t_SL g369 ( .A1(n_325), .A2(n_370), .B1(n_371), .B2(n_372), .C(n_374), .Y(n_369) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g436 ( .A(n_328), .Y(n_436) );
AOI211xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B(n_336), .C(n_340), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g411 ( .A(n_335), .Y(n_411) );
INVx1_ASAP7_75t_L g343 ( .A(n_337), .Y(n_343) );
OR2x2_ASAP7_75t_L g430 ( .A(n_337), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_SL g426 ( .A(n_338), .Y(n_426) );
AOI21xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B(n_346), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_342), .B(n_360), .Y(n_437) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_369), .Y(n_348) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_352), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
OR2x2_ASAP7_75t_L g403 ( .A(n_356), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI21xp33_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_366), .B(n_367), .Y(n_363) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
AOI31xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .A3(n_381), .B(n_383), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_380), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B1(n_406), .B2(n_407), .C(n_410), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_414), .B2(n_416), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g414 ( .A(n_415), .Y(n_414) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_427), .C(n_434), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_426), .Y(n_422) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_438), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
CKINVDCx11_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
CKINVDCx8_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_446), .B(n_782), .Y(n_445) );
INVx1_ASAP7_75t_L g783 ( .A(n_447), .Y(n_783) );
INVx2_ASAP7_75t_L g788 ( .A(n_453), .Y(n_788) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND3x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_662), .C(n_727), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_616), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_563), .B(n_589), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_527), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_479), .Y(n_458) );
AOI21xp33_ASAP7_75t_L g663 ( .A1(n_459), .A2(n_664), .B(n_675), .Y(n_663) );
AND2x2_ASAP7_75t_SL g698 ( .A(n_459), .B(n_605), .Y(n_698) );
AND2x2_ASAP7_75t_L g713 ( .A(n_459), .B(n_714), .Y(n_713) );
OR2x6_ASAP7_75t_L g723 ( .A(n_459), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g725 ( .A(n_459), .B(n_715), .Y(n_725) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g599 ( .A(n_460), .Y(n_599) );
AND2x2_ASAP7_75t_L g612 ( .A(n_460), .B(n_613), .Y(n_612) );
INVx4_ASAP7_75t_L g631 ( .A(n_460), .Y(n_631) );
AND2x2_ASAP7_75t_L g634 ( .A(n_460), .B(n_552), .Y(n_634) );
NOR2x1_ASAP7_75t_SL g637 ( .A(n_460), .B(n_567), .Y(n_637) );
AND2x4_ASAP7_75t_L g649 ( .A(n_460), .B(n_647), .Y(n_649) );
OR2x2_ASAP7_75t_L g659 ( .A(n_460), .B(n_534), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_460), .B(n_671), .Y(n_676) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVxp67_ASAP7_75t_L g502 ( .A(n_464), .Y(n_502) );
NOR2x1p5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g515 ( .A(n_467), .Y(n_515) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR2x6_ASAP7_75t_L g471 ( .A(n_468), .B(n_472), .Y(n_471) );
INVxp67_ASAP7_75t_L g492 ( .A(n_471), .Y(n_492) );
INVx2_ASAP7_75t_L g562 ( .A(n_471), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_471), .A2(n_495), .B1(n_571), .B2(n_572), .Y(n_570) );
AND2x2_ASAP7_75t_L g476 ( .A(n_472), .B(n_477), .Y(n_476) );
INVxp33_ASAP7_75t_L g514 ( .A(n_472), .Y(n_514) );
INVx1_ASAP7_75t_L g504 ( .A(n_475), .Y(n_504) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
INVx1_ASAP7_75t_L g555 ( .A(n_476), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_478), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_479), .A2(n_605), .B1(n_700), .B2(n_701), .Y(n_699) );
INVx1_ASAP7_75t_SL g743 ( .A(n_479), .Y(n_743) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_505), .Y(n_479) );
INVx2_ASAP7_75t_L g674 ( .A(n_480), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_480), .B(n_620), .Y(n_746) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_488), .Y(n_480) );
BUFx3_ASAP7_75t_L g592 ( .A(n_481), .Y(n_592) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g585 ( .A(n_482), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_482), .B(n_507), .Y(n_607) );
AND2x4_ASAP7_75t_L g624 ( .A(n_482), .B(n_625), .Y(n_624) );
INVxp67_ASAP7_75t_L g640 ( .A(n_482), .Y(n_640) );
INVx2_ASAP7_75t_L g697 ( .A(n_482), .Y(n_697) );
AND2x2_ASAP7_75t_L g615 ( .A(n_488), .B(n_581), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g661 ( .A(n_488), .B(n_584), .Y(n_661) );
AND2x2_ASAP7_75t_L g680 ( .A(n_488), .B(n_584), .Y(n_680) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g544 ( .A(n_489), .Y(n_544) );
INVx1_ASAP7_75t_L g623 ( .A(n_489), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_489), .B(n_519), .Y(n_642) );
AND2x4_ASAP7_75t_L g696 ( .A(n_489), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_498), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g655 ( .A(n_505), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_505), .B(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_518), .Y(n_505) );
AND2x2_ASAP7_75t_L g639 ( .A(n_506), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g679 ( .A(n_506), .Y(n_679) );
AND2x2_ASAP7_75t_L g684 ( .A(n_506), .B(n_584), .Y(n_684) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_507), .B(n_519), .Y(n_546) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_517), .Y(n_507) );
AO21x2_ASAP7_75t_L g581 ( .A1(n_508), .A2(n_509), .B(n_517), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_510), .B(n_516), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g620 ( .A(n_518), .Y(n_620) );
NAND2x1p5_ASAP7_75t_L g738 ( .A(n_518), .B(n_592), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_518), .B(n_544), .Y(n_759) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_519), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
OAI21xp33_ASAP7_75t_SL g527 ( .A1(n_528), .A2(n_542), .B(n_547), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_530), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g597 ( .A(n_531), .Y(n_597) );
AND2x2_ASAP7_75t_L g611 ( .A(n_531), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g645 ( .A(n_531), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g711 ( .A(n_531), .B(n_629), .Y(n_711) );
NOR3xp33_ASAP7_75t_L g757 ( .A(n_531), .B(n_758), .C(n_759), .Y(n_757) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_532), .Y(n_588) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g604 ( .A(n_534), .Y(n_604) );
AND2x2_ASAP7_75t_L g610 ( .A(n_534), .B(n_567), .Y(n_610) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_534), .Y(n_621) );
AND2x2_ASAP7_75t_L g666 ( .A(n_534), .B(n_566), .Y(n_666) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_534), .Y(n_689) );
INVx1_ASAP7_75t_L g706 ( .A(n_534), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g748 ( .A(n_542), .Y(n_748) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_543), .B(n_619), .Y(n_720) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g582 ( .A(n_544), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI211x1_ASAP7_75t_L g616 ( .A1(n_548), .A2(n_617), .B(n_626), .C(n_643), .Y(n_616) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_SL g609 ( .A(n_549), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g669 ( .A(n_549), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g605 ( .A(n_551), .B(n_566), .Y(n_605) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g565 ( .A(n_552), .B(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_552), .Y(n_630) );
INVx1_ASAP7_75t_L g647 ( .A(n_552), .Y(n_647) );
AND2x2_ASAP7_75t_L g715 ( .A(n_552), .B(n_567), .Y(n_715) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_558), .Y(n_552) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .C(n_557), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_579), .B(n_586), .Y(n_563) );
NOR2x1_ASAP7_75t_L g734 ( .A(n_564), .B(n_631), .Y(n_734) );
INVx2_ASAP7_75t_L g766 ( .A(n_564), .Y(n_766) );
INVx4_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g598 ( .A(n_565), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g671 ( .A(n_566), .Y(n_671) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g613 ( .A(n_567), .Y(n_613) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .B(n_578), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
OR2x2_ASAP7_75t_L g673 ( .A(n_580), .B(n_674), .Y(n_673) );
NAND2x1_ASAP7_75t_SL g695 ( .A(n_580), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_L g595 ( .A(n_581), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g625 ( .A(n_581), .Y(n_625) );
INVx1_ASAP7_75t_L g749 ( .A(n_582), .Y(n_749) );
AND2x2_ASAP7_75t_L g614 ( .A(n_583), .B(n_615), .Y(n_614) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx2_ASAP7_75t_L g596 ( .A(n_584), .Y(n_596) );
INVxp33_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g653 ( .A(n_588), .B(n_646), .Y(n_653) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_593), .B(n_600), .C(n_608), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g677 ( .A(n_591), .B(n_678), .Y(n_677) );
NOR2xp67_ASAP7_75t_SL g682 ( .A(n_591), .B(n_683), .Y(n_682) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_592), .B(n_679), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_598), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
AND2x2_ASAP7_75t_L g726 ( .A(n_595), .B(n_696), .Y(n_726) );
AOI222xp33_ASAP7_75t_L g744 ( .A1(n_598), .A2(n_745), .B1(n_747), .B2(n_750), .C1(n_751), .C2(n_754), .Y(n_744) );
INVx1_ASAP7_75t_L g708 ( .A(n_599), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_606), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_604), .Y(n_635) );
AND2x4_ASAP7_75t_SL g670 ( .A(n_604), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g724 ( .A(n_605), .Y(n_724) );
AND2x2_ASAP7_75t_L g769 ( .A(n_605), .B(n_621), .Y(n_769) );
AND2x2_ASAP7_75t_L g650 ( .A(n_606), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g763 ( .A(n_607), .B(n_642), .Y(n_763) );
OAI21xp33_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_611), .B(n_614), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_609), .A2(n_629), .B(n_670), .Y(n_730) );
AND2x2_ASAP7_75t_L g754 ( .A(n_610), .B(n_631), .Y(n_754) );
NOR2xp33_ASAP7_75t_SL g764 ( .A(n_610), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g702 ( .A(n_613), .Y(n_702) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_613), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g737 ( .A(n_615), .Y(n_737) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_622), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AND2x2_ASAP7_75t_L g740 ( .A(n_620), .B(n_624), .Y(n_740) );
BUFx2_ASAP7_75t_L g628 ( .A(n_621), .Y(n_628) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g651 ( .A(n_623), .Y(n_651) );
INVx2_ASAP7_75t_L g657 ( .A(n_623), .Y(n_657) );
AND2x2_ASAP7_75t_L g693 ( .A(n_623), .B(n_684), .Y(n_693) );
AND2x4_ASAP7_75t_L g660 ( .A(n_624), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g700 ( .A(n_624), .B(n_657), .Y(n_700) );
AND2x2_ASAP7_75t_L g751 ( .A(n_624), .B(n_752), .Y(n_751) );
AOI31xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_632), .A3(n_636), .B(n_638), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
AND2x2_ASAP7_75t_L g648 ( .A(n_628), .B(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_SL g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x4_ASAP7_75t_L g646 ( .A(n_631), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_634), .A2(n_686), .B1(n_717), .B2(n_720), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_634), .B(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g771 ( .A(n_634), .B(n_687), .Y(n_771) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g686 ( .A(n_637), .B(n_687), .Y(n_686) );
NAND2x1p5_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
AND2x2_ASAP7_75t_L g709 ( .A(n_639), .B(n_680), .Y(n_709) );
INVx1_ASAP7_75t_L g719 ( .A(n_641), .Y(n_719) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_652), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_648), .B(n_650), .Y(n_644) );
INVx1_ASAP7_75t_L g742 ( .A(n_645), .Y(n_742) );
AND2x2_ASAP7_75t_L g750 ( .A(n_646), .B(n_702), .Y(n_750) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_646), .Y(n_756) );
AND2x2_ASAP7_75t_L g701 ( .A(n_649), .B(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B1(n_658), .B2(n_660), .Y(n_652) );
NOR2xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_656), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_655), .A2(n_674), .B1(n_768), .B2(n_770), .Y(n_767) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g667 ( .A(n_660), .Y(n_667) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_690), .Y(n_662) );
OAI21xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B(n_668), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
OAI21xp33_ASAP7_75t_L g668 ( .A1(n_666), .A2(n_669), .B(n_672), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_669), .A2(n_693), .B1(n_694), .B2(n_698), .Y(n_692) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_681), .B2(n_685), .Y(n_675) );
INVx1_ASAP7_75t_L g710 ( .A(n_678), .Y(n_710) );
NAND2x1p5_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g690 ( .A(n_691), .B(n_703), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_699), .Y(n_691) );
INVx2_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
NAND2xp33_ASAP7_75t_SL g745 ( .A(n_695), .B(n_746), .Y(n_745) );
INVx3_ASAP7_75t_L g718 ( .A(n_696), .Y(n_718) );
INVx3_ASAP7_75t_L g732 ( .A(n_700), .Y(n_732) );
INVxp67_ASAP7_75t_L g761 ( .A(n_701), .Y(n_761) );
NAND4xp25_ASAP7_75t_L g703 ( .A(n_704), .B(n_712), .C(n_716), .D(n_721), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
AND2x2_ASAP7_75t_L g714 ( .A(n_706), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g762 ( .A(n_710), .Y(n_762) );
NAND2xp33_ASAP7_75t_SL g717 ( .A(n_718), .B(n_719), .Y(n_717) );
OAI21xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_725), .B(n_726), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AND3x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_744), .C(n_755), .Y(n_727) );
AOI221x1_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B1(n_733), .B2(n_735), .C(n_741), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp33_ASAP7_75t_SL g735 ( .A(n_736), .B(n_739), .Y(n_735) );
OR2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
NAND2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI211xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B(n_760), .C(n_767), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_760) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_773), .Y(n_787) );
CKINVDCx11_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
CKINVDCx6p67_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
CKINVDCx11_ASAP7_75t_R g785 ( .A(n_776), .Y(n_785) );
INVx3_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
BUFx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
OAI22x1_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_786), .B1(n_787), .B2(n_788), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g800 ( .A(n_790), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_SL g791 ( .A(n_792), .B(n_793), .Y(n_791) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
endmodule