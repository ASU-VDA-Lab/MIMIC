module fake_jpeg_4961_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx24_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_0),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_41),
.C(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_60),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_20),
.B1(n_19),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_20),
.B1(n_19),
.B2(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_19),
.B1(n_37),
.B2(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_61),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_20),
.B1(n_28),
.B2(n_21),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_24),
.B1(n_23),
.B2(n_25),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AND2x4_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_64),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_39),
.B(n_41),
.C(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_28),
.B1(n_23),
.B2(n_27),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_44),
.B1(n_49),
.B2(n_25),
.Y(n_90)
);

AOI32xp33_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_32),
.A3(n_37),
.B1(n_25),
.B2(n_31),
.Y(n_78)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_78),
.B(n_82),
.CI(n_32),
.CON(n_109),
.SN(n_109)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_33),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_84),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g85 ( 
.A(n_58),
.Y(n_85)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_16),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_108),
.Y(n_117)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_98),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_44),
.C(n_52),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_62),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_0),
.B(n_1),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_101),
.B(n_96),
.Y(n_118)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_105),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_109),
.Y(n_112)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_73),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_16),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_82),
.B1(n_66),
.B2(n_76),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_134),
.B1(n_32),
.B2(n_29),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_79),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_129),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_75),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_87),
.B1(n_98),
.B2(n_105),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_130),
.B(n_29),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_107),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_109),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_75),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_26),
.Y(n_158)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_133),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_80),
.B(n_69),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_132),
.CI(n_93),
.CON(n_141),
.SN(n_141)
);

BUFx2_ASAP7_75t_SL g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_67),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_65),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_62),
.B(n_73),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_29),
.C(n_26),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_110),
.A2(n_84),
.B1(n_74),
.B2(n_32),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_109),
.B1(n_103),
.B2(n_102),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_141),
.B(n_151),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_156),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_15),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_147),
.C(n_152),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_74),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_134),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_130),
.B(n_116),
.C(n_133),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_124),
.B1(n_113),
.B2(n_120),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_29),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g183 ( 
.A(n_153),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_115),
.A2(n_26),
.B1(n_22),
.B2(n_18),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_2),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_161),
.B(n_118),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_2),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_160),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_2),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_177),
.B1(n_156),
.B2(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_114),
.C(n_129),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_174),
.C(n_175),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_142),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_152),
.C(n_161),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_125),
.C(n_120),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_179),
.C(n_181),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_26),
.Y(n_177)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_150),
.B1(n_144),
.B2(n_138),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_137),
.B1(n_158),
.B2(n_141),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_22),
.C(n_18),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_22),
.B(n_18),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_180),
.Y(n_185)
);

NAND2x1_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_22),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_174),
.C(n_164),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_200),
.C(n_201),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_145),
.B1(n_141),
.B2(n_136),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_163),
.B(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_199),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_202),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_18),
.B1(n_5),
.B2(n_6),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_14),
.C(n_5),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_4),
.C(n_5),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_170),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_208),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_169),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_182),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_214),
.C(n_8),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_169),
.C(n_165),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_187),
.A2(n_168),
.B(n_162),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_216),
.A2(n_207),
.B(n_209),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_203),
.B(n_205),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_206),
.A2(n_197),
.B1(n_202),
.B2(n_195),
.Y(n_218)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_185),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_220),
.B(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_198),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_186),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_227),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_212),
.B(n_177),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_207),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_201),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_225),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_4),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_8),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_209),
.CI(n_213),
.CON(n_228),
.SN(n_228)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_235),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_233),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_219),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_240),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_203),
.Y(n_240)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_243),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_222),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_231),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_9),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_230),
.B1(n_235),
.B2(n_219),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_237),
.B1(n_241),
.B2(n_9),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_8),
.CI(n_9),
.CON(n_246),
.SN(n_246)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_10),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_248),
.C(n_247),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_250),
.A2(n_251),
.B(n_246),
.C(n_248),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_252),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_254),
.B(n_253),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_255),
.B(n_10),
.Y(n_256)
);


endmodule