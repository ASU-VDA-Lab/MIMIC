module fake_netlist_1_5496_n_547 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_547);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_547;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g76 ( .A(n_19), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_22), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_22), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_74), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_17), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_41), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_61), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_15), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_29), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_69), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_47), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_55), .Y(n_87) );
NOR2xp33_ASAP7_75t_L g88 ( .A(n_70), .B(n_17), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_58), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_24), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_18), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_23), .Y(n_92) );
INVxp67_ASAP7_75t_L g93 ( .A(n_2), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_28), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_18), .Y(n_95) );
CKINVDCx14_ASAP7_75t_R g96 ( .A(n_50), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_26), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_8), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_31), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_25), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_40), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_16), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_19), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_23), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_73), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_7), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_46), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_13), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_57), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g111 ( .A1(n_90), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_101), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_90), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_101), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
NOR2xp33_ASAP7_75t_R g116 ( .A(n_96), .B(n_37), .Y(n_116) );
INVx6_ASAP7_75t_L g117 ( .A(n_110), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_101), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_79), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_77), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_78), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_79), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_80), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_82), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_102), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_82), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_77), .B(n_3), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_84), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_119), .Y(n_135) );
NOR2xp33_ASAP7_75t_SL g136 ( .A(n_132), .B(n_99), .Y(n_136) );
NOR2xp33_ASAP7_75t_SL g137 ( .A(n_132), .B(n_86), .Y(n_137) );
INVx2_ASAP7_75t_SL g138 ( .A(n_133), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_119), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_133), .B(n_86), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_117), .B(n_87), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_119), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_129), .B(n_83), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_119), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_117), .B(n_87), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_112), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_114), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_129), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_129), .B(n_89), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_122), .Y(n_152) );
INVxp33_ASAP7_75t_L g153 ( .A(n_121), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_114), .Y(n_154) );
OR2x6_ASAP7_75t_L g155 ( .A(n_117), .B(n_83), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_134), .B(n_89), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_121), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_117), .B(n_91), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_118), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_134), .B(n_94), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_118), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_138), .B(n_123), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_151), .A2(n_123), .B1(n_98), .B2(n_111), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_153), .B(n_122), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_138), .B(n_124), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_138), .B(n_124), .Y(n_167) );
OR2x6_ASAP7_75t_L g168 ( .A(n_155), .B(n_93), .Y(n_168) );
NOR2x1_ASAP7_75t_L g169 ( .A(n_157), .B(n_125), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_157), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_155), .Y(n_172) );
CKINVDCx8_ASAP7_75t_R g173 ( .A(n_155), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_142), .B(n_125), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_136), .B(n_116), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_155), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_155), .B(n_113), .Y(n_178) );
INVx1_ASAP7_75t_SL g179 ( .A(n_155), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_137), .A2(n_115), .B(n_130), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_141), .A2(n_130), .B(n_128), .C(n_126), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_158), .B(n_126), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_151), .A2(n_100), .B1(n_93), .B2(n_76), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_136), .B(n_128), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_152), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_150), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_160), .A2(n_115), .B(n_131), .C(n_120), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_151), .A2(n_144), .B1(n_158), .B2(n_146), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_137), .B(n_94), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_150), .A2(n_144), .B1(n_158), .B2(n_142), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_144), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_147), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_146), .B(n_131), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_181), .A2(n_160), .B(n_144), .C(n_141), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_194), .A2(n_190), .B(n_195), .C(n_174), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_197), .A2(n_156), .B(n_144), .C(n_76), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_183), .A2(n_156), .B(n_159), .C(n_148), .Y(n_202) );
INVx5_ASAP7_75t_L g203 ( .A(n_168), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_173), .A2(n_150), .B1(n_159), .B2(n_161), .Y(n_204) );
AO22x1_ASAP7_75t_L g205 ( .A1(n_171), .A2(n_151), .B1(n_127), .B2(n_91), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_187), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_168), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_162), .A2(n_161), .B(n_149), .C(n_148), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_187), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_168), .Y(n_210) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_168), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_196), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_178), .B(n_151), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_189), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_171), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_178), .B(n_151), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_189), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_165), .A2(n_149), .B(n_147), .C(n_154), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_191), .B(n_151), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_182), .Y(n_220) );
BUFx2_ASAP7_75t_L g221 ( .A(n_172), .Y(n_221) );
OR2x6_ASAP7_75t_SL g222 ( .A(n_172), .B(n_151), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_166), .A2(n_147), .B(n_135), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_177), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_167), .A2(n_186), .B(n_193), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_173), .B(n_151), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_185), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_179), .B(n_154), .Y(n_228) );
INVx4_ASAP7_75t_L g229 ( .A(n_177), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_184), .B(n_154), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_196), .A2(n_135), .B(n_145), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_163), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_213), .B(n_178), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_213), .B(n_164), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_213), .A2(n_169), .B1(n_163), .B2(n_188), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_212), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_203), .A2(n_154), .B1(n_106), .B2(n_103), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_216), .A2(n_163), .B1(n_176), .B2(n_106), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_206), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_200), .Y(n_240) );
AOI211x1_ASAP7_75t_L g241 ( .A1(n_230), .A2(n_180), .B(n_107), .C(n_105), .Y(n_241) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_198), .A2(n_107), .A3(n_105), .B(n_97), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_209), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_216), .B(n_163), .Y(n_244) );
AOI221xp5_ASAP7_75t_L g245 ( .A1(n_201), .A2(n_108), .B1(n_92), .B2(n_95), .C(n_103), .Y(n_245) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_198), .A2(n_192), .B(n_175), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_216), .B(n_109), .Y(n_247) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_225), .A2(n_97), .B(n_145), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_214), .B(n_109), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_224), .B(n_108), .Y(n_250) );
OAI21x1_ASAP7_75t_SL g251 ( .A1(n_207), .A2(n_92), .B(n_95), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_212), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_221), .B(n_104), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_200), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_200), .Y(n_255) );
CKINVDCx11_ASAP7_75t_R g256 ( .A(n_222), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_215), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_207), .A2(n_104), .B1(n_88), .B2(n_143), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_203), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_240), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_246), .A2(n_218), .B(n_208), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_256), .A2(n_207), .B1(n_221), .B2(n_229), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_233), .B(n_205), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_237), .A2(n_203), .B1(n_222), .B2(n_210), .Y(n_264) );
AO21x1_ASAP7_75t_L g265 ( .A1(n_246), .A2(n_199), .B(n_202), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_256), .A2(n_224), .B1(n_229), .B2(n_203), .Y(n_266) );
OAI221xp5_ASAP7_75t_L g267 ( .A1(n_245), .A2(n_219), .B1(n_218), .B2(n_204), .C(n_210), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_239), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_239), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_236), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_248), .A2(n_223), .B(n_231), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_234), .B(n_224), .Y(n_272) );
AOI22xp33_ASAP7_75t_SL g273 ( .A1(n_251), .A2(n_203), .B1(n_229), .B2(n_211), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_236), .A2(n_228), .B(n_232), .Y(n_274) );
NAND3xp33_ASAP7_75t_L g275 ( .A(n_241), .B(n_228), .C(n_232), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g276 ( .A1(n_245), .A2(n_217), .B1(n_227), .B2(n_220), .C(n_226), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_257), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_237), .A2(n_226), .B1(n_232), .B2(n_200), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_259), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_233), .B(n_232), .Y(n_280) );
AOI22xp33_ASAP7_75t_SL g281 ( .A1(n_251), .A2(n_232), .B1(n_200), .B2(n_6), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_270), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_270), .B(n_242), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_268), .B(n_242), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_268), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_269), .B(n_243), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_270), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_260), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_265), .B(n_242), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_265), .B(n_243), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_260), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_272), .B(n_234), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_280), .B(n_242), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_260), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_271), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_275), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_278), .B(n_242), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_261), .B(n_242), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_263), .B(n_242), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_276), .B(n_242), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_275), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_294), .A2(n_264), .B1(n_278), .B2(n_250), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_283), .B(n_236), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_287), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_285), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_287), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_285), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_287), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_290), .B(n_241), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_290), .B(n_249), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_282), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_283), .B(n_254), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_299), .B(n_252), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_299), .B(n_252), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_299), .B(n_252), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_282), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_294), .A2(n_264), .B1(n_250), .B2(n_267), .Y(n_322) );
AOI211xp5_ASAP7_75t_L g323 ( .A1(n_291), .A2(n_277), .B(n_253), .C(n_259), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_297), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_284), .B(n_249), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_297), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_283), .B(n_248), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_291), .B(n_248), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_303), .A2(n_279), .B1(n_233), .B2(n_281), .Y(n_329) );
OAI33xp33_ASAP7_75t_L g330 ( .A1(n_284), .A2(n_253), .A3(n_247), .B1(n_139), .B2(n_143), .B3(n_9), .Y(n_330) );
OAI33xp33_ASAP7_75t_L g331 ( .A1(n_300), .A2(n_253), .A3(n_247), .B1(n_139), .B2(n_8), .B3(n_9), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_292), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_282), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_292), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_291), .B(n_255), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_319), .B(n_295), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_336), .B(n_302), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_319), .B(n_300), .Y(n_339) );
NAND3xp33_ASAP7_75t_SL g340 ( .A(n_323), .B(n_329), .C(n_322), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_317), .B(n_301), .Y(n_341) );
OAI33xp33_ASAP7_75t_L g342 ( .A1(n_309), .A2(n_301), .A3(n_303), .B1(n_286), .B2(n_304), .B3(n_298), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_317), .B(n_318), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_309), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_317), .B(n_295), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_318), .B(n_295), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_311), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_323), .B(n_286), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_336), .B(n_302), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_311), .B(n_289), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_334), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_318), .B(n_304), .Y(n_352) );
INVxp67_ASAP7_75t_L g353 ( .A(n_308), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_333), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_333), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_307), .B(n_289), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_312), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_320), .B(n_298), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_320), .B(n_302), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_327), .A2(n_289), .B1(n_288), .B2(n_293), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_320), .B(n_293), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_312), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_336), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_328), .B(n_293), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_316), .B(n_293), .Y(n_365) );
NOR3xp33_ASAP7_75t_L g366 ( .A(n_331), .B(n_273), .C(n_288), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_335), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_328), .B(n_296), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_313), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_313), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_321), .Y(n_371) );
NOR2xp33_ASAP7_75t_R g372 ( .A(n_307), .B(n_262), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_328), .B(n_296), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_325), .B(n_296), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_327), .B(n_288), .Y(n_375) );
OAI211xp5_ASAP7_75t_SL g376 ( .A1(n_322), .A2(n_258), .B(n_238), .C(n_235), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_327), .B(n_288), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_321), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_306), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_316), .B(n_288), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_306), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_325), .B(n_258), .Y(n_382) );
NAND4xp25_ASAP7_75t_L g383 ( .A(n_329), .B(n_238), .C(n_235), .D(n_266), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_364), .B(n_316), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_369), .B(n_335), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_364), .B(n_316), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_344), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_370), .B(n_305), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_343), .B(n_315), .Y(n_389) );
NOR2xp33_ASAP7_75t_R g390 ( .A(n_340), .B(n_4), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_347), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_375), .B(n_321), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_354), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_355), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_343), .B(n_315), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_355), .Y(n_397) );
AOI33xp33_ASAP7_75t_L g398 ( .A1(n_360), .A2(n_305), .A3(n_310), .B1(n_306), .B2(n_324), .B3(n_332), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_367), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_345), .B(n_310), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_345), .B(n_310), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_375), .B(n_326), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_367), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_377), .B(n_326), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_377), .B(n_326), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_379), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_348), .A2(n_314), .B1(n_326), .B2(n_332), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_339), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_339), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_381), .Y(n_410) );
NOR2xp67_ASAP7_75t_L g411 ( .A(n_371), .B(n_4), .Y(n_411) );
OAI21xp33_ASAP7_75t_L g412 ( .A1(n_372), .A2(n_314), .B(n_332), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_346), .B(n_324), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_346), .B(n_324), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_337), .B(n_5), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_368), .B(n_254), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_361), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_368), .B(n_254), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_373), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_363), .B(n_5), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_352), .B(n_7), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_358), .B(n_10), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_373), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_378), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_352), .B(n_10), .Y(n_425) );
NAND2x1p5_ASAP7_75t_L g426 ( .A(n_371), .B(n_240), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_351), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_353), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_361), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_358), .B(n_11), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_350), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_341), .B(n_11), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_359), .B(n_255), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_359), .B(n_255), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_341), .B(n_12), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_374), .B(n_12), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_411), .A2(n_356), .B1(n_371), .B2(n_382), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_408), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_412), .A2(n_430), .B1(n_422), .B2(n_388), .C(n_435), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_408), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_409), .Y(n_442) );
NAND4xp25_ASAP7_75t_L g443 ( .A(n_422), .B(n_383), .C(n_366), .D(n_376), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_428), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_400), .B(n_357), .Y(n_445) );
XOR2xp5_ASAP7_75t_L g446 ( .A(n_430), .B(n_380), .Y(n_446) );
XNOR2xp5_ASAP7_75t_L g447 ( .A(n_384), .B(n_380), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_409), .B(n_362), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_427), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_389), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_424), .B(n_342), .Y(n_451) );
NAND2xp33_ASAP7_75t_L g452 ( .A(n_390), .B(n_362), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_387), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_387), .Y(n_454) );
AOI32xp33_ASAP7_75t_L g455 ( .A1(n_413), .A2(n_365), .A3(n_349), .B1(n_338), .B2(n_331), .Y(n_455) );
INVx2_ASAP7_75t_SL g456 ( .A(n_396), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g457 ( .A1(n_398), .A2(n_365), .B(n_349), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_407), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_391), .Y(n_459) );
AOI211xp5_ASAP7_75t_L g460 ( .A1(n_432), .A2(n_330), .B(n_365), .C(n_338), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_396), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_431), .B(n_349), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_421), .A2(n_338), .B1(n_330), .B2(n_240), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_425), .A2(n_244), .B1(n_240), .B2(n_274), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_415), .A2(n_13), .B(n_14), .C(n_15), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_431), .A2(n_244), .B1(n_16), .B2(n_20), .C(n_21), .Y(n_466) );
OAI32xp33_ASAP7_75t_L g467 ( .A1(n_426), .A2(n_14), .A3(n_20), .B1(n_21), .B2(n_24), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_401), .A2(n_240), .B1(n_25), .B2(n_30), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_413), .Y(n_469) );
NAND4xp25_ASAP7_75t_L g470 ( .A(n_436), .B(n_192), .C(n_175), .D(n_170), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_391), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_420), .A2(n_240), .B1(n_170), .B2(n_33), .C(n_34), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_385), .A2(n_27), .B(n_32), .Y(n_473) );
OAI221xp5_ASAP7_75t_L g474 ( .A1(n_426), .A2(n_240), .B1(n_36), .B2(n_38), .C(n_39), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_410), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_414), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_419), .B(n_240), .Y(n_477) );
OAI21xp5_ASAP7_75t_SL g478 ( .A1(n_426), .A2(n_35), .B(n_42), .Y(n_478) );
AOI22x1_ASAP7_75t_L g479 ( .A1(n_414), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_475), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_475), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_453), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_440), .A2(n_419), .B1(n_423), .B2(n_384), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_458), .B(n_406), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_458), .B(n_406), .Y(n_485) );
AOI211x1_ASAP7_75t_L g486 ( .A1(n_443), .A2(n_423), .B(n_429), .C(n_386), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_461), .B(n_417), .Y(n_487) );
NOR4xp25_ASAP7_75t_L g488 ( .A(n_444), .B(n_403), .C(n_399), .D(n_394), .Y(n_488) );
OAI31xp33_ASAP7_75t_L g489 ( .A1(n_440), .A2(n_429), .A3(n_386), .B(n_395), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_451), .B(n_417), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_454), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_449), .B(n_393), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_452), .A2(n_404), .B1(n_402), .B2(n_405), .Y(n_493) );
XNOR2x1_ASAP7_75t_L g494 ( .A(n_446), .B(n_392), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_459), .Y(n_495) );
XNOR2x1_ASAP7_75t_L g496 ( .A(n_447), .B(n_392), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_438), .B(n_399), .Y(n_497) );
AOI221x1_ASAP7_75t_SL g498 ( .A1(n_457), .A2(n_403), .B1(n_397), .B2(n_410), .C(n_405), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_471), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_465), .A2(n_404), .B(n_402), .C(n_418), .Y(n_500) );
NOR2xp33_ASAP7_75t_SL g501 ( .A(n_478), .B(n_434), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_441), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_442), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_439), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_445), .B(n_418), .Y(n_505) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_437), .B(n_434), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_456), .B(n_433), .Y(n_507) );
NAND3xp33_ASAP7_75t_SL g508 ( .A(n_501), .B(n_455), .C(n_466), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_497), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_498), .A2(n_463), .B1(n_466), .B2(n_467), .C(n_448), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_480), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_SL g512 ( .A1(n_489), .A2(n_474), .B(n_473), .C(n_468), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_490), .B(n_460), .Y(n_513) );
OAI21xp5_ASAP7_75t_SL g514 ( .A1(n_500), .A2(n_474), .B(n_472), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_481), .Y(n_515) );
NAND3xp33_ASAP7_75t_L g516 ( .A(n_486), .B(n_472), .C(n_464), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_482), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_506), .A2(n_470), .B(n_479), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_493), .A2(n_476), .B1(n_469), .B2(n_462), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_496), .A2(n_450), .B1(n_477), .B2(n_416), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_484), .A2(n_416), .B(n_433), .C(n_51), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_483), .A2(n_48), .B1(n_49), .B2(n_52), .Y(n_522) );
XNOR2xp5_ASAP7_75t_L g523 ( .A(n_494), .B(n_53), .Y(n_523) );
AOI211xp5_ASAP7_75t_L g524 ( .A1(n_508), .A2(n_488), .B(n_484), .C(n_485), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_514), .A2(n_485), .B1(n_492), .B2(n_503), .C(n_502), .Y(n_525) );
OAI21xp5_ASAP7_75t_SL g526 ( .A1(n_518), .A2(n_505), .B(n_492), .Y(n_526) );
OAI221xp5_ASAP7_75t_SL g527 ( .A1(n_510), .A2(n_487), .B1(n_507), .B2(n_505), .C(n_504), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_517), .Y(n_528) );
OAI222xp33_ASAP7_75t_L g529 ( .A1(n_513), .A2(n_504), .B1(n_499), .B2(n_495), .C1(n_491), .C2(n_62), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_512), .A2(n_54), .B(n_56), .C(n_59), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_520), .B(n_60), .Y(n_531) );
OAI221xp5_ASAP7_75t_SL g532 ( .A1(n_510), .A2(n_63), .B1(n_64), .B2(n_65), .C(n_66), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_528), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_524), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_525), .B(n_509), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_527), .A2(n_516), .B1(n_519), .B2(n_515), .C(n_511), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g537 ( .A(n_530), .B(n_521), .C(n_522), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_533), .Y(n_538) );
AOI21xp33_ASAP7_75t_SL g539 ( .A1(n_534), .A2(n_526), .B(n_523), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_536), .A2(n_531), .B1(n_532), .B2(n_529), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_538), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_539), .A2(n_535), .B(n_537), .Y(n_542) );
OAI22xp5_ASAP7_75t_SL g543 ( .A1(n_541), .A2(n_540), .B1(n_531), .B2(n_71), .Y(n_543) );
OAI22x1_ASAP7_75t_L g544 ( .A1(n_543), .A2(n_542), .B1(n_68), .B2(n_72), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_544), .Y(n_545) );
INVxp67_ASAP7_75t_L g546 ( .A(n_545), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_546), .A2(n_67), .B(n_75), .Y(n_547) );
endmodule