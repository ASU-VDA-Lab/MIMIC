module fake_netlist_1_8456_n_939 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_113, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_939);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_113;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_939;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_227;
wire n_163;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_245;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx10_ASAP7_75t_L g114 ( .A(n_106), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_61), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_90), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_0), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_30), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_91), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_20), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_46), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_58), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_42), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_18), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_2), .Y(n_125) );
BUFx10_ASAP7_75t_L g126 ( .A(n_72), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_11), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_55), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_77), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_97), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_99), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_10), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_85), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_9), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_10), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g136 ( .A(n_70), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_2), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_14), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_44), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_95), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_6), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_34), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_50), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_18), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_0), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_56), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_48), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_102), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_13), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_59), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g151 ( .A(n_100), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_60), .Y(n_152) );
BUFx10_ASAP7_75t_L g153 ( .A(n_6), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_34), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_53), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_44), .Y(n_156) );
INVx1_ASAP7_75t_SL g157 ( .A(n_88), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_68), .Y(n_158) );
INVx2_ASAP7_75t_SL g159 ( .A(n_114), .Y(n_159) );
INVx5_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_136), .B(n_151), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_152), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_123), .B(n_1), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_153), .B(n_1), .Y(n_165) );
BUFx12f_ASAP7_75t_L g166 ( .A(n_114), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_132), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_132), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_123), .B(n_3), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_117), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_120), .B(n_3), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_143), .B(n_4), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_147), .B(n_4), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_150), .B(n_5), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_114), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_126), .Y(n_182) );
BUFx10_ASAP7_75t_L g183 ( .A(n_159), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_161), .A2(n_118), .B1(n_117), .B2(n_156), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g185 ( .A1(n_174), .A2(n_118), .B1(n_156), .B2(n_145), .Y(n_185) );
AO22x2_ASAP7_75t_L g186 ( .A1(n_179), .A2(n_157), .B1(n_153), .B2(n_126), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_170), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_182), .B(n_153), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_174), .A2(n_116), .B1(n_146), .B2(n_149), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_164), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_182), .B(n_126), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_170), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_174), .A2(n_124), .B1(n_154), .B2(n_125), .Y(n_194) );
OAI22xp33_ASAP7_75t_L g195 ( .A1(n_175), .A2(n_134), .B1(n_127), .B2(n_144), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g196 ( .A1(n_175), .A2(n_135), .B1(n_137), .B2(n_142), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_170), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_182), .B(n_115), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g199 ( .A1(n_175), .A2(n_138), .B1(n_139), .B2(n_141), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
XOR2xp5_ASAP7_75t_L g201 ( .A(n_161), .B(n_115), .Y(n_201) );
AO22x2_ASAP7_75t_L g202 ( .A1(n_179), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_182), .B(n_119), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_182), .B(n_119), .Y(n_204) );
OAI22xp33_ASAP7_75t_SL g205 ( .A1(n_181), .A2(n_148), .B1(n_158), .B2(n_140), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_161), .A2(n_158), .B1(n_148), .B2(n_133), .Y(n_206) );
BUFx10_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_161), .A2(n_131), .B1(n_130), .B2(n_129), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_161), .A2(n_128), .B1(n_122), .B2(n_121), .Y(n_209) );
INVxp67_ASAP7_75t_L g210 ( .A(n_165), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_166), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_181), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_166), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_164), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_182), .B(n_15), .Y(n_215) );
OAI22xp33_ASAP7_75t_SL g216 ( .A1(n_181), .A2(n_16), .B1(n_17), .B2(n_19), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_166), .A2(n_16), .B1(n_17), .B2(n_19), .Y(n_217) );
OAI22xp33_ASAP7_75t_SL g218 ( .A1(n_181), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
OAI22xp33_ASAP7_75t_L g220 ( .A1(n_176), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_166), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_221) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_179), .B(n_24), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_165), .B(n_25), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_166), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_224) );
OR2x6_ASAP7_75t_L g225 ( .A(n_165), .B(n_26), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g226 ( .A1(n_176), .A2(n_27), .B1(n_28), .B2(n_29), .Y(n_226) );
OAI22xp33_ASAP7_75t_L g227 ( .A1(n_176), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
AND2x2_ASAP7_75t_SL g229 ( .A(n_179), .B(n_164), .Y(n_229) );
OAI22xp33_ASAP7_75t_SL g230 ( .A1(n_178), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_165), .B(n_32), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_229), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_223), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_223), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_231), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_231), .B(n_165), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_210), .B(n_164), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_200), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_229), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_198), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_188), .B(n_164), .Y(n_241) );
XOR2xp5_ASAP7_75t_L g242 ( .A(n_201), .B(n_159), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_200), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_198), .B(n_159), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_219), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_219), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_219), .Y(n_248) );
INVxp67_ASAP7_75t_SL g249 ( .A(n_203), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_192), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_209), .B(n_159), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_192), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_190), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_214), .Y(n_254) );
XOR2xp5_ASAP7_75t_L g255 ( .A(n_201), .B(n_179), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_215), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_215), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_202), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_202), .Y(n_259) );
INVxp33_ASAP7_75t_L g260 ( .A(n_189), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_188), .B(n_179), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_202), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_206), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_203), .Y(n_264) );
XOR2xp5_ASAP7_75t_L g265 ( .A(n_185), .B(n_179), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_183), .Y(n_266) );
XOR2xp5_ASAP7_75t_L g267 ( .A(n_184), .B(n_179), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_191), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_204), .B(n_180), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_204), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_191), .B(n_180), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_222), .Y(n_272) );
NOR2xp67_ASAP7_75t_L g273 ( .A(n_208), .B(n_180), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_202), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_222), .B(n_180), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_183), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_183), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_207), .B(n_178), .Y(n_278) );
NAND2xp33_ASAP7_75t_SL g279 ( .A(n_212), .B(n_178), .Y(n_279) );
INVxp67_ASAP7_75t_SL g280 ( .A(n_194), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_187), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_225), .Y(n_282) );
NAND2x1p5_ASAP7_75t_L g283 ( .A(n_211), .B(n_170), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_225), .Y(n_284) );
NOR2xp33_ASAP7_75t_SL g285 ( .A(n_225), .B(n_173), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_207), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_207), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_187), .Y(n_288) );
AND2x2_ASAP7_75t_SL g289 ( .A(n_213), .B(n_173), .Y(n_289) );
INVxp33_ASAP7_75t_SL g290 ( .A(n_186), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_193), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_225), .Y(n_292) );
INVxp33_ASAP7_75t_L g293 ( .A(n_186), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_193), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_186), .Y(n_295) );
XNOR2x2_ASAP7_75t_L g296 ( .A(n_186), .B(n_173), .Y(n_296) );
XOR2xp5_ASAP7_75t_L g297 ( .A(n_205), .B(n_33), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_238), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_275), .B(n_195), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_255), .B(n_196), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_275), .B(n_199), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_243), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_281), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_236), .B(n_217), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_232), .B(n_221), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_281), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_240), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_236), .B(n_216), .Y(n_309) );
AND2x2_ASAP7_75t_SL g310 ( .A(n_285), .B(n_224), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_243), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_266), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_236), .B(n_218), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_268), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_236), .B(n_220), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_244), .Y(n_316) );
BUFx12f_ASAP7_75t_SL g317 ( .A(n_232), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_266), .B(n_197), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_244), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_246), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_246), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_271), .B(n_226), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_232), .B(n_197), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_271), .B(n_228), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_247), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_232), .B(n_228), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_232), .B(n_35), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_266), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_239), .B(n_170), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_247), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_239), .B(n_170), .Y(n_331) );
AND2x2_ASAP7_75t_SL g332 ( .A(n_258), .B(n_170), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_239), .B(n_35), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_239), .B(n_36), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_266), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_267), .B(n_230), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_266), .B(n_227), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_248), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_248), .Y(n_339) );
INVx4_ASAP7_75t_L g340 ( .A(n_292), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_288), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_239), .B(n_36), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_269), .B(n_37), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_269), .B(n_37), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_278), .Y(n_345) );
AND2x2_ASAP7_75t_SL g346 ( .A(n_258), .B(n_177), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_268), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_276), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_250), .A2(n_162), .B(n_172), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_267), .B(n_38), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_289), .B(n_38), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_249), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_299), .B(n_260), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_351), .B(n_241), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_301), .B(n_272), .Y(n_355) );
BUFx8_ASAP7_75t_SL g356 ( .A(n_327), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_351), .B(n_241), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_348), .B(n_282), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_312), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_312), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_345), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_317), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_328), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_343), .B(n_284), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_341), .Y(n_365) );
NAND2x1_ASAP7_75t_L g366 ( .A(n_312), .B(n_276), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_341), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_301), .B(n_233), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_348), .B(n_277), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_312), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_348), .B(n_345), .Y(n_371) );
BUFx8_ASAP7_75t_L g372 ( .A(n_312), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_328), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_348), .B(n_250), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_345), .B(n_252), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_299), .B(n_280), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_351), .B(n_343), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_340), .B(n_252), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_340), .B(n_264), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_312), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_300), .B(n_292), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_312), .B(n_259), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_341), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_341), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_308), .B(n_265), .Y(n_385) );
BUFx4f_ASAP7_75t_L g386 ( .A(n_312), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_371), .B(n_312), .Y(n_387) );
BUFx4_ASAP7_75t_SL g388 ( .A(n_362), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_372), .Y(n_389) );
BUFx10_ASAP7_75t_L g390 ( .A(n_371), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_365), .B(n_328), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_365), .Y(n_392) );
BUFx2_ASAP7_75t_SL g393 ( .A(n_371), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_372), .Y(n_394) );
INVx3_ASAP7_75t_SL g395 ( .A(n_371), .Y(n_395) );
INVx5_ASAP7_75t_SL g396 ( .A(n_371), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_372), .Y(n_397) );
BUFx2_ASAP7_75t_SL g398 ( .A(n_374), .Y(n_398) );
INVx5_ASAP7_75t_L g399 ( .A(n_356), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_367), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_377), .B(n_351), .Y(n_401) );
INVx6_ASAP7_75t_SL g402 ( .A(n_364), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_367), .Y(n_403) );
OR2x6_ASAP7_75t_L g404 ( .A(n_364), .B(n_259), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_377), .B(n_306), .Y(n_405) );
INVx8_ASAP7_75t_L g406 ( .A(n_356), .Y(n_406) );
INVx5_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
INVx4_ASAP7_75t_L g408 ( .A(n_374), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_372), .Y(n_409) );
BUFx4f_ASAP7_75t_SL g410 ( .A(n_372), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_361), .Y(n_411) );
INVx5_ASAP7_75t_L g412 ( .A(n_374), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_353), .A2(n_336), .B1(n_310), .B2(n_350), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_359), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_383), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_359), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_410), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_388), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_403), .Y(n_419) );
BUFx3_ASAP7_75t_L g420 ( .A(n_389), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_389), .Y(n_421) );
AOI22xp5_ASAP7_75t_SL g422 ( .A1(n_389), .A2(n_290), .B1(n_377), .B2(n_350), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_389), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_402), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_413), .A2(n_353), .B1(n_376), .B2(n_310), .Y(n_425) );
BUFx2_ASAP7_75t_SL g426 ( .A(n_389), .Y(n_426) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_408), .B(n_386), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_410), .Y(n_428) );
BUFx12f_ASAP7_75t_L g429 ( .A(n_399), .Y(n_429) );
BUFx8_ASAP7_75t_L g430 ( .A(n_403), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_413), .A2(n_376), .B1(n_310), .B2(n_357), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_401), .A2(n_310), .B1(n_357), .B2(n_354), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_401), .A2(n_310), .B1(n_357), .B2(n_354), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_398), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_398), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_401), .A2(n_354), .B1(n_336), .B2(n_385), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_398), .A2(n_364), .B1(n_385), .B2(n_361), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_406), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_394), .Y(n_440) );
CKINVDCx11_ASAP7_75t_R g441 ( .A(n_406), .Y(n_441) );
BUFx12f_ASAP7_75t_L g442 ( .A(n_399), .Y(n_442) );
AOI22xp33_ASAP7_75t_SL g443 ( .A1(n_406), .A2(n_385), .B1(n_296), .B2(n_381), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_401), .B(n_355), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_394), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_411), .Y(n_446) );
AOI22xp33_ASAP7_75t_SL g447 ( .A1(n_406), .A2(n_296), .B1(n_381), .B2(n_295), .Y(n_447) );
AOI22xp33_ASAP7_75t_SL g448 ( .A1(n_406), .A2(n_300), .B1(n_340), .B2(n_379), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_405), .A2(n_306), .B1(n_300), .B2(n_293), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_405), .A2(n_306), .B1(n_300), .B2(n_379), .Y(n_450) );
BUFx8_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_406), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_392), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_392), .Y(n_455) );
BUFx2_ASAP7_75t_SL g456 ( .A(n_399), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_405), .A2(n_306), .B1(n_379), .B2(n_289), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_392), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_402), .Y(n_459) );
INVx6_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
BUFx3_ASAP7_75t_L g461 ( .A(n_394), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_416), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_453), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_422), .A2(n_408), .B1(n_412), .B2(n_407), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_422), .A2(n_406), .B1(n_397), .B2(n_394), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_431), .A2(n_402), .B1(n_406), .B2(n_306), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_453), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_431), .A2(n_408), .B1(n_412), .B2(n_407), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_440), .Y(n_469) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_440), .Y(n_470) );
OAI21xp5_ASAP7_75t_SL g471 ( .A1(n_448), .A2(n_242), .B(n_394), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g472 ( .A1(n_438), .A2(n_399), .B1(n_407), .B2(n_412), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_425), .A2(n_443), .B1(n_433), .B2(n_432), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_455), .Y(n_474) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_430), .A2(n_406), .B1(n_397), .B2(n_394), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_428), .B(n_242), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_455), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_443), .A2(n_265), .B(n_255), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_448), .A2(n_408), .B1(n_412), .B2(n_407), .Y(n_479) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_440), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_430), .A2(n_397), .B1(n_409), .B2(n_399), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_425), .A2(n_402), .B1(n_306), .B2(n_408), .Y(n_482) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_430), .A2(n_397), .B1(n_409), .B2(n_399), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_419), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_430), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_430), .Y(n_486) );
OAI21xp5_ASAP7_75t_SL g487 ( .A1(n_447), .A2(n_409), .B(n_397), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_458), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_432), .A2(n_402), .B1(n_306), .B2(n_408), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_458), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_419), .Y(n_491) );
BUFx3_ASAP7_75t_L g492 ( .A(n_428), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_419), .B(n_400), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_433), .A2(n_402), .B1(n_408), .B2(n_412), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_438), .A2(n_407), .B1(n_412), .B2(n_399), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_436), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_451), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_447), .A2(n_297), .B(n_309), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_451), .A2(n_402), .B1(n_412), .B2(n_407), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_436), .Y(n_500) );
BUFx2_ASAP7_75t_SL g501 ( .A(n_417), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_451), .A2(n_407), .B1(n_412), .B2(n_399), .Y(n_502) );
INVx2_ASAP7_75t_SL g503 ( .A(n_451), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_451), .A2(n_407), .B1(n_412), .B2(n_399), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_437), .A2(n_407), .B1(n_412), .B2(n_399), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_437), .A2(n_407), .B1(n_412), .B2(n_399), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_436), .Y(n_507) );
OAI21xp33_ASAP7_75t_L g508 ( .A1(n_420), .A2(n_297), .B(n_309), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_426), .A2(n_397), .B1(n_409), .B2(n_393), .Y(n_509) );
BUFx12f_ASAP7_75t_L g510 ( .A(n_418), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_454), .B(n_400), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_426), .A2(n_409), .B1(n_393), .B2(n_396), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g513 ( .A1(n_420), .A2(n_456), .B1(n_421), .B2(n_423), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_457), .A2(n_409), .B1(n_379), .B2(n_378), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_444), .B(n_400), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_444), .B(n_415), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_462), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_457), .A2(n_379), .B1(n_378), .B2(n_289), .Y(n_518) );
OAI21xp33_ASAP7_75t_L g519 ( .A1(n_420), .A2(n_313), .B(n_167), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_423), .B(n_411), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_420), .A2(n_378), .B1(n_393), .B2(n_404), .Y(n_521) );
OAI21xp5_ASAP7_75t_SL g522 ( .A1(n_421), .A2(n_344), .B(n_343), .Y(n_522) );
BUFx12f_ASAP7_75t_L g523 ( .A(n_441), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_454), .B(n_415), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_460), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_450), .A2(n_378), .B1(n_404), .B2(n_313), .Y(n_526) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_456), .A2(n_396), .B1(n_390), .B2(n_340), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_454), .B(n_415), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_450), .A2(n_364), .B1(n_395), .B2(n_396), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_421), .B(n_387), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_441), .A2(n_378), .B1(n_404), .B2(n_342), .Y(n_531) );
OAI22xp33_ASAP7_75t_L g532 ( .A1(n_417), .A2(n_395), .B1(n_364), .B2(n_340), .Y(n_532) );
OAI21xp5_ASAP7_75t_SL g533 ( .A1(n_421), .A2(n_344), .B(n_343), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_421), .A2(n_396), .B1(n_390), .B2(n_340), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_439), .A2(n_364), .B1(n_395), .B2(n_396), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_449), .A2(n_404), .B1(n_342), .B2(n_327), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_423), .A2(n_396), .B1(n_390), .B2(n_340), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_478), .A2(n_417), .B1(n_429), .B2(n_442), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_471), .A2(n_449), .B1(n_452), .B2(n_439), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_529), .A2(n_429), .B1(n_442), .B2(n_460), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_473), .A2(n_429), .B1(n_442), .B2(n_460), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_465), .A2(n_452), .B1(n_460), .B2(n_435), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_508), .A2(n_460), .B1(n_461), .B2(n_440), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_475), .A2(n_460), .B1(n_434), .B2(n_435), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_485), .A2(n_434), .B1(n_461), .B2(n_427), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_498), .A2(n_461), .B1(n_445), .B2(n_459), .Y(n_546) );
AOI222xp33_ASAP7_75t_L g547 ( .A1(n_523), .A2(n_279), .B1(n_305), .B2(n_344), .C1(n_273), .C2(n_342), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_487), .B(n_167), .C(n_171), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_466), .A2(n_461), .B1(n_445), .B2(n_459), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_463), .B(n_462), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_522), .A2(n_375), .B1(n_364), .B2(n_344), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_468), .A2(n_445), .B1(n_459), .B2(n_424), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_485), .A2(n_445), .B1(n_424), .B2(n_396), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_497), .A2(n_445), .B1(n_424), .B2(n_404), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_497), .A2(n_404), .B1(n_342), .B2(n_327), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_482), .A2(n_404), .B1(n_342), .B2(n_327), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_499), .A2(n_427), .B1(n_395), .B2(n_396), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_505), .A2(n_404), .B1(n_327), .B2(n_342), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_506), .A2(n_404), .B1(n_327), .B2(n_342), .Y(n_559) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_486), .A2(n_427), .B1(n_390), .B2(n_362), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_481), .A2(n_427), .B1(n_395), .B2(n_411), .Y(n_561) );
AOI221xp5_ASAP7_75t_L g562 ( .A1(n_463), .A2(n_251), .B1(n_305), .B2(n_301), .C(n_368), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_489), .A2(n_327), .B1(n_390), .B2(n_262), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_518), .A2(n_390), .B1(n_262), .B2(n_274), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_479), .A2(n_390), .B1(n_274), .B2(n_375), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_484), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_514), .A2(n_375), .B1(n_391), .B2(n_333), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_464), .A2(n_375), .B1(n_391), .B2(n_333), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_515), .B(n_446), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_483), .A2(n_308), .B1(n_391), .B2(n_384), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_535), .A2(n_375), .B1(n_391), .B2(n_333), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_526), .A2(n_391), .B1(n_334), .B2(n_333), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_516), .B(n_446), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_474), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g575 ( .A1(n_533), .A2(n_305), .B1(n_368), .B2(n_283), .C(n_315), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_494), .A2(n_391), .B1(n_334), .B2(n_362), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_486), .A2(n_388), .B1(n_263), .B2(n_391), .Y(n_577) );
AOI22xp5_ASAP7_75t_SL g578 ( .A1(n_486), .A2(n_334), .B1(n_462), .B2(n_384), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_503), .A2(n_383), .B1(n_315), .B2(n_387), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_523), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_495), .A2(n_334), .B1(n_346), .B2(n_332), .Y(n_581) );
OAI21xp5_ASAP7_75t_SL g582 ( .A1(n_503), .A2(n_315), .B(n_283), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_502), .A2(n_352), .B1(n_386), .B2(n_322), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_531), .A2(n_346), .B1(n_332), .B2(n_283), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_536), .A2(n_355), .B1(n_352), .B2(n_337), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_467), .B(n_416), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_472), .A2(n_519), .B1(n_532), .B2(n_530), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_504), .A2(n_337), .B1(n_322), .B2(n_332), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_474), .B(n_416), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_530), .A2(n_346), .B1(n_332), .B2(n_363), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_492), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_527), .A2(n_322), .B1(n_332), .B2(n_346), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_530), .A2(n_346), .B1(n_363), .B2(n_373), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_521), .A2(n_363), .B1(n_373), .B2(n_317), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_501), .A2(n_414), .B1(n_386), .B2(n_416), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_525), .A2(n_373), .B1(n_317), .B2(n_358), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_477), .B(n_414), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_501), .A2(n_373), .B1(n_317), .B2(n_358), .Y(n_598) );
AOI21xp5_ASAP7_75t_SL g599 ( .A1(n_520), .A2(n_374), .B(n_414), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_509), .A2(n_234), .B1(n_235), .B2(n_347), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_477), .B(n_414), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_488), .B(n_414), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_512), .A2(n_513), .B1(n_537), .B2(n_534), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_492), .A2(n_373), .B1(n_358), .B2(n_257), .Y(n_604) );
OAI222xp33_ASAP7_75t_L g605 ( .A1(n_488), .A2(n_490), .B1(n_491), .B2(n_500), .C1(n_507), .C2(n_493), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_490), .B(n_414), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_476), .A2(n_386), .B1(n_347), .B2(n_314), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_493), .A2(n_314), .B1(n_358), .B2(n_270), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_511), .B(n_414), .Y(n_609) );
OA222x2_ASAP7_75t_L g610 ( .A1(n_491), .A2(n_500), .B1(n_507), .B2(n_517), .C1(n_496), .C2(n_484), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_469), .A2(n_386), .B1(n_369), .B2(n_366), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_469), .A2(n_358), .B1(n_256), .B2(n_257), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_517), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_511), .B(n_414), .Y(n_614) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_469), .A2(n_414), .B1(n_359), .B2(n_360), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g616 ( .A1(n_524), .A2(n_171), .B1(n_172), .B2(n_177), .C(n_237), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_469), .A2(n_414), .B1(n_359), .B2(n_360), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_524), .B(n_39), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_528), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_469), .A2(n_369), .B1(n_366), .B2(n_370), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_470), .A2(n_369), .B1(n_380), .B2(n_370), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_470), .A2(n_369), .B1(n_360), .B2(n_359), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_470), .A2(n_167), .B1(n_171), .B2(n_172), .C(n_177), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_528), .A2(n_256), .B1(n_321), .B2(n_311), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_470), .A2(n_382), .B1(n_320), .B2(n_325), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_470), .A2(n_382), .B1(n_320), .B2(n_325), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_496), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_480), .A2(n_320), .B1(n_325), .B2(n_339), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_510), .A2(n_302), .B1(n_311), .B2(n_319), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_480), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_480), .A2(n_320), .B1(n_325), .B2(n_339), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_480), .B(n_162), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_480), .B(n_162), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_510), .A2(n_339), .B1(n_311), .B2(n_316), .Y(n_634) );
OAI221xp5_ASAP7_75t_SL g635 ( .A1(n_471), .A2(n_177), .B1(n_171), .B2(n_172), .C(n_237), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_478), .A2(n_339), .B1(n_330), .B2(n_316), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_463), .Y(n_637) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_485), .A2(n_360), .B1(n_359), .B2(n_328), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_478), .A2(n_303), .B1(n_302), .B2(n_319), .Y(n_639) );
INVx3_ASAP7_75t_L g640 ( .A(n_486), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_471), .A2(n_303), .B1(n_319), .B2(n_321), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_641), .A2(n_167), .B1(n_171), .B2(n_172), .C(n_177), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_574), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_619), .B(n_39), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_574), .B(n_40), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_591), .B(n_177), .C(n_172), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_546), .A2(n_171), .B1(n_162), .B2(n_163), .C(n_169), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_575), .A2(n_162), .B1(n_323), .B2(n_169), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_637), .B(n_40), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_605), .A2(n_162), .B1(n_169), .B2(n_163), .C(n_160), .Y(n_650) );
NAND4xp25_ASAP7_75t_L g651 ( .A(n_547), .B(n_245), .C(n_324), .D(n_349), .Y(n_651) );
OAI21xp33_ASAP7_75t_L g652 ( .A1(n_599), .A2(n_163), .B(n_169), .Y(n_652) );
OAI21xp33_ASAP7_75t_L g653 ( .A1(n_599), .A2(n_163), .B(n_169), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_641), .A2(n_380), .B1(n_370), .B2(n_360), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_597), .B(n_163), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_597), .B(n_163), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_602), .B(n_163), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_637), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_602), .B(n_163), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_539), .A2(n_323), .B1(n_169), .B2(n_163), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_580), .B(n_41), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_550), .B(n_163), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_539), .A2(n_323), .B1(n_169), .B2(n_163), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_603), .A2(n_163), .B1(n_169), .B2(n_168), .C(n_160), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_569), .B(n_41), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_573), .B(n_42), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_550), .B(n_169), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_627), .B(n_43), .Y(n_668) );
OA211x2_ASAP7_75t_L g669 ( .A1(n_540), .A2(n_43), .B(n_318), .C(n_349), .Y(n_669) );
OA21x2_ASAP7_75t_L g670 ( .A1(n_582), .A2(n_380), .B(n_349), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_610), .B(n_169), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_610), .B(n_169), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_613), .B(n_169), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_613), .B(n_160), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_618), .B(n_160), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_566), .B(n_160), .Y(n_676) );
OAI21xp33_ASAP7_75t_L g677 ( .A1(n_587), .A2(n_328), .B(n_318), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_566), .B(n_160), .Y(n_678) );
OAI21xp33_ASAP7_75t_L g679 ( .A1(n_541), .A2(n_335), .B(n_307), .Y(n_679) );
OAI21xp33_ASAP7_75t_SL g680 ( .A1(n_542), .A2(n_261), .B(n_335), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_630), .B(n_160), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_548), .B(n_160), .C(n_168), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_630), .B(n_160), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_609), .B(n_160), .Y(n_684) );
OAI21xp5_ASAP7_75t_SL g685 ( .A1(n_577), .A2(n_261), .B(n_312), .Y(n_685) );
NOR3xp33_ASAP7_75t_L g686 ( .A(n_635), .B(n_326), .C(n_331), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_640), .B(n_160), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_640), .B(n_160), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_578), .B(n_168), .C(n_360), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_560), .B(n_168), .C(n_360), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_551), .A2(n_360), .B1(n_359), .B2(n_335), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_614), .B(n_168), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_608), .B(n_168), .Y(n_693) );
OAI211xp5_ASAP7_75t_SL g694 ( .A1(n_629), .A2(n_253), .B(n_254), .C(n_330), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_601), .B(n_168), .Y(n_695) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_551), .A2(n_335), .B(n_307), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_606), .B(n_168), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_608), .B(n_168), .Y(n_698) );
NOR2xp33_ASAP7_75t_R g699 ( .A(n_580), .B(n_335), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_543), .B(n_168), .C(n_359), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_632), .B(n_168), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_554), .B(n_168), .Y(n_702) );
OAI211xp5_ASAP7_75t_SL g703 ( .A1(n_629), .A2(n_254), .B(n_253), .C(n_330), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_624), .B(n_168), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_624), .B(n_304), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_632), .B(n_45), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_589), .B(n_304), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_586), .B(n_304), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_633), .B(n_47), .Y(n_709) );
OAI21xp5_ASAP7_75t_L g710 ( .A1(n_600), .A2(n_304), .B(n_307), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_570), .A2(n_323), .B1(n_338), .B2(n_321), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_633), .B(n_49), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_538), .A2(n_338), .B1(n_298), .B2(n_302), .C(n_303), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_549), .B(n_307), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_552), .B(n_51), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_585), .B(n_338), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_571), .A2(n_323), .B1(n_316), .B2(n_298), .Y(n_717) );
AOI211xp5_ASAP7_75t_L g718 ( .A1(n_544), .A2(n_331), .B(n_329), .C(n_326), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_585), .B(n_298), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_557), .B(n_52), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_553), .B(n_323), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_595), .B(n_335), .Y(n_722) );
OA211x2_ASAP7_75t_L g723 ( .A1(n_568), .A2(n_54), .B(n_57), .C(n_62), .Y(n_723) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_634), .A2(n_324), .B1(n_326), .B2(n_329), .C(n_331), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_588), .B(n_323), .Y(n_725) );
OAI21xp5_ASAP7_75t_SL g726 ( .A1(n_561), .A2(n_331), .B(n_329), .Y(n_726) );
OAI21xp5_ASAP7_75t_SL g727 ( .A1(n_592), .A2(n_329), .B(n_324), .Y(n_727) );
OAI221xp5_ASAP7_75t_L g728 ( .A1(n_636), .A2(n_324), .B1(n_326), .B2(n_277), .C(n_287), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_588), .B(n_579), .Y(n_729) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_607), .A2(n_294), .B1(n_291), .B2(n_288), .C(n_287), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g731 ( .A1(n_592), .A2(n_286), .B(n_294), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_545), .B(n_63), .Y(n_732) );
AOI211xp5_ASAP7_75t_L g733 ( .A1(n_583), .A2(n_286), .B(n_291), .C(n_66), .Y(n_733) );
OAI21xp5_ASAP7_75t_SL g734 ( .A1(n_638), .A2(n_64), .B(n_65), .Y(n_734) );
NOR3xp33_ASAP7_75t_L g735 ( .A(n_623), .B(n_67), .C(n_69), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_615), .B(n_71), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_565), .B(n_73), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_617), .B(n_74), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_556), .B(n_75), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_562), .B(n_113), .C(n_78), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_621), .B(n_76), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_567), .B(n_576), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_639), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_743) );
OAI21xp33_ASAP7_75t_L g744 ( .A1(n_555), .A2(n_82), .B(n_83), .Y(n_744) );
AND2x2_ASAP7_75t_SL g745 ( .A(n_581), .B(n_84), .Y(n_745) );
NAND4xp25_ASAP7_75t_L g746 ( .A(n_604), .B(n_86), .C(n_87), .D(n_89), .Y(n_746) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_620), .B(n_112), .C(n_93), .Y(n_747) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_611), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g749 ( .A(n_699), .Y(n_749) );
AOI211xp5_ASAP7_75t_L g750 ( .A1(n_671), .A2(n_616), .B(n_622), .C(n_598), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_643), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_748), .B(n_559), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_644), .B(n_594), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_643), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_658), .B(n_558), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_655), .B(n_593), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_655), .B(n_563), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_658), .B(n_572), .Y(n_758) );
OR2x2_ASAP7_75t_L g759 ( .A(n_656), .B(n_631), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_665), .B(n_612), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_666), .B(n_596), .Y(n_761) );
CKINVDCx6p67_ASAP7_75t_R g762 ( .A(n_745), .Y(n_762) );
NOR3xp33_ASAP7_75t_SL g763 ( .A(n_685), .B(n_584), .C(n_590), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_656), .B(n_564), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_657), .B(n_628), .Y(n_765) );
AND2x4_ASAP7_75t_L g766 ( .A(n_671), .B(n_625), .Y(n_766) );
INVx3_ASAP7_75t_L g767 ( .A(n_672), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_659), .B(n_626), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_659), .B(n_92), .Y(n_769) );
NAND4xp75_ASAP7_75t_L g770 ( .A(n_672), .B(n_94), .C(n_96), .D(n_98), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_662), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_662), .Y(n_772) );
NAND3xp33_ASAP7_75t_L g773 ( .A(n_664), .B(n_101), .C(n_103), .Y(n_773) );
OAI211xp5_ASAP7_75t_L g774 ( .A1(n_680), .A2(n_111), .B(n_105), .C(n_107), .Y(n_774) );
OR2x6_ASAP7_75t_L g775 ( .A(n_722), .B(n_104), .Y(n_775) );
OAI22xp5_ASAP7_75t_SL g776 ( .A1(n_745), .A2(n_108), .B1(n_109), .B2(n_110), .Y(n_776) );
OR2x2_ASAP7_75t_L g777 ( .A(n_667), .B(n_729), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_667), .B(n_676), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_673), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_668), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_674), .B(n_676), .Y(n_781) );
XNOR2xp5_ASAP7_75t_L g782 ( .A(n_718), .B(n_651), .Y(n_782) );
OR2x2_ASAP7_75t_L g783 ( .A(n_678), .B(n_707), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_674), .B(n_678), .Y(n_784) );
NOR3xp33_ASAP7_75t_L g785 ( .A(n_661), .B(n_690), .C(n_746), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_681), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_681), .B(n_683), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_670), .B(n_683), .Y(n_788) );
NOR3xp33_ASAP7_75t_SL g789 ( .A(n_734), .B(n_703), .C(n_694), .Y(n_789) );
NAND3xp33_ASAP7_75t_L g790 ( .A(n_650), .B(n_700), .C(n_733), .Y(n_790) );
NAND4xp75_ASAP7_75t_L g791 ( .A(n_669), .B(n_723), .C(n_731), .D(n_722), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_645), .Y(n_792) );
NOR2xp33_ASAP7_75t_SL g793 ( .A(n_689), .B(n_652), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_708), .B(n_725), .Y(n_794) );
AOI221x1_ASAP7_75t_SL g795 ( .A1(n_742), .A2(n_649), .B1(n_696), .B2(n_679), .C(n_677), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_670), .B(n_684), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_670), .B(n_684), .Y(n_797) );
INVx1_ASAP7_75t_SL g798 ( .A(n_699), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_695), .B(n_697), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_692), .B(n_697), .Y(n_800) );
AOI211xp5_ASAP7_75t_L g801 ( .A1(n_726), .A2(n_727), .B(n_653), .C(n_744), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_669), .A2(n_663), .B1(n_660), .B2(n_692), .Y(n_802) );
NAND4xp75_ASAP7_75t_L g803 ( .A(n_720), .B(n_715), .C(n_732), .D(n_736), .Y(n_803) );
AO21x2_ASAP7_75t_L g804 ( .A1(n_687), .A2(n_688), .B(n_720), .Y(n_804) );
NAND4xp75_ASAP7_75t_L g805 ( .A(n_715), .B(n_736), .C(n_738), .D(n_721), .Y(n_805) );
NOR3xp33_ASAP7_75t_L g806 ( .A(n_740), .B(n_642), .C(n_682), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_702), .B(n_675), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_717), .A2(n_728), .B1(n_711), .B2(n_739), .Y(n_808) );
OAI211xp5_ASAP7_75t_SL g809 ( .A1(n_648), .A2(n_698), .B(n_693), .C(n_647), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_695), .B(n_701), .Y(n_810) );
OR2x2_ASAP7_75t_L g811 ( .A(n_705), .B(n_714), .Y(n_811) );
NOR3xp33_ASAP7_75t_L g812 ( .A(n_646), .B(n_747), .C(n_713), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_716), .B(n_719), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_706), .B(n_709), .Y(n_814) );
OAI211xp5_ASAP7_75t_SL g815 ( .A1(n_704), .A2(n_737), .B(n_724), .C(n_743), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_706), .B(n_712), .Y(n_816) );
AOI221xp5_ASAP7_75t_L g817 ( .A1(n_691), .A2(n_654), .B1(n_739), .B2(n_710), .C(n_686), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_709), .B(n_712), .Y(n_818) );
AOI22xp33_ASAP7_75t_SL g819 ( .A1(n_738), .A2(n_741), .B1(n_735), .B2(n_730), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_671), .B(n_672), .C(n_664), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_748), .B(n_619), .Y(n_821) );
NAND4xp75_ASAP7_75t_L g822 ( .A(n_671), .B(n_672), .C(n_745), .D(n_669), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_643), .Y(n_823) );
NOR2x1_ASAP7_75t_L g824 ( .A(n_671), .B(n_485), .Y(n_824) );
NAND4xp25_ASAP7_75t_L g825 ( .A(n_671), .B(n_672), .C(n_664), .D(n_669), .Y(n_825) );
OAI21xp5_ASAP7_75t_L g826 ( .A1(n_685), .A2(n_745), .B(n_680), .Y(n_826) );
NOR3xp33_ASAP7_75t_L g827 ( .A(n_664), .B(n_661), .C(n_671), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_644), .B(n_591), .Y(n_828) );
XOR2x2_ASAP7_75t_L g829 ( .A(n_805), .B(n_782), .Y(n_829) );
INVx2_ASAP7_75t_SL g830 ( .A(n_824), .Y(n_830) );
NOR2xp33_ASAP7_75t_R g831 ( .A(n_762), .B(n_749), .Y(n_831) );
XOR2x2_ASAP7_75t_L g832 ( .A(n_803), .B(n_822), .Y(n_832) );
OR2x2_ASAP7_75t_L g833 ( .A(n_821), .B(n_777), .Y(n_833) );
BUFx2_ASAP7_75t_L g834 ( .A(n_749), .Y(n_834) );
NAND4xp75_ASAP7_75t_L g835 ( .A(n_826), .B(n_763), .C(n_752), .D(n_789), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_751), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_788), .B(n_796), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_754), .Y(n_838) );
NAND4xp75_ASAP7_75t_L g839 ( .A(n_763), .B(n_752), .C(n_789), .D(n_797), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_788), .B(n_796), .Y(n_840) );
XOR2x2_ASAP7_75t_L g841 ( .A(n_776), .B(n_785), .Y(n_841) );
XOR2xp5_ASAP7_75t_L g842 ( .A(n_794), .B(n_783), .Y(n_842) );
NOR4xp25_ASAP7_75t_L g843 ( .A(n_780), .B(n_792), .C(n_820), .D(n_825), .Y(n_843) );
NOR3xp33_ASAP7_75t_L g844 ( .A(n_774), .B(n_790), .C(n_791), .Y(n_844) );
NAND4xp75_ASAP7_75t_L g845 ( .A(n_797), .B(n_817), .C(n_753), .D(n_761), .Y(n_845) );
XNOR2xp5_ASAP7_75t_L g846 ( .A(n_795), .B(n_810), .Y(n_846) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_823), .Y(n_847) );
NAND4xp75_ASAP7_75t_L g848 ( .A(n_753), .B(n_761), .C(n_828), .D(n_760), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_762), .A2(n_767), .B1(n_827), .B2(n_813), .Y(n_849) );
OR2x2_ASAP7_75t_L g850 ( .A(n_772), .B(n_771), .Y(n_850) );
BUFx6f_ASAP7_75t_L g851 ( .A(n_775), .Y(n_851) );
NAND3xp33_ASAP7_75t_L g852 ( .A(n_801), .B(n_767), .C(n_828), .Y(n_852) );
NAND4xp75_ASAP7_75t_L g853 ( .A(n_760), .B(n_802), .C(n_807), .D(n_813), .Y(n_853) );
INVx1_ASAP7_75t_SL g854 ( .A(n_798), .Y(n_854) );
NAND4xp75_ASAP7_75t_L g855 ( .A(n_807), .B(n_768), .C(n_769), .D(n_756), .Y(n_855) );
AND4x1_ASAP7_75t_L g856 ( .A(n_793), .B(n_750), .C(n_812), .D(n_808), .Y(n_856) );
NAND4xp75_ASAP7_75t_L g857 ( .A(n_768), .B(n_755), .C(n_814), .D(n_765), .Y(n_857) );
NAND4xp75_ASAP7_75t_L g858 ( .A(n_814), .B(n_779), .C(n_758), .D(n_818), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_804), .B(n_816), .Y(n_859) );
NOR2xp33_ASAP7_75t_SL g860 ( .A(n_770), .B(n_775), .Y(n_860) );
NAND3xp33_ASAP7_75t_L g861 ( .A(n_806), .B(n_819), .C(n_766), .Y(n_861) );
XOR2xp5_ASAP7_75t_L g862 ( .A(n_799), .B(n_759), .Y(n_862) );
XOR2x2_ASAP7_75t_L g863 ( .A(n_808), .B(n_800), .Y(n_863) );
INVx3_ASAP7_75t_L g864 ( .A(n_775), .Y(n_864) );
NAND4xp75_ASAP7_75t_L g865 ( .A(n_757), .B(n_764), .C(n_778), .D(n_787), .Y(n_865) );
XOR2x2_ASAP7_75t_L g866 ( .A(n_766), .B(n_764), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_835), .A2(n_815), .B1(n_786), .B2(n_809), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_847), .Y(n_868) );
XOR2x2_ASAP7_75t_L g869 ( .A(n_829), .B(n_811), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_847), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_837), .B(n_840), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_856), .B(n_784), .Y(n_872) );
XOR2x2_ASAP7_75t_L g873 ( .A(n_829), .B(n_781), .Y(n_873) );
BUFx3_ASAP7_75t_L g874 ( .A(n_834), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_836), .Y(n_875) );
INVxp67_ASAP7_75t_SL g876 ( .A(n_864), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_838), .Y(n_877) );
INVx3_ASAP7_75t_L g878 ( .A(n_851), .Y(n_878) );
CKINVDCx16_ASAP7_75t_R g879 ( .A(n_831), .Y(n_879) );
INVxp67_ASAP7_75t_L g880 ( .A(n_853), .Y(n_880) );
INVx1_ASAP7_75t_SL g881 ( .A(n_854), .Y(n_881) );
INVxp67_ASAP7_75t_L g882 ( .A(n_848), .Y(n_882) );
XNOR2x1_ASAP7_75t_L g883 ( .A(n_841), .B(n_773), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_844), .A2(n_861), .B1(n_841), .B2(n_832), .Y(n_884) );
INVx1_ASAP7_75t_SL g885 ( .A(n_831), .Y(n_885) );
XNOR2x2_ASAP7_75t_L g886 ( .A(n_845), .B(n_839), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_850), .Y(n_887) );
AO22x2_ASAP7_75t_L g888 ( .A1(n_852), .A2(n_857), .B1(n_830), .B2(n_858), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_850), .Y(n_889) );
XOR2xp5_ASAP7_75t_L g890 ( .A(n_879), .B(n_832), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_887), .Y(n_891) );
AO22x2_ASAP7_75t_L g892 ( .A1(n_883), .A2(n_864), .B1(n_865), .B2(n_830), .Y(n_892) );
OAI22x1_ASAP7_75t_L g893 ( .A1(n_885), .A2(n_846), .B1(n_849), .B2(n_864), .Y(n_893) );
AOI22x1_ASAP7_75t_L g894 ( .A1(n_888), .A2(n_851), .B1(n_843), .B2(n_837), .Y(n_894) );
AO22x2_ASAP7_75t_L g895 ( .A1(n_883), .A2(n_855), .B1(n_862), .B2(n_842), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_875), .Y(n_896) );
INVxp33_ASAP7_75t_SL g897 ( .A(n_867), .Y(n_897) );
BUFx3_ASAP7_75t_L g898 ( .A(n_874), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_877), .Y(n_899) );
INVx3_ASAP7_75t_L g900 ( .A(n_878), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_874), .Y(n_901) );
OA22x2_ASAP7_75t_L g902 ( .A1(n_880), .A2(n_882), .B1(n_876), .B2(n_881), .Y(n_902) );
INVxp67_ASAP7_75t_L g903 ( .A(n_886), .Y(n_903) );
AOI22x1_ASAP7_75t_SL g904 ( .A1(n_886), .A2(n_863), .B1(n_866), .B2(n_860), .Y(n_904) );
OA22x2_ASAP7_75t_L g905 ( .A1(n_878), .A2(n_859), .B1(n_863), .B2(n_866), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_901), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_898), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_898), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_896), .Y(n_909) );
NOR2xp33_ASAP7_75t_R g910 ( .A(n_903), .B(n_884), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_899), .Y(n_911) );
OAI322xp33_ASAP7_75t_L g912 ( .A1(n_905), .A2(n_872), .A3(n_868), .B1(n_870), .B2(n_878), .C1(n_833), .C2(n_889), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_891), .Y(n_913) );
INVxp67_ASAP7_75t_L g914 ( .A(n_902), .Y(n_914) );
OA22x2_ASAP7_75t_L g915 ( .A1(n_914), .A2(n_890), .B1(n_893), .B2(n_904), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_907), .Y(n_916) );
OA22x2_ASAP7_75t_SL g917 ( .A1(n_908), .A2(n_895), .B1(n_890), .B2(n_892), .Y(n_917) );
INVx2_ASAP7_75t_SL g918 ( .A(n_906), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_914), .A2(n_895), .B1(n_905), .B2(n_892), .Y(n_919) );
O2A1O1Ixp33_ASAP7_75t_SL g920 ( .A1(n_919), .A2(n_897), .B(n_910), .C(n_895), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_915), .A2(n_897), .B1(n_893), .B2(n_902), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_917), .A2(n_892), .B1(n_894), .B2(n_888), .Y(n_922) );
AOI221xp5_ASAP7_75t_SL g923 ( .A1(n_922), .A2(n_912), .B1(n_917), .B2(n_916), .C(n_909), .Y(n_923) );
NOR4xp25_ASAP7_75t_L g924 ( .A(n_920), .B(n_918), .C(n_911), .D(n_913), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_921), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_925), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_925), .Y(n_927) );
NAND3xp33_ASAP7_75t_L g928 ( .A(n_926), .B(n_923), .C(n_924), .Y(n_928) );
NOR2x1_ASAP7_75t_L g929 ( .A(n_926), .B(n_927), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_929), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_928), .Y(n_931) );
AO22x2_ASAP7_75t_L g932 ( .A1(n_931), .A2(n_891), .B1(n_869), .B2(n_900), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_932), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_933), .A2(n_930), .B1(n_869), .B2(n_873), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_934), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_935), .A2(n_888), .B1(n_900), .B2(n_868), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_936), .Y(n_937) );
AOI221xp5_ASAP7_75t_L g938 ( .A1(n_937), .A2(n_888), .B1(n_900), .B2(n_870), .C(n_873), .Y(n_938) );
AOI211xp5_ASAP7_75t_L g939 ( .A1(n_938), .A2(n_871), .B(n_833), .C(n_889), .Y(n_939) );
endmodule