module fake_netlist_6_3475_n_170 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_170);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;

output n_170;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_21;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_39;
wire n_73;
wire n_148;
wire n_138;
wire n_22;
wire n_161;
wire n_68;
wire n_166;
wire n_28;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_24;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_23;
wire n_142;
wire n_20;
wire n_143;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVxp33_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_19),
.B(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_25),
.B(n_2),
.Y(n_46)
);

AO21x2_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_2),
.B(n_3),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_26),
.B(n_3),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_4),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_34),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_4),
.Y(n_56)
);

NOR2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_5),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_22),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR3xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_51),
.C(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2x1_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_11),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_8),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_62),
.Y(n_71)
);

OAI22x1_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_57),
.B1(n_53),
.B2(n_66),
.Y(n_72)
);

OAI21x1_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_48),
.B(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_49),
.B(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

OAI21x1_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_37),
.B(n_39),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_47),
.B1(n_36),
.B2(n_41),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_41),
.B1(n_39),
.B2(n_42),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_54),
.B(n_67),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_42),
.B(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_59),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

AOI221x1_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_50),
.B1(n_47),
.B2(n_10),
.C(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_47),
.Y(n_87)
);

OAI31xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_64),
.A3(n_70),
.B(n_77),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_69),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_64),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_64),
.B(n_77),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_76),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_76),
.B(n_82),
.Y(n_94)
);

AOI21x1_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_73),
.B(n_79),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_72),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_72),
.B(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_79),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_79),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_87),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_88),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_94),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_103),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_103),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

OAI21x1_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_91),
.B(n_95),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_85),
.C(n_92),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_92),
.B(n_85),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_92),
.B(n_104),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_102),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_105),
.B(n_104),
.C(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_101),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_105),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_105),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_107),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_108),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_131),
.B(n_118),
.Y(n_142)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_127),
.A3(n_126),
.B1(n_121),
.B2(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_127),
.B1(n_113),
.B2(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_114),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_140),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_118),
.B(n_120),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_142),
.B1(n_148),
.B2(n_143),
.C(n_139),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_118),
.B(n_123),
.Y(n_151)
);

AOI32xp33_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_129),
.A3(n_134),
.B1(n_137),
.B2(n_130),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_134),
.B1(n_113),
.B2(n_123),
.Y(n_153)
);

OAI321xp33_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_141),
.A3(n_128),
.B1(n_113),
.B2(n_135),
.C(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_152),
.Y(n_161)
);

AO22x2_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_141),
.B1(n_117),
.B2(n_123),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_122),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_161),
.A3(n_163),
.B1(n_159),
.B2(n_162),
.C1(n_158),
.C2(n_117),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_122),
.B1(n_117),
.B2(n_92),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_165),
.Y(n_168)
);

OAI21x1_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_122),
.B(n_92),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_122),
.B1(n_168),
.B2(n_164),
.Y(n_170)
);


endmodule