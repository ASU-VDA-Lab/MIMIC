module real_aes_15822_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_1404;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1544;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g1069 ( .A1(n_0), .A2(n_3), .B1(n_863), .B2(n_1070), .Y(n_1069) );
AOI22xp33_ASAP7_75t_SL g1108 ( .A1(n_0), .A2(n_239), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_1), .A2(n_220), .B1(n_1429), .B2(n_1431), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g1452 ( .A1(n_1), .A2(n_187), .B1(n_1453), .B2(n_1454), .Y(n_1452) );
INVx1_ASAP7_75t_L g438 ( .A(n_2), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_3), .A2(n_241), .B1(n_829), .B2(n_1109), .Y(n_1113) );
XNOR2xp5_ASAP7_75t_L g757 ( .A(n_4), .B(n_758), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_5), .A2(n_260), .B1(n_1110), .B2(n_1126), .Y(n_1125) );
INVxp33_ASAP7_75t_SL g1155 ( .A(n_5), .Y(n_1155) );
INVx1_ASAP7_75t_L g1514 ( .A(n_6), .Y(n_1514) );
OAI211xp5_ASAP7_75t_L g880 ( .A1(n_7), .A2(n_568), .B(n_623), .C(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g892 ( .A(n_7), .Y(n_892) );
AOI22xp5_ASAP7_75t_SL g1204 ( .A1(n_8), .A2(n_257), .B1(n_1184), .B2(n_1191), .Y(n_1204) );
INVx1_ASAP7_75t_L g294 ( .A(n_9), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_9), .B(n_304), .Y(n_458) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_9), .B(n_227), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1446 ( .A(n_9), .B(n_397), .Y(n_1446) );
INVx1_ASAP7_75t_L g1086 ( .A(n_10), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_10), .A2(n_25), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
INVx1_ASAP7_75t_L g897 ( .A(n_11), .Y(n_897) );
INVx1_ASAP7_75t_L g840 ( .A(n_12), .Y(n_840) );
OAI211xp5_ASAP7_75t_L g926 ( .A1(n_13), .A2(n_642), .B(n_927), .C(n_929), .Y(n_926) );
INVx1_ASAP7_75t_L g937 ( .A(n_13), .Y(n_937) );
INVx1_ASAP7_75t_L g1092 ( .A(n_14), .Y(n_1092) );
INVx2_ASAP7_75t_L g1179 ( .A(n_15), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_15), .B(n_1180), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_15), .B(n_100), .Y(n_1187) );
INVx1_ASAP7_75t_L g1421 ( .A(n_16), .Y(n_1421) );
OAI221xp5_ASAP7_75t_L g1462 ( .A1(n_16), .A2(n_159), .B1(n_1463), .B2(n_1467), .C(n_1472), .Y(n_1462) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_17), .A2(n_124), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
OAI22xp33_ASAP7_75t_L g1012 ( .A1(n_17), .A2(n_124), .B1(n_296), .B2(n_1013), .Y(n_1012) );
AOI22xp5_ASAP7_75t_SL g1214 ( .A1(n_18), .A2(n_132), .B1(n_1184), .B2(n_1191), .Y(n_1214) );
INVx1_ASAP7_75t_L g945 ( .A(n_19), .Y(n_945) );
OAI22xp33_ASAP7_75t_L g682 ( .A1(n_20), .A2(n_160), .B1(n_406), .B2(n_683), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g685 ( .A1(n_20), .A2(n_270), .B1(n_316), .B2(n_639), .Y(n_685) );
AOI22xp5_ASAP7_75t_SL g1224 ( .A1(n_21), .A2(n_252), .B1(n_1181), .B2(n_1186), .Y(n_1224) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_22), .Y(n_659) );
XNOR2x2_ASAP7_75t_SL g922 ( .A(n_23), .B(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g1522 ( .A(n_24), .Y(n_1522) );
INVx1_ASAP7_75t_L g1089 ( .A(n_25), .Y(n_1089) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_26), .A2(n_209), .B1(n_400), .B2(n_633), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_26), .A2(n_96), .B1(n_316), .B2(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g931 ( .A(n_27), .Y(n_931) );
OAI211xp5_ASAP7_75t_L g935 ( .A1(n_27), .A2(n_750), .B(n_904), .C(n_936), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_28), .A2(n_106), .B1(n_890), .B2(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1163 ( .A(n_28), .Y(n_1163) );
INVx1_ASAP7_75t_L g1521 ( .A(n_29), .Y(n_1521) );
INVx1_ASAP7_75t_L g422 ( .A(n_30), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g1175 ( .A1(n_31), .A2(n_179), .B1(n_1176), .B2(n_1181), .Y(n_1175) );
INVx1_ASAP7_75t_L g709 ( .A(n_32), .Y(n_709) );
INVx1_ASAP7_75t_L g777 ( .A(n_33), .Y(n_777) );
INVx1_ASAP7_75t_L g1093 ( .A(n_34), .Y(n_1093) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_35), .Y(n_665) );
INVx1_ASAP7_75t_L g978 ( .A(n_36), .Y(n_978) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_37), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g879 ( .A1(n_38), .A2(n_120), .B1(n_683), .B2(n_850), .Y(n_879) );
OAI22xp33_ASAP7_75t_L g893 ( .A1(n_38), .A2(n_49), .B1(n_358), .B2(n_639), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_39), .A2(n_97), .B1(n_1184), .B2(n_1201), .Y(n_1268) );
OAI22xp33_ASAP7_75t_L g805 ( .A1(n_40), .A2(n_163), .B1(n_406), .B2(n_633), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_40), .A2(n_114), .B1(n_316), .B2(n_354), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_41), .A2(n_278), .B1(n_316), .B2(n_355), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_41), .A2(n_43), .B1(n_683), .B2(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g765 ( .A(n_42), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_43), .A2(n_181), .B1(n_358), .B2(n_639), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g1183 ( .A1(n_44), .A2(n_180), .B1(n_1184), .B2(n_1186), .Y(n_1183) );
AOI22xp5_ASAP7_75t_L g1192 ( .A1(n_45), .A2(n_88), .B1(n_1176), .B2(n_1184), .Y(n_1192) );
INVx1_ASAP7_75t_L g802 ( .A(n_46), .Y(n_802) );
OAI211xp5_ASAP7_75t_L g808 ( .A1(n_46), .A2(n_642), .B(n_809), .C(n_810), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_47), .A2(n_131), .B1(n_314), .B2(n_323), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_47), .A2(n_131), .B1(n_296), .B2(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g320 ( .A(n_48), .Y(n_320) );
INVx1_ASAP7_75t_L g336 ( .A(n_48), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g884 ( .A1(n_49), .A2(n_213), .B1(n_633), .B2(n_885), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_50), .A2(n_75), .B1(n_863), .B2(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1107 ( .A(n_50), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_51), .A2(n_273), .B1(n_1176), .B2(n_1181), .Y(n_1194) );
INVx1_ASAP7_75t_L g782 ( .A(n_52), .Y(n_782) );
INVx1_ASAP7_75t_L g740 ( .A(n_53), .Y(n_740) );
OAI22xp33_ASAP7_75t_L g753 ( .A1(n_53), .A2(n_162), .B1(n_406), .B2(n_633), .Y(n_753) );
OAI211xp5_ASAP7_75t_L g622 ( .A1(n_54), .A2(n_477), .B(n_623), .C(n_626), .Y(n_622) );
INVx1_ASAP7_75t_L g646 ( .A(n_54), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_55), .A2(n_208), .B1(n_510), .B2(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_55), .A2(n_214), .B1(n_546), .B2(n_550), .Y(n_553) );
INVx1_ASAP7_75t_L g287 ( .A(n_56), .Y(n_287) );
INVx2_ASAP7_75t_L g322 ( .A(n_57), .Y(n_322) );
OAI22xp33_ASAP7_75t_L g1143 ( .A1(n_58), .A2(n_225), .B1(n_394), .B2(n_1020), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1151 ( .A1(n_58), .A2(n_225), .B1(n_1009), .B2(n_1152), .Y(n_1151) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_59), .A2(n_244), .B1(n_735), .B2(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_59), .A2(n_183), .B1(n_865), .B2(n_867), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g1225 ( .A1(n_60), .A2(n_71), .B1(n_1176), .B2(n_1184), .Y(n_1225) );
INVx1_ASAP7_75t_L g839 ( .A(n_61), .Y(n_839) );
INVx1_ASAP7_75t_L g883 ( .A(n_62), .Y(n_883) );
INVx1_ASAP7_75t_L g705 ( .A(n_63), .Y(n_705) );
INVx1_ASAP7_75t_L g837 ( .A(n_64), .Y(n_837) );
INVx1_ASAP7_75t_L g952 ( .A(n_65), .Y(n_952) );
OAI22xp33_ASAP7_75t_L g1054 ( .A1(n_66), .A2(n_266), .B1(n_355), .B2(n_358), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_66), .A2(n_266), .B1(n_683), .B2(n_850), .Y(n_1060) );
OAI22xp33_ASAP7_75t_SL g1048 ( .A1(n_67), .A2(n_277), .B1(n_316), .B2(n_639), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g1056 ( .A1(n_67), .A2(n_277), .B1(n_633), .B2(n_885), .Y(n_1056) );
OAI222xp33_ASAP7_75t_L g498 ( .A1(n_68), .A2(n_104), .B1(n_237), .B2(n_499), .C1(n_501), .C2(n_502), .Y(n_498) );
OAI222xp33_ASAP7_75t_L g565 ( .A1(n_68), .A2(n_104), .B1(n_237), .B2(n_388), .C1(n_566), .C2(n_568), .Y(n_565) );
INVx1_ASAP7_75t_L g900 ( .A(n_69), .Y(n_900) );
INVx1_ASAP7_75t_L g1132 ( .A(n_70), .Y(n_1132) );
INVx1_ASAP7_75t_L g1082 ( .A(n_72), .Y(n_1082) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_73), .A2(n_96), .B1(n_395), .B2(n_406), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g647 ( .A1(n_73), .A2(n_209), .B1(n_355), .B2(n_358), .Y(n_647) );
OAI211xp5_ASAP7_75t_L g1003 ( .A1(n_74), .A2(n_338), .B(n_1004), .C(n_1005), .Y(n_1003) );
INVx1_ASAP7_75t_L g1018 ( .A(n_74), .Y(n_1018) );
INVxp67_ASAP7_75t_SL g1112 ( .A(n_75), .Y(n_1112) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_76), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_77), .A2(n_279), .B1(n_519), .B2(n_522), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_77), .A2(n_129), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_78), .A2(n_129), .B1(n_530), .B2(n_531), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_78), .A2(n_279), .B1(n_546), .B2(n_550), .Y(n_545) );
INVx1_ASAP7_75t_L g1517 ( .A(n_79), .Y(n_1517) );
AOI221xp5_ASAP7_75t_L g823 ( .A1(n_80), .A2(n_276), .B1(n_531), .B2(n_824), .C(n_825), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_80), .A2(n_127), .B1(n_556), .B2(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g1031 ( .A(n_81), .Y(n_1031) );
INVx1_ASAP7_75t_L g1141 ( .A(n_82), .Y(n_1141) );
INVx1_ASAP7_75t_L g988 ( .A(n_83), .Y(n_988) );
INVx1_ASAP7_75t_L g1028 ( .A(n_84), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g1190 ( .A1(n_85), .A2(n_192), .B1(n_1181), .B2(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1087 ( .A(n_86), .Y(n_1087) );
INVx1_ASAP7_75t_L g710 ( .A(n_87), .Y(n_710) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_89), .Y(n_801) );
INVx1_ASAP7_75t_L g576 ( .A(n_90), .Y(n_576) );
INVx1_ASAP7_75t_L g975 ( .A(n_91), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g1500 ( .A1(n_92), .A2(n_228), .B1(n_562), .B2(n_1501), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g1504 ( .A1(n_92), .A2(n_228), .B1(n_1505), .B2(n_1506), .Y(n_1504) );
INVx1_ASAP7_75t_L g430 ( .A(n_93), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_94), .A2(n_117), .B1(n_1110), .B2(n_1136), .Y(n_1427) );
AOI221xp5_ASAP7_75t_L g1448 ( .A1(n_94), .A2(n_248), .B1(n_1449), .B2(n_1450), .C(n_1451), .Y(n_1448) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_95), .Y(n_289) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_95), .B(n_287), .Y(n_1177) );
INVx1_ASAP7_75t_L g951 ( .A(n_98), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g1199 ( .A1(n_99), .A2(n_158), .B1(n_1176), .B2(n_1181), .Y(n_1199) );
INVx1_ASAP7_75t_L g1180 ( .A(n_100), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_100), .B(n_1179), .Y(n_1185) );
AOI22xp5_ASAP7_75t_L g1205 ( .A1(n_101), .A2(n_190), .B1(n_1176), .B2(n_1181), .Y(n_1205) );
XOR2x2_ASAP7_75t_L g1390 ( .A(n_101), .B(n_1391), .Y(n_1390) );
AOI22xp5_ASAP7_75t_L g1487 ( .A1(n_101), .A2(n_1488), .B1(n_1537), .B2(n_1539), .Y(n_1487) );
INVx1_ASAP7_75t_L g776 ( .A(n_102), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_103), .A2(n_1490), .B1(n_1491), .B2(n_1492), .Y(n_1489) );
CKINVDCx5p33_ASAP7_75t_R g1490 ( .A(n_103), .Y(n_1490) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_105), .Y(n_661) );
INVx1_ASAP7_75t_L g1156 ( .A(n_106), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_107), .A2(n_229), .B1(n_495), .B2(n_496), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_107), .A2(n_229), .B1(n_562), .B2(n_563), .Y(n_561) );
INVx2_ASAP7_75t_L g365 ( .A(n_108), .Y(n_365) );
INVx1_ASAP7_75t_L g446 ( .A(n_108), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_108), .B(n_322), .Y(n_1397) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_109), .Y(n_584) );
INVx1_ASAP7_75t_L g903 ( .A(n_110), .Y(n_903) );
INVx1_ASAP7_75t_L g947 ( .A(n_111), .Y(n_947) );
XOR2xp5_ASAP7_75t_L g969 ( .A(n_112), .B(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g1037 ( .A(n_113), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_114), .A2(n_121), .B1(n_562), .B2(n_804), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g1403 ( .A1(n_115), .A2(n_142), .B1(n_1404), .B2(n_1408), .Y(n_1403) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_116), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_117), .A2(n_261), .B1(n_1454), .B2(n_1478), .Y(n_1477) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_118), .A2(n_187), .B1(n_531), .B2(n_1429), .Y(n_1428) );
AOI21xp33_ASAP7_75t_L g1474 ( .A1(n_118), .A2(n_1450), .B(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g490 ( .A(n_119), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g887 ( .A1(n_120), .A2(n_213), .B1(n_316), .B2(n_355), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_121), .A2(n_163), .B1(n_323), .B2(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g452 ( .A(n_122), .Y(n_452) );
INVx1_ASAP7_75t_L g907 ( .A(n_123), .Y(n_907) );
INVx1_ASAP7_75t_L g713 ( .A(n_125), .Y(n_713) );
INVx1_ASAP7_75t_L g985 ( .A(n_126), .Y(n_985) );
AOI221xp5_ASAP7_75t_L g826 ( .A1(n_127), .A2(n_222), .B1(n_531), .B2(n_824), .C(n_827), .Y(n_826) );
OAI22xp33_ASAP7_75t_L g932 ( .A1(n_128), .A2(n_235), .B1(n_316), .B2(n_933), .Y(n_932) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_128), .A2(n_235), .B1(n_406), .B2(n_633), .Y(n_940) );
INVx1_ASAP7_75t_L g1035 ( .A(n_130), .Y(n_1035) );
XOR2xp5_ASAP7_75t_L g486 ( .A(n_133), .B(n_487), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_134), .Y(n_678) );
INVx1_ASAP7_75t_L g1123 ( .A(n_135), .Y(n_1123) );
INVx1_ASAP7_75t_L g1267 ( .A(n_136), .Y(n_1267) );
CKINVDCx5p33_ASAP7_75t_R g1402 ( .A(n_137), .Y(n_1402) );
INVx1_ASAP7_75t_L g958 ( .A(n_138), .Y(n_958) );
INVx1_ASAP7_75t_L g905 ( .A(n_139), .Y(n_905) );
AOI31xp33_ASAP7_75t_L g818 ( .A1(n_140), .A2(n_819), .A3(n_833), .B(n_843), .Y(n_818) );
NAND2xp33_ASAP7_75t_SL g860 ( .A(n_140), .B(n_861), .Y(n_860) );
INVxp67_ASAP7_75t_SL g874 ( .A(n_140), .Y(n_874) );
INVx1_ASAP7_75t_L g1053 ( .A(n_141), .Y(n_1053) );
OAI211xp5_ASAP7_75t_L g1057 ( .A1(n_141), .A2(n_623), .B(n_662), .C(n_1058), .Y(n_1057) );
OAI211xp5_ASAP7_75t_L g1443 ( .A1(n_142), .A2(n_1444), .B(n_1447), .C(n_1456), .Y(n_1443) );
INVx1_ASAP7_75t_L g738 ( .A(n_143), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_143), .A2(n_258), .B1(n_562), .B2(n_747), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g1200 ( .A1(n_144), .A2(n_185), .B1(n_1184), .B2(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g733 ( .A(n_145), .Y(n_733) );
OA211x2_ASAP7_75t_L g749 ( .A1(n_145), .A2(n_568), .B(n_750), .C(n_751), .Y(n_749) );
BUFx3_ASAP7_75t_L g318 ( .A(n_146), .Y(n_318) );
INVx1_ASAP7_75t_L g1029 ( .A(n_147), .Y(n_1029) );
INVx1_ASAP7_75t_L g1032 ( .A(n_148), .Y(n_1032) );
INVx1_ASAP7_75t_L g898 ( .A(n_149), .Y(n_898) );
INVx1_ASAP7_75t_L g420 ( .A(n_150), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_151), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_152), .Y(n_666) );
INVx1_ASAP7_75t_L g1068 ( .A(n_153), .Y(n_1068) );
OAI22xp5_ASAP7_75t_SL g693 ( .A1(n_154), .A2(n_694), .B1(n_744), .B2(n_755), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_154), .B(n_695), .C(n_715), .D(n_727), .Y(n_694) );
INVx1_ASAP7_75t_L g1007 ( .A(n_155), .Y(n_1007) );
OAI211xp5_ASAP7_75t_L g1014 ( .A1(n_155), .A2(n_378), .B(n_1015), .C(n_1017), .Y(n_1014) );
CKINVDCx5p33_ASAP7_75t_R g1052 ( .A(n_156), .Y(n_1052) );
OAI22xp33_ASAP7_75t_L g1138 ( .A1(n_157), .A2(n_253), .B1(n_296), .B2(n_406), .Y(n_1138) );
OAI22xp33_ASAP7_75t_L g1145 ( .A1(n_157), .A2(n_253), .B1(n_323), .B2(n_1146), .Y(n_1145) );
XNOR2x1_ASAP7_75t_L g1023 ( .A(n_158), .B(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1416 ( .A(n_159), .Y(n_1416) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_160), .A2(n_275), .B1(n_355), .B2(n_358), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g663 ( .A(n_161), .Y(n_663) );
INVx1_ASAP7_75t_L g737 ( .A(n_162), .Y(n_737) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_164), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_165), .A2(n_214), .B1(n_510), .B2(n_516), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_165), .A2(n_208), .B1(n_538), .B2(n_542), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_166), .Y(n_654) );
INVx1_ASAP7_75t_L g1133 ( .A(n_167), .Y(n_1133) );
INVx1_ASAP7_75t_L g780 ( .A(n_168), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g1195 ( .A1(n_169), .A2(n_218), .B1(n_1184), .B2(n_1191), .Y(n_1195) );
XOR2x2_ASAP7_75t_L g876 ( .A(n_170), .B(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g426 ( .A(n_171), .Y(n_426) );
INVx1_ASAP7_75t_L g1142 ( .A(n_172), .Y(n_1142) );
OAI211xp5_ASAP7_75t_L g1147 ( .A1(n_172), .A2(n_338), .B(n_789), .C(n_1148), .Y(n_1147) );
OAI211xp5_ASAP7_75t_L g798 ( .A1(n_173), .A2(n_750), .B(n_799), .C(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g811 ( .A(n_173), .Y(n_811) );
OAI22xp33_ASAP7_75t_L g1502 ( .A1(n_174), .A2(n_207), .B1(n_296), .B2(n_406), .Y(n_1502) );
OAI22xp33_ASAP7_75t_L g1510 ( .A1(n_174), .A2(n_207), .B1(n_314), .B2(n_323), .Y(n_1510) );
INVx1_ASAP7_75t_L g348 ( .A(n_175), .Y(n_348) );
INVx1_ASAP7_75t_L g831 ( .A(n_176), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_176), .A2(n_244), .B1(n_543), .B2(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g955 ( .A(n_177), .Y(n_955) );
INVx1_ASAP7_75t_L g959 ( .A(n_178), .Y(n_959) );
INVxp67_ASAP7_75t_SL g847 ( .A(n_181), .Y(n_847) );
INVx1_ASAP7_75t_L g1083 ( .A(n_182), .Y(n_1083) );
INVx1_ASAP7_75t_L g830 ( .A(n_183), .Y(n_830) );
INVx1_ASAP7_75t_L g767 ( .A(n_184), .Y(n_767) );
OAI211xp5_ASAP7_75t_L g1049 ( .A1(n_186), .A2(n_642), .B(n_1050), .C(n_1051), .Y(n_1049) );
INVx1_ASAP7_75t_L g1059 ( .A(n_186), .Y(n_1059) );
OAI22xp33_ASAP7_75t_L g1434 ( .A1(n_188), .A2(n_249), .B1(n_1435), .B2(n_1438), .Y(n_1434) );
INVx1_ASAP7_75t_L g1457 ( .A(n_188), .Y(n_1457) );
INVx1_ASAP7_75t_L g700 ( .A(n_189), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g925 ( .A1(n_191), .A2(n_204), .B1(n_355), .B2(n_356), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_191), .A2(n_204), .B1(n_395), .B2(n_804), .Y(n_939) );
CKINVDCx20_ASAP7_75t_R g1527 ( .A(n_193), .Y(n_1527) );
INVx1_ASAP7_75t_L g908 ( .A(n_194), .Y(n_908) );
OAI211xp5_ASAP7_75t_SL g1495 ( .A1(n_195), .A2(n_750), .B(n_1015), .C(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1509 ( .A(n_195), .Y(n_1509) );
INVx1_ASAP7_75t_L g1515 ( .A(n_196), .Y(n_1515) );
OAI211xp5_ASAP7_75t_SL g330 ( .A1(n_197), .A2(n_331), .B(n_338), .C(n_342), .Y(n_330) );
INVx1_ASAP7_75t_L g392 ( .A(n_197), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_198), .Y(n_658) );
INVx1_ASAP7_75t_L g702 ( .A(n_199), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_200), .Y(n_587) );
INVx1_ASAP7_75t_L g983 ( .A(n_201), .Y(n_983) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_202), .A2(n_264), .B1(n_354), .B2(n_356), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_202), .A2(n_264), .B1(n_394), .B2(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g699 ( .A(n_203), .Y(n_699) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_205), .Y(n_300) );
INVx1_ASAP7_75t_L g987 ( .A(n_206), .Y(n_987) );
INVx1_ASAP7_75t_L g680 ( .A(n_210), .Y(n_680) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_210), .A2(n_449), .B(n_642), .C(n_687), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_211), .Y(n_582) );
INVx1_ASAP7_75t_L g882 ( .A(n_212), .Y(n_882) );
INVx1_ASAP7_75t_L g956 ( .A(n_215), .Y(n_956) );
OAI211xp5_ASAP7_75t_L g1139 ( .A1(n_216), .A2(n_373), .B(n_378), .C(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g1150 ( .A(n_216), .Y(n_1150) );
INVx1_ASAP7_75t_L g1034 ( .A(n_217), .Y(n_1034) );
INVx1_ASAP7_75t_L g901 ( .A(n_219), .Y(n_901) );
INVx1_ASAP7_75t_L g1473 ( .A(n_220), .Y(n_1473) );
INVx1_ASAP7_75t_L g1498 ( .A(n_221), .Y(n_1498) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_222), .A2(n_276), .B1(n_865), .B2(n_867), .Y(n_864) );
INVx1_ASAP7_75t_L g979 ( .A(n_223), .Y(n_979) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_224), .Y(n_628) );
INVx1_ASAP7_75t_L g1519 ( .A(n_226), .Y(n_1519) );
BUFx3_ASAP7_75t_L g304 ( .A(n_227), .Y(n_304) );
INVx1_ASAP7_75t_L g397 ( .A(n_227), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_230), .A2(n_259), .B1(n_354), .B2(n_1009), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_230), .A2(n_259), .B1(n_562), .B2(n_1020), .Y(n_1019) );
XOR2x2_ASAP7_75t_L g310 ( .A(n_231), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g732 ( .A(n_232), .Y(n_732) );
INVx1_ASAP7_75t_L g714 ( .A(n_233), .Y(n_714) );
OAI211xp5_ASAP7_75t_L g676 ( .A1(n_234), .A2(n_477), .B(n_623), .C(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g688 ( .A(n_234), .Y(n_688) );
INVx1_ASAP7_75t_L g440 ( .A(n_236), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_238), .Y(n_595) );
INVxp67_ASAP7_75t_SL g1072 ( .A(n_239), .Y(n_1072) );
INVx1_ASAP7_75t_L g1038 ( .A(n_240), .Y(n_1038) );
INVxp67_ASAP7_75t_SL g1073 ( .A(n_241), .Y(n_1073) );
INVx1_ASAP7_75t_L g370 ( .A(n_242), .Y(n_370) );
INVx1_ASAP7_75t_L g445 ( .A(n_242), .Y(n_445) );
INVx2_ASAP7_75t_L g457 ( .A(n_242), .Y(n_457) );
INVx1_ASAP7_75t_L g762 ( .A(n_243), .Y(n_762) );
INVx1_ASAP7_75t_L g930 ( .A(n_245), .Y(n_930) );
INVx1_ASAP7_75t_L g1006 ( .A(n_246), .Y(n_1006) );
INVx1_ASAP7_75t_L g1067 ( .A(n_247), .Y(n_1067) );
AOI22xp33_ASAP7_75t_SL g1433 ( .A1(n_248), .A2(n_261), .B1(n_1110), .B2(n_1136), .Y(n_1433) );
INVx1_ASAP7_75t_L g1460 ( .A(n_249), .Y(n_1460) );
XNOR2x1_ASAP7_75t_L g1118 ( .A(n_250), .B(n_1119), .Y(n_1118) );
AOI22xp5_ASAP7_75t_L g1213 ( .A1(n_251), .A2(n_268), .B1(n_1176), .B2(n_1181), .Y(n_1213) );
XNOR2xp5_ASAP7_75t_L g1063 ( .A(n_254), .B(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1265 ( .A(n_254), .Y(n_1265) );
INVx1_ASAP7_75t_L g1499 ( .A(n_255), .Y(n_1499) );
OAI211xp5_ASAP7_75t_L g1507 ( .A1(n_255), .A2(n_331), .B(n_338), .C(n_1508), .Y(n_1507) );
INVx1_ASAP7_75t_L g771 ( .A(n_256), .Y(n_771) );
INVx1_ASAP7_75t_L g742 ( .A(n_258), .Y(n_742) );
INVxp67_ASAP7_75t_SL g1161 ( .A(n_260), .Y(n_1161) );
INVx1_ASAP7_75t_L g974 ( .A(n_262), .Y(n_974) );
INVx1_ASAP7_75t_L g1124 ( .A(n_263), .Y(n_1124) );
INVx1_ASAP7_75t_L g448 ( .A(n_265), .Y(n_448) );
INVx1_ASAP7_75t_L g734 ( .A(n_267), .Y(n_734) );
XNOR2xp5_ASAP7_75t_L g649 ( .A(n_268), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g352 ( .A(n_269), .Y(n_352) );
OAI211xp5_ASAP7_75t_L g372 ( .A1(n_269), .A2(n_373), .B(n_378), .C(n_383), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_270), .A2(n_275), .B1(n_400), .B2(n_633), .Y(n_681) );
INVx1_ASAP7_75t_L g492 ( .A(n_271), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_272), .Y(n_603) );
INVx1_ASAP7_75t_L g1525 ( .A(n_274), .Y(n_1525) );
INVx1_ASAP7_75t_L g845 ( .A(n_278), .Y(n_845) );
INVx1_ASAP7_75t_L g631 ( .A(n_280), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g641 ( .A1(n_280), .A2(n_449), .B(n_642), .C(n_643), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_305), .B(n_1167), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_290), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g1486 ( .A(n_284), .B(n_293), .Y(n_1486) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g1538 ( .A(n_286), .B(n_289), .Y(n_1538) );
INVx1_ASAP7_75t_L g1543 ( .A(n_286), .Y(n_1543) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g1545 ( .A(n_289), .B(n_1543), .Y(n_1545) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g411 ( .A(n_293), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g480 ( .A(n_294), .B(n_304), .Y(n_480) );
AND2x4_ASAP7_75t_L g1476 ( .A(n_294), .B(n_303), .Y(n_1476) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_295), .A2(n_407), .B1(n_490), .B2(n_492), .Y(n_559) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_295), .A2(n_407), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
AND2x4_ASAP7_75t_SL g1485 ( .A(n_295), .B(n_1486), .Y(n_1485) );
INVx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_302), .Y(n_296) );
OR2x6_ASAP7_75t_L g395 ( .A(n_297), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g683 ( .A(n_297), .B(n_396), .Y(n_683) );
BUFx4f_ASAP7_75t_L g721 ( .A(n_297), .Y(n_721) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx4f_ASAP7_75t_L g463 ( .A(n_298), .Y(n_463) );
INVx3_ASAP7_75t_L g634 ( .A(n_298), .Y(n_634) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2x1_ASAP7_75t_L g377 ( .A(n_300), .B(n_301), .Y(n_377) );
AND2x2_ASAP7_75t_L g382 ( .A(n_300), .B(n_301), .Y(n_382) );
INVx1_ASAP7_75t_L g391 ( .A(n_300), .Y(n_391) );
INVx2_ASAP7_75t_L g404 ( .A(n_300), .Y(n_404) );
AND2x2_ASAP7_75t_L g408 ( .A(n_300), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g472 ( .A(n_300), .Y(n_472) );
BUFx2_ASAP7_75t_L g386 ( .A(n_301), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_301), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g409 ( .A(n_301), .Y(n_409) );
OR2x2_ASAP7_75t_L g471 ( .A(n_301), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g541 ( .A(n_301), .Y(n_541) );
AND2x2_ASAP7_75t_L g544 ( .A(n_301), .B(n_404), .Y(n_544) );
OR2x6_ASAP7_75t_L g633 ( .A(n_302), .B(n_634), .Y(n_633) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g380 ( .A(n_303), .Y(n_380) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g385 ( .A(n_304), .Y(n_385) );
AND2x4_ASAP7_75t_L g389 ( .A(n_304), .B(n_390), .Y(n_389) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B1(n_917), .B2(n_918), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
XNOR2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_571), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_310), .B1(n_484), .B2(n_485), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND3xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_371), .C(n_414), .Y(n_311) );
OAI31xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_330), .A3(n_353), .B(n_361), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_315), .A2(n_324), .B1(n_1092), .B2(n_1093), .Y(n_1100) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_SL g491 ( .A(n_316), .Y(n_491) );
INVx1_ASAP7_75t_L g741 ( .A(n_316), .Y(n_741) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_316), .Y(n_1001) );
OR2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_321), .Y(n_316) );
OR2x4_ASAP7_75t_L g355 ( .A(n_317), .B(n_325), .Y(n_355) );
BUFx3_ASAP7_75t_L g421 ( .A(n_317), .Y(n_421) );
BUFx4f_ASAP7_75t_L g583 ( .A(n_317), .Y(n_583) );
INVx2_ASAP7_75t_L g600 ( .A(n_317), .Y(n_600) );
BUFx3_ASAP7_75t_L g788 ( .A(n_317), .Y(n_788) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g329 ( .A(n_318), .Y(n_329) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_318), .Y(n_337) );
AND2x4_ASAP7_75t_L g340 ( .A(n_318), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_318), .B(n_336), .Y(n_360) );
INVx1_ASAP7_75t_L g515 ( .A(n_319), .Y(n_515) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVxp67_ASAP7_75t_L g328 ( .A(n_320), .Y(n_328) );
INVx1_ASAP7_75t_L g325 ( .A(n_321), .Y(n_325) );
AND2x4_ASAP7_75t_L g339 ( .A(n_321), .B(n_340), .Y(n_339) );
OR2x6_ASAP7_75t_L g358 ( .A(n_321), .B(n_359), .Y(n_358) );
NAND3x1_ASAP7_75t_L g443 ( .A(n_321), .B(n_444), .C(n_446), .Y(n_443) );
NAND2x1p5_ASAP7_75t_L g605 ( .A(n_321), .B(n_446), .Y(n_605) );
AND2x4_ASAP7_75t_L g1410 ( .A(n_321), .B(n_1411), .Y(n_1410) );
INVx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g346 ( .A(n_322), .Y(n_346) );
NAND2xp33_ASAP7_75t_SL g418 ( .A(n_322), .B(n_365), .Y(n_418) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_324), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_489) );
INVx2_ASAP7_75t_L g933 ( .A(n_324), .Y(n_933) );
INVx1_ASAP7_75t_L g1002 ( .A(n_324), .Y(n_1002) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g640 ( .A(n_325), .B(n_326), .Y(n_640) );
INVx2_ASAP7_75t_L g588 ( .A(n_326), .Y(n_588) );
INVx2_ASAP7_75t_L g793 ( .A(n_326), .Y(n_793) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_326), .Y(n_824) );
INVx1_ASAP7_75t_L g984 ( .A(n_326), .Y(n_984) );
INVx2_ASAP7_75t_L g1106 ( .A(n_326), .Y(n_1106) );
BUFx6f_ASAP7_75t_L g1131 ( .A(n_326), .Y(n_1131) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_327), .Y(n_429) );
INVx2_ASAP7_75t_L g521 ( .A(n_327), .Y(n_521) );
BUFx8_ASAP7_75t_L g708 ( .A(n_327), .Y(n_708) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x4_ASAP7_75t_L g514 ( .A(n_329), .B(n_515), .Y(n_514) );
OAI22xp33_ASAP7_75t_L g1534 ( .A1(n_331), .A2(n_1515), .B1(n_1522), .B2(n_1535), .Y(n_1534) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g501 ( .A(n_332), .Y(n_501) );
INVx1_ASAP7_75t_L g789 ( .A(n_332), .Y(n_789) );
INVx1_ASAP7_75t_L g809 ( .A(n_332), .Y(n_809) );
INVx1_ASAP7_75t_L g915 ( .A(n_332), .Y(n_915) );
INVx4_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx3_ASAP7_75t_L g424 ( .A(n_333), .Y(n_424) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_333), .Y(n_669) );
OR2x2_ASAP7_75t_L g1405 ( .A(n_333), .B(n_1396), .Y(n_1405) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx2_ASAP7_75t_L g451 ( .A(n_334), .Y(n_451) );
BUFx3_ASAP7_75t_L g602 ( .A(n_334), .Y(n_602) );
NAND2x1p5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
BUFx2_ASAP7_75t_L g351 ( .A(n_335), .Y(n_351) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g341 ( .A(n_336), .Y(n_341) );
BUFx2_ASAP7_75t_L g347 ( .A(n_337), .Y(n_347) );
AND2x4_ASAP7_75t_L g524 ( .A(n_337), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g1419 ( .A(n_337), .Y(n_1419) );
CKINVDCx8_ASAP7_75t_R g338 ( .A(n_339), .Y(n_338) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_339), .B(n_494), .C(n_498), .Y(n_493) );
CKINVDCx8_ASAP7_75t_R g642 ( .A(n_339), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_339), .B(n_730), .Y(n_729) );
AOI211xp5_ASAP7_75t_L g1095 ( .A1(n_339), .A2(n_1087), .B(n_1096), .C(n_1097), .Y(n_1095) );
INVx2_ASAP7_75t_L g517 ( .A(n_340), .Y(n_517) );
BUFx2_ASAP7_75t_L g528 ( .A(n_340), .Y(n_528) );
BUFx2_ASAP7_75t_L g735 ( .A(n_340), .Y(n_735) );
BUFx3_ASAP7_75t_L g829 ( .A(n_340), .Y(n_829) );
BUFx2_ASAP7_75t_L g890 ( .A(n_340), .Y(n_890) );
BUFx2_ASAP7_75t_L g1110 ( .A(n_340), .Y(n_1110) );
INVx1_ASAP7_75t_L g525 ( .A(n_341), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_348), .B1(n_349), .B2(n_352), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_343), .A2(n_349), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
BUFx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g1149 ( .A(n_344), .Y(n_1149) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
AND2x4_ASAP7_75t_L g350 ( .A(n_345), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g500 ( .A(n_345), .B(n_347), .Y(n_500) );
AND2x4_ASAP7_75t_L g644 ( .A(n_345), .B(n_347), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_345), .B(n_351), .Y(n_645) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND3x4_ASAP7_75t_L g507 ( .A(n_346), .B(n_365), .C(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_348), .A2(n_384), .B1(n_387), .B2(n_392), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_349), .A2(n_1141), .B1(n_1149), .B2(n_1150), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1508 ( .A1(n_349), .A2(n_1149), .B1(n_1498), .B2(n_1509), .Y(n_1508) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g502 ( .A(n_350), .Y(n_502) );
AOI222xp33_ASAP7_75t_L g731 ( .A1(n_350), .A2(n_644), .B1(n_732), .B2(n_733), .C1(n_734), .C2(n_735), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_350), .A2(n_500), .B1(n_801), .B2(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_350), .A2(n_500), .B1(n_930), .B2(n_931), .Y(n_929) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g495 ( .A(n_355), .Y(n_495) );
INVx2_ASAP7_75t_SL g743 ( .A(n_355), .Y(n_743) );
BUFx2_ASAP7_75t_L g1505 ( .A(n_355), .Y(n_1505) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_357), .A2(n_640), .B1(n_737), .B2(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g497 ( .A(n_358), .Y(n_497) );
BUFx3_ASAP7_75t_L g813 ( .A(n_358), .Y(n_813) );
INVx1_ASAP7_75t_L g1010 ( .A(n_358), .Y(n_1010) );
BUFx3_ASAP7_75t_L g439 ( .A(n_359), .Y(n_439) );
INVx1_ASAP7_75t_L g597 ( .A(n_359), .Y(n_597) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g433 ( .A(n_360), .Y(n_433) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI31xp33_ASAP7_75t_L g1144 ( .A1(n_362), .A2(n_1145), .A3(n_1147), .B(n_1151), .Y(n_1144) );
OAI31xp33_ASAP7_75t_L g1503 ( .A1(n_362), .A2(n_1504), .A3(n_1507), .B(n_1510), .Y(n_1503) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_363), .B(n_366), .Y(n_362) );
AND2x4_ASAP7_75t_L g504 ( .A(n_363), .B(n_366), .Y(n_504) );
AND2x2_ASAP7_75t_L g648 ( .A(n_363), .B(n_366), .Y(n_648) );
AND2x2_ASAP7_75t_L g814 ( .A(n_363), .B(n_366), .Y(n_814) );
AND2x2_ASAP7_75t_L g842 ( .A(n_363), .B(n_366), .Y(n_842) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g1411 ( .A(n_365), .Y(n_1411) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g417 ( .A(n_368), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g482 ( .A(n_368), .Y(n_482) );
AND2x2_ASAP7_75t_SL g620 ( .A(n_368), .B(n_480), .Y(n_620) );
OR2x2_ASAP7_75t_L g1396 ( .A(n_368), .B(n_1397), .Y(n_1396) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g413 ( .A(n_369), .Y(n_413) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI31xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_393), .A3(n_405), .B(n_410), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_375), .A2(n_616), .B1(n_951), .B2(n_955), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_375), .A2(n_616), .B1(n_947), .B2(n_959), .Y(n_965) );
BUFx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_SL g569 ( .A(n_376), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_376), .A2(n_584), .B1(n_603), .B2(n_616), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_376), .A2(n_613), .B1(n_658), .B2(n_659), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_376), .A2(n_975), .B1(n_988), .B2(n_996), .Y(n_995) );
BUFx2_ASAP7_75t_SL g1159 ( .A(n_376), .Y(n_1159) );
OAI22xp5_ASAP7_75t_L g1520 ( .A1(n_376), .A2(n_996), .B1(n_1521), .B2(n_1522), .Y(n_1520) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_377), .Y(n_475) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_379), .B(n_561), .C(n_565), .Y(n_560) );
INVx3_ASAP7_75t_L g750 ( .A(n_379), .Y(n_750) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AND2x2_ASAP7_75t_L g624 ( .A(n_380), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g627 ( .A(n_380), .B(n_386), .Y(n_627) );
OR2x2_ASAP7_75t_L g850 ( .A(n_380), .B(n_402), .Y(n_850) );
BUFx3_ASAP7_75t_L g867 ( .A(n_381), .Y(n_867) );
BUFx6f_ASAP7_75t_L g1090 ( .A(n_381), .Y(n_1090) );
BUFx3_ASAP7_75t_L g1449 ( .A(n_381), .Y(n_1449) );
AND2x6_ASAP7_75t_L g1455 ( .A(n_381), .B(n_1401), .Y(n_1455) );
AND2x4_ASAP7_75t_SL g1466 ( .A(n_381), .B(n_1446), .Y(n_1466) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g552 ( .A(n_382), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g936 ( .A1(n_384), .A2(n_930), .B1(n_937), .B2(n_938), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_384), .A2(n_629), .B1(n_1052), .B2(n_1059), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_384), .A2(n_389), .B1(n_1141), .B2(n_1142), .Y(n_1140) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
OR2x2_ASAP7_75t_L g401 ( .A(n_385), .B(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g567 ( .A(n_385), .B(n_386), .Y(n_567) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_385), .B(n_872), .Y(n_1081) );
INVx1_ASAP7_75t_L g1470 ( .A(n_386), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_387), .A2(n_567), .B1(n_732), .B2(n_734), .Y(n_751) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g938 ( .A(n_388), .Y(n_938) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g630 ( .A(n_389), .Y(n_630) );
BUFx3_ASAP7_75t_L g679 ( .A(n_389), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_389), .A2(n_627), .B1(n_837), .B2(n_839), .Y(n_852) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_389), .A2(n_567), .B1(n_1006), .B2(n_1018), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1407 ( .A(n_390), .B(n_1401), .Y(n_1407) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_395), .Y(n_562) );
AND2x4_ASAP7_75t_L g407 ( .A(n_396), .B(n_408), .Y(n_407) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g1080 ( .A1(n_399), .A2(n_1081), .B1(n_1082), .B2(n_1083), .C(n_1084), .Y(n_1080) );
INVx2_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
HB1xp67_ASAP7_75t_L g1501 ( .A(n_400), .Y(n_1501) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g564 ( .A(n_401), .Y(n_564) );
INVx2_ASAP7_75t_L g748 ( .A(n_401), .Y(n_748) );
INVx8_ASAP7_75t_L g466 ( .A(n_402), .Y(n_466) );
BUFx2_ASAP7_75t_L g722 ( .A(n_402), .Y(n_722) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_407), .A2(n_845), .B1(n_846), .B2(n_847), .Y(n_844) );
INVx4_ASAP7_75t_L g885 ( .A(n_407), .Y(n_885) );
INVx3_ASAP7_75t_SL g1013 ( .A(n_407), .Y(n_1013) );
INVx2_ASAP7_75t_L g549 ( .A(n_408), .Y(n_549) );
BUFx6f_ASAP7_75t_L g866 ( .A(n_408), .Y(n_866) );
BUFx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g570 ( .A(n_411), .Y(n_570) );
BUFx2_ASAP7_75t_L g636 ( .A(n_411), .Y(n_636) );
OAI31xp33_ASAP7_75t_L g878 ( .A1(n_411), .A2(n_879), .A3(n_880), .B(n_884), .Y(n_878) );
BUFx2_ASAP7_75t_SL g941 ( .A(n_411), .Y(n_941) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g1406 ( .A(n_413), .B(n_1407), .Y(n_1406) );
INVxp67_ASAP7_75t_L g1412 ( .A(n_413), .Y(n_1412) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_453), .Y(n_414) );
OAI33xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_419), .A3(n_425), .B1(n_434), .B2(n_441), .B3(n_447), .Y(n_415) );
OAI33xp33_ASAP7_75t_L g696 ( .A1(n_416), .A2(n_697), .A3(n_701), .B1(n_706), .B2(n_711), .B3(n_712), .Y(n_696) );
OAI33xp33_ASAP7_75t_L g943 ( .A1(n_416), .A2(n_711), .A3(n_944), .B1(n_950), .B2(n_953), .B3(n_957), .Y(n_943) );
OAI22xp33_ASAP7_75t_L g1104 ( .A1(n_416), .A2(n_1105), .B1(n_1111), .B2(n_1114), .Y(n_1104) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx4f_ASAP7_75t_L g580 ( .A(n_417), .Y(n_580) );
BUFx8_ASAP7_75t_L g784 ( .A(n_417), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_420), .A2(n_448), .B1(n_460), .B2(n_464), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g447 ( .A1(n_421), .A2(n_448), .B1(n_449), .B2(n_452), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g712 ( .A1(n_421), .A2(n_669), .B1(n_713), .B2(n_714), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g973 ( .A1(n_421), .A2(n_974), .B1(n_975), .B2(n_976), .Y(n_973) );
OAI22xp33_ASAP7_75t_L g986 ( .A1(n_421), .A2(n_915), .B1(n_987), .B2(n_988), .Y(n_986) );
OAI22xp33_ASAP7_75t_L g1529 ( .A1(n_421), .A2(n_1514), .B1(n_1521), .B2(n_1530), .Y(n_1529) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_422), .A2(n_452), .B1(n_468), .B2(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx3_ASAP7_75t_L g585 ( .A(n_424), .Y(n_585) );
INVx2_ASAP7_75t_L g796 ( .A(n_424), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_430), .B2(n_431), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_426), .A2(n_438), .B1(n_468), .B2(n_473), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_427), .A2(n_978), .B1(n_979), .B2(n_980), .Y(n_977) );
BUFx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx8_ASAP7_75t_L g1429 ( .A(n_428), .Y(n_1429) );
INVx5_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g437 ( .A(n_429), .Y(n_437) );
INVx2_ASAP7_75t_SL g672 ( .A(n_429), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_430), .A2(n_440), .B1(n_460), .B2(n_464), .Y(n_483) );
OAI22xp33_ASAP7_75t_SL g792 ( .A1(n_431), .A2(n_771), .B1(n_782), .B2(n_793), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_431), .A2(n_983), .B1(n_984), .B2(n_985), .Y(n_982) );
CKINVDCx8_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g590 ( .A(n_432), .Y(n_590) );
INVx3_ASAP7_75t_L g673 ( .A(n_432), .Y(n_673) );
INVx3_ASAP7_75t_L g913 ( .A(n_432), .Y(n_913) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g704 ( .A(n_433), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_438), .B1(n_439), .B2(n_440), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_437), .A2(n_590), .B1(n_900), .B2(n_907), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_437), .A2(n_913), .B1(n_1028), .B2(n_1029), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_439), .A2(n_767), .B1(n_780), .B2(n_791), .Y(n_790) );
OAI221xp5_ASAP7_75t_L g1105 ( .A1(n_439), .A2(n_1067), .B1(n_1106), .B2(n_1107), .C(n_1108), .Y(n_1105) );
OAI221xp5_ASAP7_75t_L g1122 ( .A1(n_439), .A2(n_791), .B1(n_1123), .B2(n_1124), .C(n_1125), .Y(n_1122) );
OAI221xp5_ASAP7_75t_L g1129 ( .A1(n_439), .A2(n_1130), .B1(n_1132), .B2(n_1133), .C(n_1134), .Y(n_1129) );
OAI22xp5_ASAP7_75t_L g1531 ( .A1(n_439), .A2(n_1517), .B1(n_1525), .B2(n_1532), .Y(n_1531) );
OAI22xp5_ASAP7_75t_L g1533 ( .A1(n_439), .A2(n_588), .B1(n_1519), .B2(n_1527), .Y(n_1533) );
INVx1_ASAP7_75t_L g532 ( .A(n_441), .Y(n_532) );
OAI33xp33_ASAP7_75t_L g972 ( .A1(n_441), .A2(n_784), .A3(n_973), .B1(n_977), .B2(n_982), .B3(n_986), .Y(n_972) );
OAI33xp33_ASAP7_75t_L g1528 ( .A1(n_441), .A2(n_784), .A3(n_1529), .B1(n_1531), .B2(n_1533), .B3(n_1534), .Y(n_1528) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g794 ( .A(n_442), .Y(n_794) );
INVx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx3_ASAP7_75t_L g1116 ( .A(n_443), .Y(n_1116) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g1399 ( .A(n_445), .Y(n_1399) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g949 ( .A(n_451), .Y(n_949) );
OAI33xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_459), .A3(n_467), .B1(n_476), .B2(n_478), .B3(n_483), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g536 ( .A(n_455), .Y(n_536) );
INVx2_ASAP7_75t_L g607 ( .A(n_455), .Y(n_607) );
INVx4_ASAP7_75t_L g719 ( .A(n_455), .Y(n_719) );
AND2x4_ASAP7_75t_L g455 ( .A(n_456), .B(n_458), .Y(n_455) );
OR2x2_ASAP7_75t_L g604 ( .A(n_456), .B(n_605), .Y(n_604) );
OR2x6_ASAP7_75t_L g711 ( .A(n_456), .B(n_605), .Y(n_711) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g508 ( .A(n_457), .Y(n_508) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx4_ASAP7_75t_L g609 ( .A(n_463), .Y(n_609) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_463), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g998 ( .A1(n_464), .A2(n_779), .B1(n_979), .B2(n_985), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_464), .A2(n_779), .B1(n_1124), .B2(n_1133), .Y(n_1164) );
OAI22xp33_ASAP7_75t_L g1513 ( .A1(n_464), .A2(n_779), .B1(n_1514), .B2(n_1515), .Y(n_1513) );
INVx6_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx5_ASAP7_75t_L g1157 ( .A(n_465), .Y(n_1157) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g611 ( .A(n_466), .Y(n_611) );
INVx4_ASAP7_75t_L g618 ( .A(n_466), .Y(n_618) );
INVx2_ASAP7_75t_SL g655 ( .A(n_466), .Y(n_655) );
INVx2_ASAP7_75t_L g781 ( .A(n_466), .Y(n_781) );
INVx1_ASAP7_75t_L g992 ( .A(n_466), .Y(n_992) );
INVx1_ASAP7_75t_L g1041 ( .A(n_466), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_468), .A2(n_700), .B1(n_714), .B2(n_724), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_468), .A2(n_1161), .B1(n_1162), .B2(n_1163), .Y(n_1160) );
INVx4_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g613 ( .A(n_470), .Y(n_613) );
INVx2_ASAP7_75t_L g1518 ( .A(n_470), .Y(n_1518) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g616 ( .A(n_471), .Y(n_616) );
BUFx2_ASAP7_75t_L g770 ( .A(n_471), .Y(n_770) );
INVx1_ASAP7_75t_L g775 ( .A(n_471), .Y(n_775) );
AND2x2_ASAP7_75t_L g540 ( .A(n_472), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g477 ( .A(n_474), .Y(n_477) );
INVx2_ASAP7_75t_L g614 ( .A(n_474), .Y(n_614) );
INVx1_ASAP7_75t_L g724 ( .A(n_474), .Y(n_724) );
INVx2_ASAP7_75t_L g799 ( .A(n_474), .Y(n_799) );
INVx4_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_475), .Y(n_662) );
BUFx4f_ASAP7_75t_L g772 ( .A(n_475), .Y(n_772) );
BUFx4f_ASAP7_75t_L g904 ( .A(n_475), .Y(n_904) );
BUFx4f_ASAP7_75t_L g1162 ( .A(n_475), .Y(n_1162) );
OAI33xp33_ASAP7_75t_L g760 ( .A1(n_478), .A2(n_719), .A3(n_761), .B1(n_766), .B2(n_773), .B3(n_778), .Y(n_760) );
OA33x2_ASAP7_75t_L g1153 ( .A1(n_478), .A2(n_535), .A3(n_1154), .B1(n_1158), .B2(n_1160), .B3(n_1164), .Y(n_1153) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
AOI33xp33_ASAP7_75t_L g533 ( .A1(n_479), .A2(n_534), .A3(n_537), .B1(n_545), .B2(n_553), .B3(n_554), .Y(n_533) );
INVx2_ASAP7_75t_L g997 ( .A(n_479), .Y(n_997) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_480), .B(n_481), .Y(n_1078) );
INVx1_ASAP7_75t_SL g1451 ( .A(n_480), .Y(n_1451) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND4xp25_ASAP7_75t_SL g487 ( .A(n_488), .B(n_505), .C(n_533), .D(n_558), .Y(n_487) );
AO21x1_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_493), .B(n_503), .Y(n_488) );
INVx2_ASAP7_75t_SL g1146 ( .A(n_491), .Y(n_1146) );
INVx1_ASAP7_75t_L g1102 ( .A(n_495), .Y(n_1102) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g1101 ( .A1(n_497), .A2(n_1082), .B1(n_1083), .B2(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1506 ( .A(n_497), .Y(n_1506) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI31xp33_ASAP7_75t_L g728 ( .A1(n_503), .A2(n_729), .A3(n_736), .B(n_739), .Y(n_728) );
CKINVDCx14_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
AOI33xp33_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_509), .A3(n_518), .B1(n_526), .B2(n_529), .B3(n_532), .Y(n_505) );
BUFx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g825 ( .A(n_507), .Y(n_825) );
AOI33xp33_ASAP7_75t_L g1426 ( .A1(n_507), .A2(n_1427), .A3(n_1428), .B1(n_1430), .B2(n_1432), .B3(n_1433), .Y(n_1426) );
INVx1_ASAP7_75t_L g1482 ( .A(n_508), .Y(n_1482) );
BUFx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g827 ( .A1(n_512), .A2(n_828), .B1(n_830), .B2(n_831), .C(n_832), .Y(n_827) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
BUFx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx8_ASAP7_75t_L g822 ( .A(n_514), .Y(n_822) );
BUFx3_ASAP7_75t_L g1127 ( .A(n_514), .Y(n_1127) );
NAND2x1p5_ASAP7_75t_L g1409 ( .A(n_514), .B(n_1410), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_516), .B(n_837), .Y(n_836) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g1096 ( .A(n_517), .Y(n_1096) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_520), .A2(n_702), .B1(n_703), .B2(n_705), .Y(n_701) );
BUFx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g530 ( .A(n_521), .Y(n_530) );
INVx3_ASAP7_75t_L g594 ( .A(n_521), .Y(n_594) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g531 ( .A(n_523), .Y(n_531) );
INVx2_ASAP7_75t_R g1431 ( .A(n_523), .Y(n_1431) );
INVx5_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g1425 ( .A(n_525), .Y(n_1425) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g1441 ( .A(n_528), .B(n_1420), .Y(n_1441) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI33xp33_ASAP7_75t_L g989 ( .A1(n_535), .A2(n_990), .A3(n_993), .B1(n_995), .B2(n_997), .B3(n_998), .Y(n_989) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_535), .A2(n_1066), .B1(n_1071), .B2(n_1078), .Y(n_1065) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI33xp33_ASAP7_75t_L g652 ( .A1(n_536), .A2(n_619), .A3(n_653), .B1(n_657), .B2(n_660), .B3(n_664), .Y(n_652) );
OAI33xp33_ASAP7_75t_L g895 ( .A1(n_536), .A2(n_619), .A3(n_896), .B1(n_899), .B2(n_902), .B3(n_906), .Y(n_895) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_SL g555 ( .A(n_539), .Y(n_555) );
INVx2_ASAP7_75t_L g863 ( .A(n_539), .Y(n_863) );
INVx2_ASAP7_75t_L g1453 ( .A(n_539), .Y(n_1453) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx6f_ASAP7_75t_L g872 ( .A(n_540), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_540), .B(n_1401), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_540), .B(n_1446), .Y(n_1459) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g557 ( .A(n_544), .Y(n_557) );
BUFx6f_ASAP7_75t_L g1077 ( .A(n_544), .Y(n_1077) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g1450 ( .A(n_547), .Y(n_1450) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g625 ( .A(n_552), .Y(n_625) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g1070 ( .A(n_557), .Y(n_1070) );
AO21x1_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B(n_570), .Y(n_558) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_567), .A2(n_629), .B1(n_801), .B2(n_802), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_567), .A2(n_679), .B1(n_882), .B2(n_883), .Y(n_881) );
BUFx3_ASAP7_75t_L g1497 ( .A(n_567), .Y(n_1497) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_568), .A2(n_774), .B1(n_776), .B2(n_777), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g1516 ( .A1(n_568), .A2(n_1517), .B1(n_1518), .B2(n_1519), .Y(n_1516) );
INVx5_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AO21x1_ASAP7_75t_L g843 ( .A1(n_570), .A2(n_844), .B(n_848), .Y(n_843) );
AOI21xp33_ASAP7_75t_L g1079 ( .A1(n_570), .A2(n_1080), .B(n_1091), .Y(n_1079) );
XOR2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_690), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
XNOR2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_649), .Y(n_574) );
XNOR2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND3x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_621), .C(n_637), .Y(n_577) );
NOR2xp33_ASAP7_75t_SL g578 ( .A(n_579), .B(n_606), .Y(n_578) );
OAI33xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .A3(n_586), .B1(n_591), .B2(n_598), .B3(n_604), .Y(n_579) );
OAI33xp33_ASAP7_75t_L g667 ( .A1(n_580), .A2(n_604), .A3(n_668), .B1(n_670), .B2(n_671), .B3(n_674), .Y(n_667) );
OAI33xp33_ASAP7_75t_L g909 ( .A1(n_580), .A2(n_604), .A3(n_910), .B1(n_911), .B2(n_912), .B3(n_914), .Y(n_909) );
OAI33xp33_ASAP7_75t_L g1026 ( .A1(n_580), .A2(n_604), .A3(n_1027), .B1(n_1030), .B2(n_1033), .B3(n_1036), .Y(n_1026) );
BUFx3_ASAP7_75t_L g1128 ( .A(n_580), .Y(n_1128) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B1(n_584), .B2(n_585), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_582), .A2(n_601), .B1(n_609), .B2(n_610), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g914 ( .A1(n_583), .A2(n_898), .B1(n_905), .B2(n_915), .Y(n_914) );
OAI22xp5_ASAP7_75t_SL g1030 ( .A1(n_583), .A2(n_585), .B1(n_1031), .B2(n_1032), .Y(n_1030) );
OAI22xp33_ASAP7_75t_L g1033 ( .A1(n_583), .A2(n_602), .B1(n_1034), .B2(n_1035), .Y(n_1033) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_585), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_589), .B2(n_590), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_587), .A2(n_592), .B1(n_613), .B2(n_614), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_588), .A2(n_590), .B1(n_658), .B2(n_665), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_588), .A2(n_901), .B1(n_908), .B2(n_913), .Y(n_912) );
OAI221xp5_ASAP7_75t_L g1111 ( .A1(n_588), .A2(n_913), .B1(n_1068), .B2(n_1112), .C(n_1113), .Y(n_1111) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_589), .A2(n_595), .B1(n_609), .B2(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B1(n_595), .B2(n_596), .Y(n_591) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g791 ( .A(n_594), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_596), .A2(n_672), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx2_ASAP7_75t_L g981 ( .A(n_597), .Y(n_981) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B1(n_602), .B2(n_603), .Y(n_598) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_599), .A2(n_654), .B1(n_661), .B2(n_669), .Y(n_668) );
OAI22xp33_ASAP7_75t_L g674 ( .A1(n_599), .A2(n_602), .B1(n_656), .B2(n_663), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g910 ( .A1(n_599), .A2(n_602), .B1(n_897), .B2(n_903), .Y(n_910) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_599), .B(n_1436), .Y(n_1435) );
INVx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g698 ( .A(n_600), .Y(n_698) );
INVx2_ASAP7_75t_L g928 ( .A(n_602), .Y(n_928) );
OAI22xp33_ASAP7_75t_L g957 ( .A1(n_602), .A2(n_698), .B1(n_958), .B2(n_959), .Y(n_957) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_602), .Y(n_976) );
BUFx6f_ASAP7_75t_L g1050 ( .A(n_602), .Y(n_1050) );
HB1xp67_ASAP7_75t_L g1530 ( .A(n_602), .Y(n_1530) );
OAI33xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .A3(n_612), .B1(n_615), .B2(n_617), .B3(n_619), .Y(n_606) );
OAI33xp33_ASAP7_75t_L g1039 ( .A1(n_607), .A2(n_1040), .A3(n_1042), .B1(n_1043), .B2(n_1045), .B3(n_1046), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_609), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_609), .A2(n_610), .B1(n_665), .B2(n_666), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_609), .A2(n_610), .B1(n_897), .B2(n_898), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_609), .A2(n_655), .B1(n_907), .B2(n_908), .Y(n_906) );
OAI22xp33_ASAP7_75t_L g1040 ( .A1(n_609), .A2(n_1031), .B1(n_1034), .B2(n_1041), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_609), .A2(n_618), .B1(n_1029), .B2(n_1038), .Y(n_1046) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_613), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_613), .A2(n_662), .B1(n_900), .B2(n_901), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_613), .A2(n_903), .B1(n_904), .B2(n_905), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_614), .A2(n_1032), .B1(n_1035), .B2(n_1044), .Y(n_1043) );
OAI22xp5_ASAP7_75t_SL g723 ( .A1(n_616), .A2(n_702), .B1(n_709), .B2(n_724), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_616), .A2(n_904), .B1(n_1028), .B2(n_1037), .Y(n_1042) );
OAI33xp33_ASAP7_75t_L g716 ( .A1(n_619), .A2(n_717), .A3(n_720), .B1(n_723), .B2(n_725), .B3(n_726), .Y(n_716) );
OAI33xp33_ASAP7_75t_L g960 ( .A1(n_619), .A2(n_719), .A3(n_961), .B1(n_964), .B2(n_965), .B3(n_966), .Y(n_960) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI33xp33_ASAP7_75t_L g861 ( .A1(n_620), .A2(n_718), .A3(n_862), .B1(n_864), .B2(n_868), .B3(n_869), .Y(n_861) );
INVx2_ASAP7_75t_L g1045 ( .A(n_620), .Y(n_1045) );
OAI31xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_632), .A3(n_635), .B(n_636), .Y(n_621) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g856 ( .A(n_624), .Y(n_856) );
INVx1_ASAP7_75t_L g855 ( .A(n_625), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_629), .B2(n_631), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_627), .A2(n_678), .B1(n_679), .B2(n_680), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g1085 ( .A1(n_627), .A2(n_629), .B1(n_1086), .B2(n_1087), .Y(n_1085) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_628), .A2(n_644), .B1(n_645), .B2(n_646), .Y(n_643) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g846 ( .A(n_633), .Y(n_846) );
BUFx3_ASAP7_75t_L g779 ( .A(n_634), .Y(n_779) );
INVx2_ASAP7_75t_SL g963 ( .A(n_634), .Y(n_963) );
OAI31xp33_ASAP7_75t_L g675 ( .A1(n_636), .A2(n_676), .A3(n_681), .B(n_682), .Y(n_675) );
INVx1_ASAP7_75t_L g754 ( .A(n_636), .Y(n_754) );
OAI31xp33_ASAP7_75t_L g797 ( .A1(n_636), .A2(n_798), .A3(n_803), .B(n_805), .Y(n_797) );
OAI31xp33_ASAP7_75t_SL g1055 ( .A1(n_636), .A2(n_1056), .A3(n_1057), .B(n_1060), .Y(n_1055) );
OAI31xp33_ASAP7_75t_SL g1137 ( .A1(n_636), .A2(n_1138), .A3(n_1139), .B(n_1143), .Y(n_1137) );
OAI31xp33_ASAP7_75t_L g1494 ( .A1(n_636), .A2(n_1495), .A3(n_1500), .B(n_1502), .Y(n_1494) );
OAI31xp33_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_641), .A3(n_647), .B(n_648), .Y(n_637) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND3xp33_ASAP7_75t_SL g835 ( .A(n_642), .B(n_836), .C(n_838), .Y(n_835) );
NAND3xp33_ASAP7_75t_SL g888 ( .A(n_642), .B(n_889), .C(n_891), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_644), .A2(n_645), .B1(n_678), .B2(n_688), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_644), .A2(n_645), .B1(n_839), .B2(n_840), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_644), .A2(n_645), .B1(n_882), .B2(n_892), .Y(n_891) );
AOI22xp33_ASAP7_75t_SL g1051 ( .A1(n_644), .A2(n_645), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
INVx1_ASAP7_75t_L g1098 ( .A(n_644), .Y(n_1098) );
INVxp67_ASAP7_75t_L g1099 ( .A(n_645), .Y(n_1099) );
OAI31xp33_ASAP7_75t_SL g684 ( .A1(n_648), .A2(n_685), .A3(n_686), .B(n_689), .Y(n_684) );
OAI31xp33_ASAP7_75t_L g1047 ( .A1(n_648), .A2(n_1048), .A3(n_1049), .B(n_1054), .Y(n_1047) );
AND3x1_ASAP7_75t_L g650 ( .A(n_651), .B(n_675), .C(n_684), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_667), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_655), .A2(n_705), .B1(n_710), .B2(n_721), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g761 ( .A1(n_655), .A2(n_762), .B1(n_763), .B2(n_765), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_655), .A2(n_952), .B1(n_956), .B2(n_962), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_659), .A2(n_666), .B1(n_672), .B2(n_673), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g1071 ( .A1(n_662), .A2(n_996), .B1(n_1072), .B2(n_1073), .C(n_1074), .Y(n_1071) );
OAI22xp5_ASAP7_75t_L g950 ( .A1(n_673), .A2(n_791), .B1(n_951), .B2(n_952), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1496 ( .A1(n_679), .A2(n_1497), .B1(n_1498), .B2(n_1499), .Y(n_1496) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B1(n_816), .B2(n_916), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_756), .B1(n_757), .B2(n_815), .Y(n_692) );
INVx1_ASAP7_75t_L g815 ( .A(n_693), .Y(n_815) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR4xp25_ASAP7_75t_L g755 ( .A(n_696), .B(n_716), .C(n_728), .D(n_744), .Y(n_755) );
BUFx4f_ASAP7_75t_SL g946 ( .A(n_698), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g720 ( .A1(n_699), .A2(n_713), .B1(n_721), .B2(n_722), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_703), .A2(n_707), .B1(n_709), .B2(n_710), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_703), .A2(n_954), .B1(n_955), .B2(n_956), .Y(n_953) );
BUFx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g1395 ( .A(n_704), .B(n_1396), .Y(n_1395) );
INVx3_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g954 ( .A(n_708), .Y(n_954) );
AND2x4_ASAP7_75t_L g1439 ( .A(n_708), .B(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g832 ( .A(n_711), .Y(n_832) );
INVx1_ASAP7_75t_L g1432 ( .A(n_711), .Y(n_1432) );
INVxp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
OAI33xp33_ASAP7_75t_L g1512 ( .A1(n_719), .A2(n_997), .A3(n_1513), .B1(n_1516), .B2(n_1520), .B3(n_1523), .Y(n_1512) );
OAI22xp33_ASAP7_75t_L g1154 ( .A1(n_721), .A2(n_1155), .B1(n_1156), .B2(n_1157), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_722), .A2(n_945), .B1(n_958), .B2(n_962), .Y(n_961) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B1(n_742), .B2(n_743), .Y(n_739) );
INVx2_ASAP7_75t_L g1152 ( .A(n_743), .Y(n_1152) );
AOI31xp67_ASAP7_75t_SL g744 ( .A1(n_745), .A2(n_749), .A3(n_752), .B(n_754), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVxp67_ASAP7_75t_SL g804 ( .A(n_748), .Y(n_804) );
INVx1_ASAP7_75t_L g1020 ( .A(n_748), .Y(n_1020) );
INVxp67_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND3xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_797), .C(n_806), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_783), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g785 ( .A1(n_762), .A2(n_776), .B1(n_786), .B2(n_789), .Y(n_785) );
INVx3_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g991 ( .A(n_764), .Y(n_991) );
INVx2_ASAP7_75t_L g1524 ( .A(n_764), .Y(n_1524) );
OAI22xp33_ASAP7_75t_L g795 ( .A1(n_765), .A2(n_777), .B1(n_786), .B2(n_796), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_771), .B2(n_772), .Y(n_766) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx4_ASAP7_75t_L g994 ( .A(n_769), .Y(n_994) );
INVx2_ASAP7_75t_L g996 ( .A(n_769), .Y(n_996) );
INVx4_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g1016 ( .A(n_772), .Y(n_1016) );
OAI221xp5_ASAP7_75t_L g1066 ( .A1(n_774), .A2(n_904), .B1(n_1067), .B2(n_1068), .C(n_1069), .Y(n_1066) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g1044 ( .A(n_775), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B1(n_781), .B2(n_782), .Y(n_778) );
OAI33xp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .A3(n_790), .B1(n_792), .B2(n_794), .B3(n_795), .Y(n_783) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g1536 ( .A(n_788), .Y(n_1536) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_794), .A2(n_1122), .B1(n_1128), .B2(n_1129), .Y(n_1121) );
OAI211xp5_ASAP7_75t_SL g1472 ( .A1(n_799), .A2(n_1473), .B(n_1474), .C(n_1477), .Y(n_1472) );
OAI31xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .A3(n_812), .B(n_814), .Y(n_806) );
OAI31xp33_ASAP7_75t_L g999 ( .A1(n_814), .A2(n_1000), .A3(n_1003), .B(n_1008), .Y(n_999) );
INVx2_ASAP7_75t_L g916 ( .A(n_816), .Y(n_916) );
XNOR2x1_ASAP7_75t_L g816 ( .A(n_817), .B(n_876), .Y(n_816) );
OR2x2_ASAP7_75t_L g817 ( .A(n_818), .B(n_857), .Y(n_817) );
INVx1_ASAP7_75t_L g859 ( .A(n_819), .Y(n_859) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_823), .B(n_826), .Y(n_819) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx3_ASAP7_75t_L g1109 ( .A(n_822), .Y(n_1109) );
INVx8_ASAP7_75t_L g1136 ( .A(n_822), .Y(n_1136) );
INVx1_ASAP7_75t_L g1532 ( .A(n_824), .Y(n_1532) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_833), .B(n_843), .Y(n_858) );
OAI31xp33_ASAP7_75t_SL g833 ( .A1(n_834), .A2(n_835), .A3(n_841), .B(n_842), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_840), .B(n_854), .Y(n_853) );
OAI31xp33_ASAP7_75t_SL g886 ( .A1(n_842), .A2(n_887), .A3(n_888), .B(n_893), .Y(n_886) );
OAI31xp33_ASAP7_75t_L g924 ( .A1(n_842), .A2(n_925), .A3(n_926), .B(n_932), .Y(n_924) );
INVx1_ASAP7_75t_L g1103 ( .A(n_842), .Y(n_1103) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_851), .Y(n_848) );
NAND3xp33_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .C(n_856), .Y(n_851) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NAND3xp33_ASAP7_75t_L g1084 ( .A(n_856), .B(n_1085), .C(n_1088), .Y(n_1084) );
OAI31xp33_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_859), .A3(n_860), .B(n_873), .Y(n_857) );
INVx1_ASAP7_75t_L g875 ( .A(n_861), .Y(n_875) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AND2x4_ASAP7_75t_L g1461 ( .A(n_866), .B(n_1446), .Y(n_1461) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx3_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
BUFx6f_ASAP7_75t_L g1478 ( .A(n_872), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
NAND3xp33_ASAP7_75t_SL g877 ( .A(n_878), .B(n_886), .C(n_894), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_883), .B(n_890), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_895), .B(n_909), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_904), .A2(n_978), .B1(n_983), .B2(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
XOR2xp5_ASAP7_75t_L g918 ( .A(n_919), .B(n_1021), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_920), .A2(n_921), .B1(n_967), .B2(n_968), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
NAND3xp33_ASAP7_75t_L g923 ( .A(n_924), .B(n_934), .C(n_942), .Y(n_923) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
OAI31xp33_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_939), .A3(n_940), .B(n_941), .Y(n_934) );
OAI31xp33_ASAP7_75t_L g1011 ( .A1(n_941), .A2(n_1012), .A3(n_1014), .B(n_1019), .Y(n_1011) );
NOR2xp33_ASAP7_75t_L g942 ( .A(n_943), .B(n_960), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_946), .B1(n_947), .B2(n_948), .Y(n_944) );
INVxp67_ASAP7_75t_SL g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g1004 ( .A(n_949), .Y(n_1004) );
INVx2_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
NAND3xp33_ASAP7_75t_L g970 ( .A(n_971), .B(n_999), .C(n_1011), .Y(n_970) );
NOR2xp33_ASAP7_75t_L g971 ( .A(n_972), .B(n_989), .Y(n_971) );
OAI22xp33_ASAP7_75t_L g990 ( .A1(n_974), .A2(n_987), .B1(n_991), .B2(n_992), .Y(n_990) );
INVx3_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g1158 ( .A1(n_996), .A2(n_1123), .B1(n_1132), .B2(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
AOI22xp5_ASAP7_75t_L g1021 ( .A1(n_1022), .A2(n_1023), .B1(n_1061), .B2(n_1166), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
AND3x1_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1047), .C(n_1055), .Y(n_1024) );
NOR2xp33_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1039), .Y(n_1025) );
BUFx3_ASAP7_75t_L g1526 ( .A(n_1041), .Y(n_1526) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1061), .Y(n_1166) );
OA22x2_ASAP7_75t_L g1061 ( .A1(n_1062), .A2(n_1117), .B1(n_1118), .B2(n_1165), .Y(n_1061) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1062), .Y(n_1165) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
NOR4xp25_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1079), .C(n_1094), .D(n_1104), .Y(n_1064) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
AND2x4_ASAP7_75t_L g1445 ( .A(n_1077), .B(n_1446), .Y(n_1445) );
HB1xp67_ASAP7_75t_L g1454 ( .A(n_1077), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1090), .Y(n_1088) );
AOI31xp33_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1100), .A3(n_1101), .B(n_1103), .Y(n_1094) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
NAND4xp75_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1137), .C(n_1144), .D(n_1153), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
BUFx2_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx2_ASAP7_75t_SL g1130 ( .A(n_1131), .Y(n_1130) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
OAI221xp5_ASAP7_75t_L g1167 ( .A1(n_1168), .A2(n_1387), .B1(n_1389), .B2(n_1483), .C(n_1487), .Y(n_1167) );
AND4x1_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1290), .C(n_1341), .D(n_1372), .Y(n_1168) );
O2A1O1Ixp33_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1226), .B(n_1260), .C(n_1269), .Y(n_1169) );
OAI221xp5_ASAP7_75t_L g1170 ( .A1(n_1171), .A2(n_1196), .B1(n_1206), .B2(n_1209), .C(n_1215), .Y(n_1170) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1171), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1171), .B(n_1366), .Y(n_1365) );
OR2x2_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1188), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1172), .B(n_1333), .Y(n_1340) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_1173), .Y(n_1172) );
NOR2xp33_ASAP7_75t_L g1228 ( .A(n_1173), .B(n_1229), .Y(n_1228) );
O2A1O1Ixp33_ASAP7_75t_L g1249 ( .A1(n_1173), .A2(n_1250), .B(n_1251), .C(n_1255), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1173), .B(n_1246), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1173), .B(n_1231), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1173), .B(n_1283), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1173), .B(n_1370), .Y(n_1369) );
INVx4_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx4_ASAP7_75t_L g1236 ( .A(n_1174), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1174), .B(n_1272), .Y(n_1271) );
NAND2xp5_ASAP7_75t_SL g1281 ( .A(n_1174), .B(n_1193), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1287 ( .A(n_1174), .B(n_1193), .Y(n_1287) );
NOR2xp33_ASAP7_75t_L g1300 ( .A(n_1174), .B(n_1301), .Y(n_1300) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_1174), .B(n_1254), .Y(n_1312) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_1174), .B(n_1324), .Y(n_1357) );
AND2x4_ASAP7_75t_SL g1174 ( .A(n_1175), .B(n_1183), .Y(n_1174) );
AND2x4_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1178), .Y(n_1176) );
AND2x6_ASAP7_75t_L g1181 ( .A(n_1177), .B(n_1182), .Y(n_1181) );
AND2x6_ASAP7_75t_L g1184 ( .A(n_1177), .B(n_1185), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1177), .B(n_1187), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1177), .B(n_1187), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1177), .B(n_1187), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1177), .B(n_1178), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1180), .Y(n_1178) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1181), .Y(n_1266) );
HB1xp67_ASAP7_75t_L g1542 ( .A(n_1182), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1188), .B(n_1237), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1193), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1189), .B(n_1212), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1189), .B(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1189), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1189), .B(n_1238), .Y(n_1248) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1189), .B(n_1212), .Y(n_1254) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1189), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1192), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1193), .B(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1193), .Y(n_1232) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1193), .B(n_1212), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1193), .B(n_1217), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1193), .B(n_1217), .Y(n_1321) );
OR2x2_ASAP7_75t_L g1381 ( .A(n_1193), .B(n_1299), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1195), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1194), .B(n_1195), .Y(n_1238) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1202), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1198), .B(n_1208), .Y(n_1207) );
INVx3_ASAP7_75t_L g1220 ( .A(n_1198), .Y(n_1220) );
NOR2xp33_ASAP7_75t_SL g1289 ( .A(n_1198), .B(n_1262), .Y(n_1289) );
A2O1A1Ixp33_ASAP7_75t_L g1290 ( .A1(n_1198), .A2(n_1291), .B(n_1313), .C(n_1326), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1198), .B(n_1202), .Y(n_1304) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1198), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1200), .Y(n_1198) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1202), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1202), .B(n_1222), .Y(n_1241) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1202), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1202), .B(n_1220), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1202), .B(n_1285), .Y(n_1298) );
OR2x2_ASAP7_75t_L g1324 ( .A(n_1202), .B(n_1223), .Y(n_1324) );
INVx2_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
OR2x2_ASAP7_75t_L g1221 ( .A(n_1203), .B(n_1222), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1205), .Y(n_1203) );
OAI222xp33_ASAP7_75t_L g1318 ( .A1(n_1206), .A2(n_1255), .B1(n_1319), .B2(n_1320), .C1(n_1322), .C2(n_1325), .Y(n_1318) );
AOI21xp33_ASAP7_75t_SL g1384 ( .A1(n_1206), .A2(n_1385), .B(n_1386), .Y(n_1384) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
NOR2xp33_ASAP7_75t_L g1275 ( .A(n_1208), .B(n_1236), .Y(n_1275) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1208), .Y(n_1371) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
O2A1O1Ixp33_ASAP7_75t_L g1335 ( .A1(n_1210), .A2(n_1336), .B(n_1337), .C(n_1338), .Y(n_1335) );
NAND2x1_ASAP7_75t_L g1386 ( .A(n_1210), .B(n_1236), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1211), .B(n_1280), .Y(n_1279) );
OAI221xp5_ASAP7_75t_L g1305 ( .A1(n_1211), .A2(n_1281), .B1(n_1306), .B2(n_1307), .C(n_1309), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1211), .B(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1211), .Y(n_1339) );
OAI21xp5_ASAP7_75t_L g1375 ( .A1(n_1211), .A2(n_1252), .B(n_1376), .Y(n_1375) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1212), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1212), .B(n_1240), .Y(n_1239) );
NAND2x1p5_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1214), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1218), .Y(n_1215) );
NAND3xp33_ASAP7_75t_L g1257 ( .A(n_1216), .B(n_1258), .C(n_1259), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1216), .B(n_1232), .Y(n_1272) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1216), .Y(n_1306) );
NOR2xp33_ASAP7_75t_L g1231 ( .A(n_1217), .B(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1221), .Y(n_1219) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1220), .B(n_1246), .Y(n_1255) );
CKINVDCx14_ASAP7_75t_R g1259 ( .A(n_1220), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1220), .B(n_1285), .Y(n_1292) );
O2A1O1Ixp33_ASAP7_75t_L g1341 ( .A1(n_1220), .A2(n_1342), .B(n_1353), .C(n_1358), .Y(n_1341) );
CKINVDCx5p33_ASAP7_75t_R g1333 ( .A(n_1221), .Y(n_1333) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1222), .Y(n_1246) );
NOR2xp33_ASAP7_75t_L g1345 ( .A(n_1222), .B(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1223), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1225), .Y(n_1223) );
A2O1A1Ixp33_ASAP7_75t_L g1226 ( .A1(n_1227), .A2(n_1233), .B(n_1241), .C(n_1242), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
HB1xp67_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1232), .B(n_1253), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1325 ( .A(n_1232), .B(n_1254), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1232), .B(n_1350), .Y(n_1349) );
OR2x2_ASAP7_75t_L g1352 ( .A(n_1232), .B(n_1239), .Y(n_1352) );
OAI211xp5_ASAP7_75t_L g1353 ( .A1(n_1233), .A2(n_1273), .B(n_1354), .C(n_1356), .Y(n_1353) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
NOR2xp33_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1237), .Y(n_1234) );
NOR2xp33_ASAP7_75t_L g1296 ( .A(n_1235), .B(n_1297), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1235), .B(n_1253), .Y(n_1309) );
CKINVDCx5p33_ASAP7_75t_R g1235 ( .A(n_1236), .Y(n_1235) );
NOR2xp33_ASAP7_75t_L g1247 ( .A(n_1236), .B(n_1248), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1236), .B(n_1285), .Y(n_1308) );
NOR2x1_ASAP7_75t_L g1350 ( .A(n_1236), .B(n_1339), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1236), .B(n_1364), .Y(n_1363) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1236), .B(n_1263), .Y(n_1383) );
NOR2xp33_ASAP7_75t_L g1355 ( .A(n_1237), .B(n_1307), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1239), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1238), .B(n_1312), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1239), .B(n_1281), .Y(n_1319) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1239), .Y(n_1364) );
CKINVDCx5p33_ASAP7_75t_R g1283 ( .A(n_1241), .Y(n_1283) );
AOI211xp5_ASAP7_75t_L g1242 ( .A1(n_1243), .A2(n_1244), .B(n_1249), .C(n_1256), .Y(n_1242) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1243), .Y(n_1273) );
A2O1A1Ixp33_ASAP7_75t_L g1342 ( .A1(n_1243), .A2(n_1343), .B(n_1344), .C(n_1348), .Y(n_1342) );
AOI32xp33_ASAP7_75t_L g1379 ( .A1(n_1243), .A2(n_1298), .A3(n_1310), .B1(n_1380), .B2(n_1382), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1247), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1245), .B(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
NOR2xp33_ASAP7_75t_L g1368 ( .A(n_1246), .B(n_1369), .Y(n_1368) );
INVxp67_ASAP7_75t_L g1370 ( .A(n_1248), .Y(n_1370) );
AOI21xp5_ASAP7_75t_L g1338 ( .A1(n_1250), .A2(n_1339), .B(n_1340), .Y(n_1338) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1253), .B(n_1280), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1253), .B(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1286 ( .A(n_1254), .B(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_1259), .B(n_1262), .Y(n_1328) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_1260), .A2(n_1359), .B1(n_1361), .B2(n_1367), .Y(n_1358) );
AOI221xp5_ASAP7_75t_L g1361 ( .A1(n_1260), .A2(n_1333), .B1(n_1362), .B2(n_1363), .C(n_1365), .Y(n_1361) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1260), .Y(n_1373) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
AOI211xp5_ASAP7_75t_SL g1302 ( .A1(n_1261), .A2(n_1303), .B(n_1305), .C(n_1310), .Y(n_1302) );
OAI21xp33_ASAP7_75t_L g1315 ( .A1(n_1261), .A2(n_1283), .B(n_1316), .Y(n_1315) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
OAI221xp5_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1265), .B1(n_1266), .B2(n_1267), .C(n_1268), .Y(n_1263) );
CKINVDCx20_ASAP7_75t_R g1388 ( .A(n_1266), .Y(n_1388) );
O2A1O1Ixp33_ASAP7_75t_SL g1269 ( .A1(n_1270), .A2(n_1273), .B(n_1274), .C(n_1288), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
OAI31xp33_ASAP7_75t_L g1367 ( .A1(n_1271), .A2(n_1345), .A3(n_1368), .B(n_1371), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1272), .B(n_1283), .Y(n_1282) );
AOI211xp5_ASAP7_75t_L g1274 ( .A1(n_1275), .A2(n_1276), .B(n_1277), .C(n_1284), .Y(n_1274) );
NAND2xp33_ASAP7_75t_SL g1277 ( .A(n_1278), .B(n_1282), .Y(n_1277) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1279), .Y(n_1343) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
OAI21xp5_ASAP7_75t_SL g1348 ( .A1(n_1283), .A2(n_1349), .B(n_1351), .Y(n_1348) );
NOR2xp33_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1286), .Y(n_1284) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1285), .Y(n_1337) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1287), .Y(n_1317) );
AOI21xp5_ASAP7_75t_L g1314 ( .A1(n_1288), .A2(n_1315), .B(n_1318), .Y(n_1314) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
A2O1A1Ixp33_ASAP7_75t_L g1291 ( .A1(n_1292), .A2(n_1293), .B(n_1295), .C(n_1302), .Y(n_1291) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
AOI21xp5_ASAP7_75t_L g1295 ( .A1(n_1296), .A2(n_1299), .B(n_1300), .Y(n_1295) );
NOR2xp33_ASAP7_75t_L g1334 ( .A(n_1297), .B(n_1319), .Y(n_1334) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
AOI221xp5_ASAP7_75t_SL g1329 ( .A1(n_1298), .A2(n_1330), .B1(n_1332), .B2(n_1333), .C(n_1334), .Y(n_1329) );
CKINVDCx14_ASAP7_75t_R g1303 ( .A(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1312), .Y(n_1331) );
INVxp67_ASAP7_75t_SL g1313 ( .A(n_1314), .Y(n_1313) );
OAI211xp5_ASAP7_75t_L g1326 ( .A1(n_1314), .A2(n_1327), .B(n_1329), .C(n_1335), .Y(n_1326) );
CKINVDCx14_ASAP7_75t_R g1320 ( .A(n_1321), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1321), .B(n_1357), .Y(n_1356) );
A2O1A1Ixp33_ASAP7_75t_L g1377 ( .A1(n_1322), .A2(n_1325), .B(n_1378), .C(n_1379), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1324), .Y(n_1322) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1324), .Y(n_1362) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1332), .Y(n_1366) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1337), .Y(n_1385) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1340), .Y(n_1376) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1349), .Y(n_1378) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVxp67_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
AOI211xp5_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1374), .B(n_1377), .C(n_1384), .Y(n_1372) );
INVxp67_ASAP7_75t_SL g1374 ( .A(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
CKINVDCx20_ASAP7_75t_R g1387 ( .A(n_1388), .Y(n_1387) );
HB1xp67_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
NAND3xp33_ASAP7_75t_SL g1391 ( .A(n_1392), .B(n_1413), .C(n_1442), .Y(n_1391) );
AOI21xp33_ASAP7_75t_L g1392 ( .A1(n_1393), .A2(n_1402), .B(n_1403), .Y(n_1392) );
INVx8_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
AND2x4_ASAP7_75t_L g1394 ( .A(n_1395), .B(n_1398), .Y(n_1394) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1396), .Y(n_1437) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1396), .Y(n_1440) );
OR2x2_ASAP7_75t_L g1398 ( .A(n_1399), .B(n_1400), .Y(n_1398) );
AND2x4_ASAP7_75t_L g1420 ( .A(n_1399), .B(n_1410), .Y(n_1420) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1401), .Y(n_1471) );
AND2x4_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1406), .Y(n_1404) );
OR2x2_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1412), .Y(n_1408) );
NOR3xp33_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1434), .C(n_1441), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1426), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g1415 ( .A1(n_1416), .A2(n_1417), .B1(n_1421), .B2(n_1422), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1420), .Y(n_1417) );
INVx3_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
AND2x4_ASAP7_75t_L g1422 ( .A(n_1420), .B(n_1423), .Y(n_1422) );
INVx2_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVxp67_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx2_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
OAI21xp5_ASAP7_75t_L g1442 ( .A1(n_1443), .A2(n_1462), .B(n_1479), .Y(n_1442) );
INVx2_ASAP7_75t_SL g1444 ( .A(n_1445), .Y(n_1444) );
AOI21xp5_ASAP7_75t_L g1447 ( .A1(n_1448), .A2(n_1452), .B(n_1455), .Y(n_1447) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_1457), .A2(n_1458), .B1(n_1460), .B2(n_1461), .Y(n_1456) );
BUFx6f_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx4_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
INVx2_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
BUFx2_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
INVx2_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
NOR2x1_ASAP7_75t_L g1469 ( .A(n_1470), .B(n_1471), .Y(n_1469) );
INVx3_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
BUFx2_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx2_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
BUFx3_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
INVxp33_ASAP7_75t_SL g1488 ( .A(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
HB1xp67_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
NAND3xp33_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1503), .C(n_1511), .Y(n_1493) );
NOR2xp33_ASAP7_75t_SL g1511 ( .A(n_1512), .B(n_1528), .Y(n_1511) );
OAI22xp5_ASAP7_75t_L g1523 ( .A1(n_1524), .A2(n_1525), .B1(n_1526), .B2(n_1527), .Y(n_1523) );
INVx2_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
BUFx3_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx2_ASAP7_75t_SL g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
OAI21xp5_ASAP7_75t_L g1541 ( .A1(n_1542), .A2(n_1543), .B(n_1544), .Y(n_1541) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
endmodule