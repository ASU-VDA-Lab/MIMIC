module fake_jpeg_15002_n_356 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_356);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_27),
.Y(n_71)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_56),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_35),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_65),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_57),
.C(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_72),
.Y(n_96)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_76),
.Y(n_98)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_20),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_55),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_53),
.B1(n_50),
.B2(n_42),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_88),
.A2(n_94),
.B1(n_61),
.B2(n_64),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_104),
.Y(n_145)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_92),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_46),
.B1(n_34),
.B2(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_111),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_62),
.A2(n_34),
.B1(n_40),
.B2(n_44),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_69),
.B(n_61),
.Y(n_126)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_27),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_39),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_68),
.B(n_34),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_117),
.B(n_32),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_71),
.A2(n_34),
.B(n_20),
.C(n_36),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_40),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_80),
.B(n_21),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_138),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_37),
.C(n_31),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_102),
.C(n_28),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_29),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_125),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_74),
.B1(n_23),
.B2(n_30),
.Y(n_129)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_91),
.Y(n_134)
);

INVx6_ASAP7_75t_SL g164 ( 
.A(n_134),
.Y(n_164)
);

OAI22x1_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_26),
.B1(n_30),
.B2(n_37),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_110),
.B(n_92),
.Y(n_151)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_74),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_149),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_31),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_70),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_88),
.Y(n_143)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_SL g193 ( 
.A(n_151),
.B(n_156),
.C(n_157),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_138),
.B(n_98),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_171),
.Y(n_181)
);

NAND2x1p5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_116),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_21),
.B(n_39),
.C(n_36),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_167),
.B(n_174),
.C(n_29),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_165),
.B(n_140),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_0),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_102),
.C(n_60),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_172),
.Y(n_179)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_104),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_59),
.C(n_101),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_126),
.B(n_145),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_176),
.A2(n_185),
.B(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_178),
.B(n_180),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_158),
.B(n_128),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_123),
.Y(n_183)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_135),
.B(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_129),
.B1(n_147),
.B2(n_121),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_153),
.B(n_141),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_175),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_146),
.B1(n_90),
.B2(n_103),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_161),
.B1(n_146),
.B2(n_90),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_170),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_130),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_194),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_121),
.B1(n_110),
.B2(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_181),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_156),
.B1(n_161),
.B2(n_160),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_224),
.B(n_201),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_167),
.B(n_174),
.C(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_218),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_209),
.B(n_214),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_210),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_SL g211 ( 
.A1(n_176),
.A2(n_151),
.B(n_173),
.C(n_168),
.Y(n_211)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_136),
.B1(n_127),
.B2(n_148),
.Y(n_247)
);

CKINVDCx12_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_172),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_184),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_136),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_170),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_217),
.B(n_190),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_222),
.B(n_187),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_151),
.B1(n_157),
.B2(n_165),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_225),
.B(n_235),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_179),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_232),
.C(n_233),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_227),
.A2(n_202),
.B(n_211),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_118),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_229),
.B(n_242),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_179),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_195),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_242),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_220),
.B(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_173),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_130),
.Y(n_239)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_241),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_159),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_249),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_59),
.C(n_118),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_209),
.C(n_221),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_247),
.A2(n_214),
.B1(n_200),
.B2(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_256),
.C(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_215),
.C(n_204),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_248),
.B(n_223),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_265),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_211),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_223),
.B1(n_211),
.B2(n_202),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_247),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_262),
.A2(n_238),
.B(n_3),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_211),
.C(n_210),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_269),
.C(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_18),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_2),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_64),
.C(n_30),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_26),
.C(n_100),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_26),
.C(n_33),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_254),
.Y(n_275)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_266),
.B(n_231),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_252),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_284),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_231),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_278),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_246),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_252),
.C(n_33),
.Y(n_294)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_108),
.B1(n_5),
.B2(n_6),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_259),
.A2(n_243),
.B(n_234),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_247),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_269),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_230),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_17),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_24),
.B(n_5),
.Y(n_296)
);

AOI21x1_ASAP7_75t_SL g288 ( 
.A1(n_267),
.A2(n_258),
.B(n_260),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_288),
.A2(n_289),
.B1(n_270),
.B2(n_271),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_2),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_304),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_299),
.C(n_301),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_277),
.Y(n_319)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_28),
.C(n_24),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_289),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_4),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_273),
.B(n_4),
.C(n_6),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_281),
.C(n_290),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_7),
.Y(n_304)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_290),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_314),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_297),
.A2(n_288),
.B(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_272),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_311),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_278),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_316),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_306),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_280),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_301),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_292),
.C(n_295),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_9),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_324),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_328),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_314),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_317),
.B(n_294),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_308),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_7),
.C(n_8),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_8),
.Y(n_337)
);

O2A1O1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_308),
.B(n_309),
.C(n_307),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_332),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_333),
.B(n_334),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_323),
.A2(n_7),
.B(n_8),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_331),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_335),
.A2(n_337),
.B1(n_321),
.B2(n_330),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_12),
.C(n_13),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_10),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_11),
.Y(n_341)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_341),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_342),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_344),
.C(n_345),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_12),
.C(n_13),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_338),
.B1(n_346),
.B2(n_336),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_350),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_347),
.B(n_341),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_352),
.B(n_351),
.CI(n_348),
.CON(n_353),
.SN(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_15),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_353),
.B1(n_16),
.B2(n_17),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_15),
.Y(n_356)
);


endmodule