module real_jpeg_11439_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_43),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_3),
.A2(n_25),
.B(n_31),
.C(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_3),
.B(n_88),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_78),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_3),
.B(n_51),
.C(n_65),
.Y(n_126)
);

NAND2x1_ASAP7_75t_SL g130 ( 
.A(n_3),
.B(n_24),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_3),
.A2(n_55),
.B(n_136),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_78),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_70),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_70),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_8),
.A2(n_34),
.B1(n_50),
.B2(n_51),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_12),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_12),
.A2(n_37),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_115),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_82),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_19),
.B(n_82),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_61),
.C(n_74),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_20),
.A2(n_21),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_40),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_41),
.C(n_48),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_30),
.B(n_35),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_23),
.A2(n_30),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2x1_ASAP7_75t_R g38 ( 
.A(n_24),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_24),
.B(n_36),
.Y(n_163)
);

AO22x1_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_26),
.A2(n_27),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_26),
.A2(n_29),
.B(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_27),
.B(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_32),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_31),
.A2(n_46),
.A3(n_89),
.B1(n_92),
.B2(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_32),
.B(n_45),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_44),
.B(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_45),
.A2(n_46),
.B1(n_88),
.B2(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_55),
.B1(n_58),
.B2(n_60),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_60),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_57),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_51),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_50),
.B(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_58),
.B1(n_60),
.B2(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_55),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_56),
.A2(n_57),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_57),
.B(n_81),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_60),
.A2(n_80),
.B(n_141),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_60),
.B(n_78),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_61),
.A2(n_74),
.B1(n_75),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_61),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_68),
.B(n_71),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_62),
.A2(n_71),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_73),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_63),
.A2(n_69),
.B1(n_72),
.B2(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_67),
.A2(n_102),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_67),
.B(n_78),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_76),
.B(n_79),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_89),
.B(n_91),
.C(n_93),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_104),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_95),
.B2(n_103),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_97),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_169),
.B(n_175),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_156),
.B(n_168),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_137),
.B(n_155),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_132),
.C(n_134),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_145),
.B(n_154),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_139),
.B(n_143),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_149),
.B(n_153),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_147),
.B(n_148),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_157),
.B(n_158),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_164),
.C(n_167),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_170),
.B(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);


endmodule