module fake_jpeg_14411_n_613 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_613);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_613;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_66),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_36),
.A2(n_38),
.B1(n_18),
.B2(n_39),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_67),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_22),
.B(n_10),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_68),
.B(n_84),
.Y(n_167)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_71),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_75),
.Y(n_180)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_77),
.Y(n_181)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_79),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_80),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_81),
.Y(n_208)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_9),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_87),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_25),
.B(n_9),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_123),
.Y(n_127)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_89),
.Y(n_174)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_91),
.Y(n_193)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_93),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_36),
.B(n_11),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_121),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_38),
.B(n_11),
.Y(n_96)
);

NAND2x1p5_ASAP7_75t_L g190 ( 
.A(n_96),
.B(n_0),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_18),
.A2(n_11),
.B1(n_15),
.B2(n_13),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_50),
.B1(n_28),
.B2(n_27),
.Y(n_132)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_98),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_8),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_103),
.B(n_106),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_26),
.B(n_12),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_18),
.Y(n_109)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_109),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_110),
.Y(n_198)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_119),
.B(n_120),
.Y(n_201)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_23),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_124),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_26),
.B(n_12),
.Y(n_124)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_46),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_125),
.A2(n_44),
.B1(n_23),
.B2(n_30),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_44),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_132),
.A2(n_138),
.B1(n_165),
.B2(n_172),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_136),
.A2(n_155),
.B1(n_170),
.B2(n_176),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_23),
.B1(n_45),
.B2(n_31),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_44),
.B1(n_43),
.B2(n_57),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_149),
.A2(n_153),
.B(n_158),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_112),
.A2(n_44),
.B1(n_43),
.B2(n_57),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_61),
.A2(n_31),
.B1(n_55),
.B2(n_45),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_157),
.B(n_190),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_21),
.B1(n_37),
.B2(n_51),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_68),
.B(n_32),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_159),
.B(n_160),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_84),
.B(n_106),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_119),
.A2(n_40),
.B1(n_37),
.B2(n_51),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_103),
.A2(n_32),
.B1(n_58),
.B2(n_33),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_122),
.A2(n_40),
.B1(n_24),
.B2(n_48),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_97),
.A2(n_29),
.B1(n_58),
.B2(n_33),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_175),
.A2(n_179),
.B1(n_183),
.B2(n_192),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_64),
.A2(n_47),
.B1(n_35),
.B2(n_29),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_83),
.B(n_35),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_178),
.B(n_206),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_78),
.A2(n_48),
.B1(n_24),
.B2(n_55),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_72),
.A2(n_47),
.B1(n_60),
.B2(n_30),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_182),
.A2(n_79),
.B(n_99),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_73),
.A2(n_60),
.B1(n_1),
.B2(n_2),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_75),
.A2(n_60),
.B1(n_13),
.B2(n_7),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_187),
.A2(n_202),
.B1(n_191),
.B2(n_169),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_82),
.A2(n_7),
.B1(n_13),
.B2(n_15),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_95),
.A2(n_16),
.B(n_15),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_15),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_77),
.A2(n_86),
.B1(n_85),
.B2(n_102),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_SL g203 ( 
.A(n_125),
.Y(n_203)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_123),
.B(n_7),
.Y(n_206)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_150),
.Y(n_209)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_210),
.B(n_219),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_167),
.A2(n_81),
.B1(n_80),
.B2(n_100),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_211),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_213),
.Y(n_330)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_215),
.Y(n_288)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_216),
.Y(n_289)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_129),
.Y(n_218)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_218),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_143),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_143),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_220),
.B(n_223),
.Y(n_301)
);

INVx11_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g304 ( 
.A(n_221),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_127),
.B(n_89),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_222),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_16),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_16),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_224),
.B(n_231),
.Y(n_295)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_225),
.Y(n_321)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_128),
.Y(n_227)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_227),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_92),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_228),
.Y(n_327)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_145),
.Y(n_229)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_229),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_230),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_16),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_133),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_233),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_154),
.Y(n_234)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_234),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_131),
.B(n_120),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_235),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_134),
.B(n_0),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_236),
.B(n_253),
.Y(n_302)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_238),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_143),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_239),
.Y(n_316)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_240),
.Y(n_299)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_140),
.Y(n_241)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_241),
.Y(n_307)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_142),
.Y(n_242)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_133),
.Y(n_243)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_162),
.Y(n_244)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_201),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_245),
.Y(n_318)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_133),
.Y(n_247)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_247),
.Y(n_293)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_152),
.Y(n_250)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_250),
.Y(n_322)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_146),
.Y(n_252)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_252),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_190),
.B(n_0),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_0),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_255),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_155),
.B(n_1),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_110),
.C(n_1),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_146),
.Y(n_258)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_258),
.Y(n_323)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_148),
.Y(n_259)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_154),
.Y(n_261)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_128),
.Y(n_262)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_262),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_147),
.Y(n_263)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_151),
.B(n_2),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_148),
.Y(n_265)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_265),
.Y(n_334)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_141),
.Y(n_266)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_193),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_267),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_201),
.B(n_2),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_279),
.Y(n_315)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_141),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_271),
.B1(n_272),
.B2(n_275),
.Y(n_286)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_174),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_156),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_274),
.A2(n_281),
.B1(n_139),
.B2(n_195),
.Y(n_319)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_161),
.Y(n_275)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_135),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_144),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_144),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_156),
.B(n_194),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_174),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_183),
.A2(n_138),
.B1(n_172),
.B2(n_165),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_217),
.A2(n_158),
.B1(n_179),
.B2(n_149),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_291),
.A2(n_292),
.B1(n_300),
.B2(n_309),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_217),
.A2(n_153),
.B1(n_137),
.B2(n_192),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_274),
.A2(n_191),
.B1(n_169),
.B2(n_208),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_214),
.A2(n_135),
.B1(n_139),
.B2(n_195),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_319),
.A2(n_320),
.B1(n_335),
.B2(n_338),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_211),
.A2(n_208),
.B1(n_171),
.B2(n_180),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_237),
.B(n_189),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_226),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_214),
.A2(n_181),
.B1(n_188),
.B2(n_171),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_248),
.A2(n_251),
.B1(n_270),
.B2(n_268),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_336),
.A2(n_198),
.B1(n_204),
.B2(n_265),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_248),
.A2(n_147),
.B1(n_180),
.B2(n_181),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_340),
.A2(n_230),
.B1(n_256),
.B2(n_273),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_342),
.A2(n_350),
.B1(n_352),
.B2(n_376),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_330),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_343),
.B(n_374),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_344),
.B(n_366),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_313),
.A2(n_226),
.B(n_268),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_345),
.A2(n_294),
.B(n_330),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_331),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_347),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_316),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_283),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_348),
.B(n_349),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_254),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_305),
.A2(n_267),
.B1(n_260),
.B2(n_188),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_313),
.A2(n_263),
.B1(n_258),
.B2(n_252),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_282),
.Y(n_353)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_254),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_359),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_275),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_355),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_290),
.A2(n_215),
.B(n_209),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_356),
.A2(n_361),
.B(n_380),
.Y(n_411)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_358),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_315),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_315),
.B(n_240),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_360),
.B(n_379),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_317),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_361),
.B(n_371),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_362),
.Y(n_401)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_333),
.Y(n_363)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_363),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_364),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_277),
.C(n_241),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_365),
.B(n_299),
.C(n_322),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_301),
.B(n_242),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_309),
.A2(n_216),
.B1(n_271),
.B2(n_259),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_368),
.A2(n_212),
.B1(n_289),
.B2(n_299),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_308),
.B(n_250),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_369),
.B(n_375),
.Y(n_412)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_370),
.Y(n_425)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_372),
.B(n_373),
.Y(n_406)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_339),
.Y(n_373)
);

O2A1O1Ixp33_ASAP7_75t_L g374 ( 
.A1(n_335),
.A2(n_221),
.B(n_334),
.C(n_287),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_294),
.B(n_280),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_302),
.A2(n_276),
.B1(n_227),
.B2(n_262),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_296),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_378),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_295),
.B(n_198),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_302),
.B(n_243),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_321),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_380),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_286),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_381),
.B(n_383),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_300),
.A2(n_334),
.B1(n_323),
.B2(n_289),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_295),
.B(n_233),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_384),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_287),
.B(n_213),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_385),
.B(n_324),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_166),
.B1(n_232),
.B2(n_204),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_386),
.A2(n_332),
.B1(n_324),
.B2(n_212),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_388),
.A2(n_420),
.B(n_381),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_328),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_407),
.C(n_413),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_359),
.B(n_298),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_396),
.B(n_407),
.Y(n_440)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_398),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_357),
.A2(n_314),
.B1(n_323),
.B2(n_298),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_424),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_342),
.A2(n_314),
.B1(n_296),
.B2(n_325),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_405),
.A2(n_421),
.B1(n_367),
.B2(n_371),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_349),
.B(n_329),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_411),
.B(n_375),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_354),
.B(n_284),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_373),
.C(n_377),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_352),
.A2(n_293),
.B1(n_306),
.B2(n_285),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_357),
.A2(n_325),
.B1(n_288),
.B2(n_284),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_385),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_367),
.A2(n_288),
.B1(n_322),
.B2(n_312),
.Y(n_424)
);

OAI32xp33_ASAP7_75t_L g427 ( 
.A1(n_402),
.A2(n_344),
.A3(n_360),
.B1(n_366),
.B2(n_383),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_427),
.B(n_432),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_428),
.A2(n_436),
.B(n_449),
.Y(n_480)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_430),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_397),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_416),
.Y(n_433)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_395),
.A2(n_345),
.B1(n_379),
.B2(n_378),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_434),
.A2(n_442),
.B1(n_456),
.B2(n_400),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_387),
.B(n_347),
.Y(n_435)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_435),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_414),
.A2(n_374),
.B(n_356),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_437),
.B(n_457),
.Y(n_466)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_399),
.Y(n_439)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_439),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_440),
.B(n_404),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_402),
.B(n_365),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_441),
.B(n_453),
.C(n_412),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_395),
.A2(n_358),
.B1(n_376),
.B2(n_341),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_443),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_406),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_447),
.Y(n_474)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_389),
.Y(n_445)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_445),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_446),
.Y(n_487)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_389),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_406),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_448),
.B(n_451),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_414),
.A2(n_411),
.B(n_388),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_415),
.C(n_405),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_423),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_452),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_396),
.B(n_413),
.C(n_394),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_419),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_458),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_397),
.A2(n_369),
.B(n_353),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_455),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_421),
.A2(n_350),
.B1(n_343),
.B2(n_386),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_419),
.B(n_372),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_397),
.A2(n_306),
.B(n_285),
.Y(n_458)
);

OAI32xp33_ASAP7_75t_L g459 ( 
.A1(n_403),
.A2(n_363),
.A3(n_364),
.B1(n_362),
.B2(n_384),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_460),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_416),
.B(n_364),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_482),
.C(n_450),
.Y(n_492)
);

BUFx5_ASAP7_75t_L g468 ( 
.A(n_439),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g503 ( 
.A(n_468),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_438),
.A2(n_417),
.B1(n_403),
.B2(n_420),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_469),
.A2(n_472),
.B1(n_479),
.B2(n_484),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_470),
.A2(n_476),
.B1(n_436),
.B2(n_426),
.Y(n_495)
);

OA22x2_ASAP7_75t_L g471 ( 
.A1(n_432),
.A2(n_438),
.B1(n_451),
.B2(n_444),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_471),
.B(n_370),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_446),
.A2(n_410),
.B1(n_390),
.B2(n_408),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_435),
.B(n_393),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_473),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_442),
.A2(n_424),
.B1(n_398),
.B2(n_392),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_449),
.A2(n_410),
.B1(n_408),
.B2(n_412),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_457),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_483),
.A2(n_486),
.B1(n_490),
.B2(n_443),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_460),
.A2(n_391),
.B1(n_393),
.B2(n_396),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_433),
.A2(n_391),
.B1(n_418),
.B2(n_401),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_437),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_425),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_492),
.B(n_504),
.C(n_506),
.Y(n_533)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_493),
.Y(n_522)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_478),
.Y(n_494)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_494),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_495),
.A2(n_496),
.B1(n_499),
.B2(n_500),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_463),
.A2(n_470),
.B1(n_488),
.B2(n_462),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_480),
.A2(n_428),
.B(n_454),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_497),
.A2(n_481),
.B(n_464),
.Y(n_529)
);

AOI21xp33_ASAP7_75t_L g498 ( 
.A1(n_487),
.A2(n_448),
.B(n_455),
.Y(n_498)
);

NAND3xp33_ASAP7_75t_L g528 ( 
.A(n_498),
.B(n_507),
.C(n_515),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_463),
.A2(n_426),
.B1(n_453),
.B2(n_434),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_488),
.A2(n_427),
.B1(n_431),
.B2(n_458),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_478),
.Y(n_501)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_501),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_462),
.A2(n_431),
.B1(n_430),
.B2(n_429),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_502),
.A2(n_510),
.B1(n_469),
.B2(n_472),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_465),
.B(n_441),
.C(n_440),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_466),
.Y(n_505)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_505),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_447),
.C(n_445),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_490),
.B(n_459),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_474),
.Y(n_508)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_508),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_474),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_517),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_475),
.A2(n_418),
.B1(n_401),
.B2(n_456),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_512),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_425),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_422),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_513),
.B(n_491),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_467),
.B(n_422),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_467),
.B(n_362),
.Y(n_516)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_516),
.Y(n_541)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_473),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_519),
.B(n_473),
.Y(n_521)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_521),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_514),
.A2(n_464),
.B1(n_475),
.B2(n_480),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_525),
.A2(n_527),
.B1(n_538),
.B2(n_510),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_514),
.A2(n_507),
.B1(n_509),
.B2(n_501),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_532),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_477),
.Y(n_534)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_534),
.Y(n_548)
);

MAJx2_ASAP7_75t_L g559 ( 
.A(n_535),
.B(n_536),
.C(n_531),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_504),
.B(n_479),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_506),
.B(n_466),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_537),
.B(n_540),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_494),
.A2(n_476),
.B1(n_485),
.B2(n_477),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_500),
.B(n_483),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_492),
.B(n_481),
.C(n_471),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_542),
.B(n_512),
.C(n_511),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_543),
.A2(n_549),
.B1(n_530),
.B2(n_520),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_546),
.B(n_558),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_527),
.A2(n_496),
.B1(n_495),
.B2(n_502),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_534),
.Y(n_550)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_550),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_533),
.B(n_499),
.C(n_513),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_551),
.B(n_552),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_526),
.A2(n_508),
.B1(n_485),
.B2(n_486),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_521),
.Y(n_553)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_553),
.Y(n_576)
);

BUFx24_ASAP7_75t_SL g554 ( 
.A(n_536),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_554),
.B(n_555),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_542),
.B(n_503),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_532),
.B(n_468),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_556),
.B(n_557),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_531),
.B(n_497),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_517),
.C(n_471),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_559),
.B(n_535),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_522),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_560),
.B(n_561),
.Y(n_564)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_541),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_548),
.A2(n_529),
.B(n_524),
.Y(n_563)
);

AOI21x1_ASAP7_75t_SL g588 ( 
.A1(n_563),
.A2(n_567),
.B(n_569),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_558),
.A2(n_523),
.B(n_539),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_568),
.A2(n_575),
.B1(n_562),
.B2(n_571),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_545),
.A2(n_520),
.B(n_530),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_547),
.A2(n_528),
.B(n_519),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_570),
.B(n_574),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_572),
.B(n_577),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_551),
.B(n_468),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_549),
.A2(n_518),
.B1(n_525),
.B2(n_515),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_556),
.A2(n_471),
.B(n_461),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_576),
.A2(n_560),
.B1(n_516),
.B2(n_544),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_578),
.B(n_580),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_566),
.B(n_546),
.C(n_544),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_563),
.A2(n_471),
.B1(n_461),
.B2(n_557),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_581),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_565),
.B(n_567),
.C(n_568),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_582),
.A2(n_589),
.B(n_579),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_571),
.B(n_572),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_307),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_569),
.A2(n_489),
.B1(n_484),
.B2(n_559),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_585),
.B(n_587),
.Y(n_591)
);

INVx6_ASAP7_75t_L g586 ( 
.A(n_573),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_582),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_577),
.A2(n_489),
.B(n_304),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_583),
.A2(n_564),
.B1(n_575),
.B2(n_304),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_592),
.B(n_594),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_587),
.A2(n_304),
.B1(n_293),
.B2(n_297),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_595),
.B(n_597),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_SL g596 ( 
.A1(n_580),
.A2(n_304),
.B(n_307),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_596),
.A2(n_589),
.B(n_579),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_598),
.B(n_585),
.Y(n_604)
);

NAND4xp25_ASAP7_75t_L g605 ( 
.A(n_599),
.B(n_603),
.C(n_588),
.D(n_601),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_593),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_600),
.B(n_604),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_591),
.A2(n_584),
.B(n_581),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_602),
.A2(n_588),
.B(n_591),
.Y(n_607)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_605),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_607),
.B(n_590),
.C(n_595),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_608),
.A2(n_606),
.B(n_586),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g611 ( 
.A(n_610),
.B(n_609),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_594),
.Y(n_612)
);

AOI321xp33_ASAP7_75t_L g613 ( 
.A1(n_612),
.A2(n_185),
.A3(n_247),
.B1(n_297),
.B2(n_312),
.C(n_598),
.Y(n_613)
);


endmodule