module fake_jpeg_2882_n_470 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_470);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_470;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_45),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_51),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_52),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_18),
.B(n_7),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_56),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_7),
.Y(n_56)
);

INVxp67_ASAP7_75t_SL g57 ( 
.A(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_18),
.B(n_7),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_30),
.B(n_8),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_76),
.Y(n_123)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_8),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_16),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_41),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_104),
.B(n_113),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_41),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_36),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_121),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_57),
.B(n_22),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_94),
.A2(n_22),
.B1(n_31),
.B2(n_24),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_133),
.B1(n_28),
.B2(n_29),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_44),
.A2(n_24),
.B1(n_31),
.B2(n_29),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_61),
.B(n_15),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_134),
.B(n_148),
.Y(n_192)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_59),
.B(n_42),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_138),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_72),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_62),
.B(n_15),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_64),
.B(n_42),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_28),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_152),
.B(n_155),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_100),
.B(n_79),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_153),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_101),
.A2(n_16),
.B1(n_52),
.B2(n_50),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_157),
.A2(n_191),
.B1(n_95),
.B2(n_126),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_108),
.B1(n_120),
.B2(n_103),
.Y(n_206)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

BUFx4f_ASAP7_75t_SL g208 ( 
.A(n_160),
.Y(n_208)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_165),
.B(n_173),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_101),
.A2(n_75),
.B1(n_82),
.B2(n_45),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_168),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_170),
.Y(n_218)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_86),
.C(n_85),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_183),
.Y(n_196)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_175),
.B(n_177),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_98),
.A2(n_47),
.B1(n_49),
.B2(n_55),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_184),
.B1(n_128),
.B2(n_133),
.Y(n_200)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_178),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g179 ( 
.A(n_97),
.B(n_84),
.Y(n_179)
);

NAND2xp33_ASAP7_75t_SL g201 ( 
.A(n_179),
.B(n_180),
.Y(n_201)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_87),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_98),
.A2(n_83),
.B(n_43),
.C(n_38),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_123),
.A2(n_53),
.B1(n_93),
.B2(n_43),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_187),
.Y(n_211)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_189),
.Y(n_223)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

NAND2xp67_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_125),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_122),
.A2(n_38),
.B1(n_8),
.B2(n_9),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_145),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_205),
.B1(n_217),
.B2(n_227),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_106),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_131),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_156),
.A2(n_124),
.B1(n_111),
.B2(n_110),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_SL g249 ( 
.A1(n_206),
.A2(n_226),
.B(n_179),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_137),
.B1(n_151),
.B2(n_129),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_212),
.A2(n_187),
.B1(n_97),
.B2(n_159),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_119),
.B1(n_112),
.B2(n_102),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_219),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_127),
.B1(n_141),
.B2(n_118),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_127),
.B1(n_126),
.B2(n_95),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_179),
.B1(n_189),
.B2(n_188),
.Y(n_251)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_186),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_232),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_169),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_198),
.A2(n_154),
.B1(n_169),
.B2(n_153),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_260)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_237),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_183),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_241),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_207),
.B(n_172),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_224),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_243),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_196),
.B(n_176),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_245),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_198),
.B(n_164),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_248),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_201),
.A2(n_179),
.B(n_153),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_247),
.A2(n_201),
.B(n_246),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_218),
.B(n_161),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_256),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_200),
.A2(n_177),
.B1(n_174),
.B2(n_141),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_255),
.B1(n_197),
.B2(n_227),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_217),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_215),
.A2(n_170),
.B1(n_167),
.B2(n_166),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_280),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_216),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_259),
.C(n_261),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_218),
.C(n_210),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_241),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_247),
.A2(n_215),
.B(n_218),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_270),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_243),
.A2(n_206),
.B(n_209),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_277),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_238),
.A2(n_244),
.B1(n_230),
.B2(n_233),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_274),
.B1(n_255),
.B2(n_226),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_238),
.A2(n_226),
.B1(n_229),
.B2(n_206),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_202),
.C(n_205),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_279),
.B1(n_234),
.B2(n_252),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_226),
.B1(n_199),
.B2(n_206),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_202),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_231),
.B(n_209),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_260),
.A2(n_251),
.B1(n_234),
.B2(n_253),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_286),
.A2(n_297),
.B1(n_300),
.B2(n_301),
.Y(n_333)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_294),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_273),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_291),
.B(n_293),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_256),
.Y(n_292)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_281),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_262),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_250),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_296),
.C(n_298),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_258),
.B(n_219),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_228),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_299),
.A2(n_302),
.B1(n_277),
.B2(n_271),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_260),
.A2(n_279),
.B1(n_282),
.B2(n_262),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_226),
.B1(n_206),
.B2(n_199),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_237),
.B1(n_197),
.B2(n_235),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_276),
.Y(n_303)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_L g305 ( 
.A1(n_270),
.A2(n_214),
.B(n_208),
.C(n_222),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_208),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_237),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_301),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_222),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_259),
.C(n_276),
.Y(n_331)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_308),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_309),
.B(n_221),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_337),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_267),
.B(n_257),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_311),
.A2(n_328),
.B(n_336),
.Y(n_357)
);

OAI22x1_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_269),
.B1(n_278),
.B2(n_283),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_313),
.A2(n_323),
.B1(n_325),
.B2(n_334),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_261),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_320),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_306),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_318),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_290),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_319),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_288),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_285),
.B(n_283),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_321),
.B(n_298),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_292),
.A2(n_265),
.B1(n_263),
.B2(n_280),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_324),
.A2(n_327),
.B1(n_296),
.B2(n_288),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_302),
.A2(n_265),
.B1(n_263),
.B2(n_280),
.Y(n_325)
);

XOR2x2_ASAP7_75t_L g326 ( 
.A(n_285),
.B(n_261),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_331),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_305),
.Y(n_327)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_284),
.A2(n_275),
.B1(n_235),
.B2(n_203),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_300),
.A2(n_220),
.B(n_275),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_355),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_328),
.A2(n_295),
.B(n_289),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_337),
.A2(n_294),
.B(n_308),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_347),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_349),
.B1(n_352),
.B2(n_356),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_307),
.Y(n_345)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_345),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_313),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_333),
.A2(n_286),
.B1(n_303),
.B2(n_275),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_350),
.A2(n_358),
.B1(n_359),
.B2(n_363),
.Y(n_382)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_330),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_353),
.Y(n_385)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_325),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_208),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_333),
.A2(n_171),
.B1(n_220),
.B2(n_178),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_320),
.B(n_160),
.C(n_162),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_360),
.B(n_346),
.C(n_355),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_221),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_331),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_322),
.A2(n_208),
.B1(n_173),
.B2(n_175),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_366),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_361),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_376),
.Y(n_401)
);

XNOR2x1_ASAP7_75t_SL g366 ( 
.A(n_362),
.B(n_311),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_368),
.C(n_373),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_329),
.C(n_321),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_348),
.B(n_323),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_372),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_329),
.C(n_310),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_338),
.C(n_342),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_378),
.C(n_379),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_335),
.Y(n_376)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_349),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_377),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_337),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_340),
.C(n_339),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_312),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_312),
.C(n_336),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_383),
.C(n_386),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_334),
.C(n_315),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_357),
.B(n_315),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_190),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_387),
.B(n_0),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_371),
.A2(n_350),
.B1(n_343),
.B2(n_352),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_385),
.A2(n_356),
.B1(n_358),
.B2(n_180),
.Y(n_390)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_390),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_370),
.A2(n_109),
.B1(n_114),
.B2(n_10),
.Y(n_392)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_382),
.Y(n_394)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_394),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_369),
.A2(n_384),
.B1(n_378),
.B2(n_379),
.Y(n_395)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_381),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_397)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_400),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_374),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_14),
.B(n_13),
.Y(n_402)
);

AOI21xp33_ASAP7_75t_L g422 ( 
.A1(n_402),
.A2(n_0),
.B(n_1),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_366),
.A2(n_14),
.B(n_11),
.Y(n_403)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_11),
.C(n_10),
.Y(n_421)
);

NAND2x1_ASAP7_75t_SL g405 ( 
.A(n_375),
.B(n_0),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_405),
.B(n_367),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_373),
.Y(n_408)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_408),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_416),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_364),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_413),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_407),
.B(n_368),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_38),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_393),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_417),
.B(n_424),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_421),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_423),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_388),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_1),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_415),
.A2(n_394),
.B(n_395),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_425),
.A2(n_405),
.B(n_406),
.Y(n_443)
);

INVx11_ASAP7_75t_L g427 ( 
.A(n_418),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_433),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_419),
.A2(n_399),
.B(n_396),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_428),
.A2(n_434),
.B(n_38),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_407),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_414),
.A2(n_396),
.B(n_401),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_409),
.A2(n_390),
.B1(n_404),
.B2(n_402),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_435),
.B(n_436),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_389),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_416),
.C(n_410),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_405),
.C(n_421),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_412),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_442),
.Y(n_451)
);

OAI21xp33_ASAP7_75t_L g440 ( 
.A1(n_429),
.A2(n_403),
.B(n_393),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_440),
.A2(n_438),
.B(n_447),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_434),
.B(n_392),
.Y(n_442)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_444),
.B(n_447),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_437),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_428),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_1),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_449),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_441),
.Y(n_450)
);

AOI211xp5_ASAP7_75t_L g459 ( 
.A1(n_450),
.A2(n_426),
.B(n_427),
.C(n_3),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_454),
.A2(n_455),
.B(n_444),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_446),
.A2(n_431),
.B(n_425),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_456),
.B(n_426),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_459),
.B(n_460),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_453),
.A2(n_1),
.B(n_2),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_461),
.B(n_462),
.C(n_457),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_451),
.A2(n_2),
.B(n_3),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_464),
.B(n_463),
.C(n_5),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_460),
.Y(n_465)
);

AOI21x1_ASAP7_75t_SL g466 ( 
.A1(n_465),
.A2(n_452),
.B(n_3),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_466),
.A2(n_467),
.B(n_2),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_5),
.C(n_6),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_5),
.Y(n_470)
);


endmodule