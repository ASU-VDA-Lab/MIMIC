module fake_jpeg_403_n_185 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_185);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_59),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_50),
.B1(n_54),
.B2(n_51),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_66),
.B1(n_23),
.B2(n_24),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_64),
.B1(n_50),
.B2(n_54),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_82),
.B1(n_74),
.B2(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_60),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_64),
.B1(n_51),
.B2(n_55),
.Y(n_82)
);

OA22x2_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_55),
.B1(n_57),
.B2(n_61),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_58),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_58),
.B1(n_57),
.B2(n_53),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_86),
.B1(n_63),
.B2(n_65),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_58),
.B1(n_57),
.B2(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_78),
.B1(n_5),
.B2(n_6),
.Y(n_111)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_77),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_100),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_93),
.B1(n_26),
.B2(n_43),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_2),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_96),
.Y(n_105)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_76),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_22),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_3),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_104),
.Y(n_107)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_3),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_4),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_118),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_121),
.B1(n_12),
.B2(n_13),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_17),
.Y(n_143)
);

NOR2x1p5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_20),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_14),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_4),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_119),
.C(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_5),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_7),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_8),
.B(n_11),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_95),
.C(n_99),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_36),
.C(n_27),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_89),
.B(n_101),
.Y(n_125)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_17),
.B(n_18),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_136),
.B1(n_140),
.B2(n_18),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_14),
.B(n_15),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_130),
.C(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_15),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_45),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_107),
.B1(n_121),
.B2(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_16),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_34),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_16),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_35),
.B1(n_41),
.B2(n_19),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_143),
.A2(n_32),
.B(n_40),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_155),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_154),
.C(n_140),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_28),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_29),
.B1(n_37),
.B2(n_39),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_136),
.C(n_134),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_147),
.C(n_151),
.Y(n_170)
);

OAI321xp33_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_130),
.A3(n_141),
.B1(n_126),
.B2(n_132),
.C(n_42),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_158),
.B1(n_153),
.B2(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_169),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_173),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_163),
.C(n_161),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_170),
.C(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_172),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_178),
.B(n_175),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_174),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_180),
.B(n_167),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_159),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_149),
.B(n_152),
.Y(n_183)
);

XOR2x2_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_149),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_160),
.Y(n_185)
);


endmodule