module fake_aes_6203_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_1), .Y(n_11) );
NOR2xp33_ASAP7_75t_R g12 ( .A(n_10), .B(n_0), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_8), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_2), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_7), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_0), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_6), .Y(n_17) );
OR2x6_ASAP7_75t_L g18 ( .A(n_12), .B(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_11), .B(n_16), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_9), .B(n_3), .Y(n_20) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_14), .A2(n_2), .B(n_3), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_18), .A2(n_12), .B1(n_15), .B2(n_4), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_18), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_19), .B(n_4), .Y(n_25) );
INVx2_ASAP7_75t_SL g26 ( .A(n_25), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
BUFx2_ASAP7_75t_L g28 ( .A(n_24), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_23), .B1(n_19), .B2(n_22), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_26), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_28), .B1(n_27), .B2(n_21), .Y(n_31) );
NOR2xp33_ASAP7_75t_R g32 ( .A(n_29), .B(n_28), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g33 ( .A(n_32), .Y(n_33) );
BUFx6f_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
XNOR2xp5_ASAP7_75t_L g36 ( .A(n_35), .B(n_27), .Y(n_36) );
OAI222xp33_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_5), .B1(n_20), .B2(n_21), .C1(n_34), .C2(n_33), .Y(n_37) );
endmodule