module fake_netlist_6_3495_n_96 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_96);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_96;

wire n_52;
wire n_91;
wire n_46;
wire n_88;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_77;
wire n_92;
wire n_42;
wire n_90;
wire n_24;
wire n_54;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_78;
wire n_84;
wire n_23;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_40;
wire n_25;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVxp67_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NAND2xp33_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_6),
.Y(n_29)
);

AND2x4_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_8),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_8),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_7),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_9),
.Y(n_44)
);

CKINVDCx11_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2x1p5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

OAI21x1_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_48),
.B(n_44),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AO31x2_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_29),
.A3(n_39),
.B(n_27),
.Y(n_53)
);

OAI21x1_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_33),
.B(n_27),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_24),
.B(n_23),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

OA21x2_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_30),
.B(n_39),
.Y(n_58)
);

OAI21x1_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_41),
.B(n_35),
.Y(n_59)
);

OAI21x1_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_55),
.B(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_52),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_52),
.Y(n_65)
);

AND2x4_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_62),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_45),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_62),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_66),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_62),
.B(n_63),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_34),
.A3(n_29),
.B1(n_31),
.B2(n_69),
.C1(n_51),
.C2(n_63),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_38),
.C(n_59),
.Y(n_78)
);

AOI221xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_63),
.B1(n_67),
.B2(n_57),
.C(n_61),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_71),
.C(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_59),
.Y(n_81)
);

NAND4xp75_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_58),
.C(n_57),
.D(n_53),
.Y(n_82)
);

NAND4xp25_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_57),
.C(n_53),
.D(n_28),
.Y(n_83)
);

NOR2xp67_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

NOR3x2_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_60),
.C(n_58),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_60),
.C(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

AOI322xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_25),
.A3(n_28),
.B1(n_83),
.B2(n_58),
.C1(n_84),
.C2(n_60),
.Y(n_89)
);

OAI211xp5_ASAP7_75t_SL g90 ( 
.A1(n_86),
.A2(n_25),
.B(n_28),
.C(n_58),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

OAI22x1_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_58),
.B1(n_25),
.B2(n_28),
.Y(n_92)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_90),
.B(n_89),
.Y(n_93)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_88),
.B(n_93),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

OR2x6_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_94),
.Y(n_96)
);


endmodule