module fake_netlist_1_9861_n_644 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_644);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_644;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
HB1xp67_ASAP7_75t_L g76 ( .A(n_55), .Y(n_76) );
CKINVDCx16_ASAP7_75t_R g77 ( .A(n_13), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_35), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_27), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_62), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_72), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_10), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_54), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_53), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_63), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_56), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_65), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_57), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_17), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_24), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_31), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_42), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_71), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_36), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_18), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_17), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_15), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_15), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_5), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_32), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_50), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_25), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_4), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_73), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_48), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_34), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_21), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_28), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_30), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_23), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_19), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_40), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_3), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_18), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_0), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_111), .B(n_0), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_77), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_108), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_111), .B(n_77), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_79), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_76), .B(n_1), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_89), .B(n_2), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_96), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_79), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_108), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_93), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_78), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_116), .B(n_4), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_93), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_89), .B(n_5), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_87), .B(n_6), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_90), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_81), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_95), .B(n_7), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_87), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_82), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_95), .B(n_7), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_87), .Y(n_146) );
NAND2xp33_ASAP7_75t_R g147 ( .A(n_103), .B(n_8), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_93), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_93), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_92), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_93), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_84), .Y(n_154) );
INVx1_ASAP7_75t_SL g155 ( .A(n_143), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_123), .B(n_83), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_152), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
BUFx4f_ASAP7_75t_L g159 ( .A(n_136), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_136), .B(n_97), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_136), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_136), .Y(n_162) );
AND2x6_ASAP7_75t_L g163 ( .A(n_136), .B(n_94), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_143), .B(n_109), .Y(n_164) );
INVx1_ASAP7_75t_SL g165 ( .A(n_131), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_152), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_127), .B(n_100), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_122), .B(n_118), .Y(n_168) );
INVx1_ASAP7_75t_SL g169 ( .A(n_131), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_122), .A2(n_117), .B1(n_114), .B2(n_97), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_122), .B(n_99), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_146), .B(n_85), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_119), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_130), .B(n_105), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_130), .B(n_105), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_146), .B(n_106), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_121), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_146), .B(n_106), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_132), .A2(n_117), .B1(n_114), .B2(n_115), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_119), .B(n_102), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_133), .B(n_113), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_133), .B(n_113), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_142), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_119), .B(n_88), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_137), .B(n_139), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_142), .Y(n_190) );
NAND2xp33_ASAP7_75t_SL g191 ( .A(n_132), .B(n_101), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_137), .B(n_102), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_121), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_121), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_139), .B(n_91), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_121), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_183), .B(n_144), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_187), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_155), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_159), .B(n_132), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_183), .B(n_144), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_183), .B(n_154), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_159), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_179), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_160), .A2(n_145), .B1(n_147), .B2(n_154), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_159), .B(n_124), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_155), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_163), .A2(n_145), .B1(n_124), .B2(n_128), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_173), .B(n_145), .Y(n_210) );
NOR3xp33_ASAP7_75t_SL g211 ( .A(n_191), .B(n_120), .C(n_147), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_179), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_183), .B(n_140), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_187), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_187), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_163), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_193), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_160), .B(n_140), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_188), .B(n_128), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_173), .B(n_128), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_160), .B(n_125), .Y(n_222) );
OR2x2_ASAP7_75t_L g223 ( .A(n_169), .B(n_120), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_157), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_157), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_163), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_189), .B(n_128), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_178), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_182), .A2(n_171), .B1(n_168), .B2(n_162), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_160), .B(n_125), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_164), .B(n_135), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_195), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_163), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_157), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_163), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_170), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_157), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_157), .Y(n_239) );
NAND2x1p5_ASAP7_75t_L g240 ( .A(n_161), .B(n_162), .Y(n_240) );
INVx1_ASAP7_75t_SL g241 ( .A(n_163), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_163), .B(n_135), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_161), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_174), .A2(n_142), .B1(n_153), .B2(n_91), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_195), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_197), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_186), .A2(n_153), .B1(n_152), .B2(n_88), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_178), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_156), .B(n_104), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_198), .Y(n_250) );
NOR2xp67_ASAP7_75t_SL g251 ( .A(n_234), .B(n_180), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_200), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_200), .B(n_167), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_222), .B(n_196), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_202), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_243), .A2(n_192), .B(n_197), .C(n_176), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_208), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_203), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_243), .A2(n_181), .B(n_190), .C(n_175), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_221), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_220), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_212), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_210), .Y(n_264) );
NAND2x2_ASAP7_75t_L g265 ( .A(n_223), .B(n_150), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_219), .A2(n_172), .B(n_180), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_205), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_222), .A2(n_138), .B1(n_184), .B2(n_190), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_213), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_206), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_229), .B(n_180), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_210), .B(n_126), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_213), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_206), .A2(n_80), .B1(n_86), .B2(n_112), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_222), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_223), .B(n_153), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_218), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_237), .B(n_9), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g279 ( .A1(n_214), .A2(n_104), .B(n_107), .C(n_110), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_222), .B(n_107), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_234), .B(n_110), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_230), .A2(n_194), .B1(n_185), .B2(n_177), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_218), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_248), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_230), .A2(n_194), .B1(n_185), .B2(n_177), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_232), .Y(n_286) );
AOI222xp33_ASAP7_75t_L g287 ( .A1(n_231), .A2(n_148), .B1(n_134), .B2(n_151), .C1(n_149), .C2(n_129), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_234), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_226), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_232), .Y(n_290) );
NOR2xp67_ASAP7_75t_SL g291 ( .A(n_226), .B(n_166), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_230), .B(n_9), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_230), .B(n_10), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_211), .B(n_11), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_242), .B(n_11), .Y(n_295) );
AO31x2_ASAP7_75t_L g296 ( .A1(n_256), .A2(n_129), .A3(n_141), .B(n_148), .Y(n_296) );
AO31x2_ASAP7_75t_L g297 ( .A1(n_256), .A2(n_129), .A3(n_141), .B(n_148), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_250), .B(n_242), .Y(n_298) );
BUFx4f_ASAP7_75t_SL g299 ( .A(n_257), .Y(n_299) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_259), .A2(n_244), .B(n_166), .Y(n_300) );
NAND2xp33_ASAP7_75t_L g301 ( .A(n_254), .B(n_241), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_252), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_271), .A2(n_233), .B(n_246), .Y(n_303) );
CKINVDCx11_ASAP7_75t_R g304 ( .A(n_265), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_262), .Y(n_305) );
BUFx12f_ASAP7_75t_L g306 ( .A(n_252), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_295), .A2(n_225), .B(n_224), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_270), .A2(n_242), .B1(n_209), .B2(n_201), .Y(n_308) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_266), .A2(n_239), .B(n_225), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_275), .B(n_204), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g311 ( .A1(n_270), .A2(n_204), .B1(n_244), .B2(n_217), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_289), .Y(n_312) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_259), .A2(n_227), .B(n_158), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_271), .A2(n_233), .B(n_245), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_263), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_267), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_269), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_272), .B(n_242), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_273), .A2(n_224), .B(n_235), .Y(n_319) );
BUFx8_ASAP7_75t_L g320 ( .A(n_255), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_258), .B(n_240), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_277), .A2(n_224), .B(n_235), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_283), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_286), .A2(n_249), .B(n_207), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_289), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_288), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_321), .B(n_260), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_320), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_302), .A2(n_264), .B1(n_274), .B2(n_294), .C(n_253), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_326), .B(n_316), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_316), .Y(n_332) );
OR2x6_ASAP7_75t_L g333 ( .A(n_321), .B(n_288), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_316), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_305), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_320), .A2(n_265), .B1(n_278), .B2(n_253), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_320), .A2(n_253), .B1(n_261), .B2(n_281), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_320), .A2(n_281), .B1(n_276), .B2(n_292), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_305), .Y(n_339) );
CKINVDCx11_ASAP7_75t_R g340 ( .A(n_306), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_317), .B(n_290), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_312), .Y(n_342) );
AOI322xp5_ASAP7_75t_L g343 ( .A1(n_315), .A2(n_268), .A3(n_280), .B1(n_293), .B2(n_247), .C1(n_281), .C2(n_12), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_317), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_323), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_299), .A2(n_204), .B1(n_284), .B2(n_245), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_326), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_323), .Y(n_348) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_306), .A2(n_204), .B1(n_217), .B2(n_236), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_312), .B(n_240), .Y(n_350) );
O2A1O1Ixp33_ASAP7_75t_L g351 ( .A1(n_311), .A2(n_279), .B(n_285), .C(n_240), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_318), .A2(n_246), .B1(n_236), .B2(n_248), .Y(n_352) );
OA21x2_ASAP7_75t_L g353 ( .A1(n_307), .A2(n_134), .B(n_141), .Y(n_353) );
A2O1A1Ixp33_ASAP7_75t_L g354 ( .A1(n_303), .A2(n_314), .B(n_325), .C(n_298), .Y(n_354) );
INVxp67_ASAP7_75t_SL g355 ( .A(n_332), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_332), .B(n_296), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_334), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_347), .Y(n_358) );
NOR2x1p5_ASAP7_75t_L g359 ( .A(n_329), .B(n_306), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_334), .B(n_296), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_331), .Y(n_361) );
AOI221x1_ASAP7_75t_SL g362 ( .A1(n_339), .A2(n_304), .B1(n_13), .B2(n_14), .C(n_16), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_335), .B(n_296), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_335), .B(n_296), .Y(n_365) );
AO21x2_ASAP7_75t_L g366 ( .A1(n_354), .A2(n_313), .B(n_314), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_345), .B(n_296), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_345), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_348), .Y(n_369) );
AND3x2_ASAP7_75t_L g370 ( .A(n_341), .B(n_327), .C(n_303), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_353), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_348), .B(n_296), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_331), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_353), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_328), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_333), .B(n_297), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_333), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_333), .B(n_297), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_341), .B(n_297), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_344), .B(n_297), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_353), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_340), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_328), .B(n_297), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_362), .A2(n_330), .B1(n_336), .B2(n_318), .C(n_328), .Y(n_385) );
OAI31xp33_ASAP7_75t_SL g386 ( .A1(n_362), .A2(n_349), .A3(n_329), .B(n_337), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_379), .B(n_297), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_361), .B(n_343), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_363), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_358), .A2(n_308), .B1(n_325), .B2(n_346), .C(n_338), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_379), .B(n_313), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_359), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_361), .B(n_342), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_355), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_371), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_373), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_363), .Y(n_398) );
AOI21xp33_ASAP7_75t_SL g399 ( .A1(n_383), .A2(n_342), .B(n_350), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_371), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_376), .A2(n_352), .B1(n_298), .B2(n_351), .C(n_350), .Y(n_401) );
INVx4_ASAP7_75t_L g402 ( .A(n_364), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_368), .B(n_327), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_371), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_368), .A2(n_310), .B1(n_313), .B2(n_134), .C(n_149), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_365), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_373), .B(n_313), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_384), .A2(n_310), .B1(n_300), .B2(n_301), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_364), .B(n_324), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_379), .B(n_300), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_356), .B(n_309), .Y(n_411) );
INVx2_ASAP7_75t_SL g412 ( .A(n_359), .Y(n_412) );
NOR3xp33_ASAP7_75t_SL g413 ( .A(n_369), .B(n_12), .C(n_16), .Y(n_413) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_377), .B(n_300), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_384), .B(n_300), .Y(n_415) );
AOI33xp33_ASAP7_75t_L g416 ( .A1(n_370), .A2(n_369), .A3(n_380), .B1(n_367), .B2(n_372), .B3(n_365), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_374), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_365), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_375), .Y(n_419) );
NOR2x1p5_ASAP7_75t_L g420 ( .A(n_376), .B(n_324), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_384), .B(n_324), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_367), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_356), .B(n_309), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_370), .B(n_287), .C(n_149), .Y(n_425) );
NOR3xp33_ASAP7_75t_L g426 ( .A(n_380), .B(n_151), .C(n_158), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_367), .B(n_324), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_389), .B(n_372), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_389), .B(n_372), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_394), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_393), .Y(n_432) );
INVx1_ASAP7_75t_SL g433 ( .A(n_394), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_395), .B(n_377), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_419), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_395), .B(n_380), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_420), .B(n_360), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_403), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_396), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_398), .B(n_357), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_398), .B(n_360), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_406), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_418), .B(n_357), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_418), .B(n_360), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_422), .B(n_356), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_425), .A2(n_378), .B1(n_355), .B2(n_381), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_396), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_422), .B(n_356), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_387), .B(n_356), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_427), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_425), .A2(n_378), .B(n_381), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_388), .B(n_366), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_416), .B(n_382), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_427), .B(n_382), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_421), .B(n_382), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g457 ( .A1(n_392), .A2(n_381), .B1(n_374), .B2(n_366), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_420), .B(n_366), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_400), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g460 ( .A(n_386), .B(n_151), .C(n_324), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_411), .B(n_366), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_400), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_404), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_404), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_387), .B(n_307), .Y(n_465) );
NOR2xp33_ASAP7_75t_SL g466 ( .A(n_392), .B(n_324), .Y(n_466) );
NOR2xp67_ASAP7_75t_L g467 ( .A(n_399), .B(n_20), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_391), .B(n_307), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_415), .B(n_322), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_411), .B(n_322), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_399), .B(n_310), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_415), .B(n_322), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_421), .B(n_319), .Y(n_473) );
AND3x2_ASAP7_75t_L g474 ( .A(n_385), .B(n_426), .C(n_412), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_412), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_417), .Y(n_476) );
NOR2xp67_ASAP7_75t_L g477 ( .A(n_402), .B(n_22), .Y(n_477) );
OR2x6_ASAP7_75t_L g478 ( .A(n_402), .B(n_319), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_391), .B(n_319), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_411), .B(n_424), .Y(n_480) );
INVx5_ASAP7_75t_L g481 ( .A(n_402), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_417), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_390), .B(n_282), .C(n_310), .D(n_248), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_481), .B(n_402), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_438), .B(n_410), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_431), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_442), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_481), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_432), .B(n_410), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_450), .B(n_424), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_443), .Y(n_491) );
AOI211xp5_ASAP7_75t_SL g492 ( .A1(n_467), .A2(n_401), .B(n_424), .C(n_411), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_481), .B(n_409), .Y(n_493) );
NOR2xp33_ASAP7_75t_SL g494 ( .A(n_481), .B(n_423), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_450), .B(n_424), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_439), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_429), .B(n_414), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_481), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_482), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_440), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_429), .B(n_414), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_453), .B(n_407), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_430), .B(n_414), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_430), .B(n_407), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_436), .B(n_423), .Y(n_505) );
AOI211xp5_ASAP7_75t_L g506 ( .A1(n_454), .A2(n_405), .B(n_413), .C(n_251), .Y(n_506) );
BUFx2_ASAP7_75t_L g507 ( .A(n_462), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_475), .Y(n_508) );
NOR3xp33_ASAP7_75t_SL g509 ( .A(n_483), .B(n_408), .C(n_29), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_444), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_445), .B(n_26), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_436), .B(n_33), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_439), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_441), .B(n_37), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_475), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_474), .A2(n_291), .B1(n_228), .B2(n_235), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_441), .B(n_38), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_446), .B(n_39), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_448), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_435), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_448), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_428), .B(n_41), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_463), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_451), .B(n_43), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_463), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_446), .B(n_44), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_464), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_433), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_449), .B(n_45), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_471), .B(n_46), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_480), .B(n_47), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_464), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_476), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_449), .B(n_49), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_465), .B(n_51), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_471), .B(n_52), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_465), .B(n_58), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_480), .B(n_461), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_509), .A2(n_477), .B(n_454), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_490), .B(n_480), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_515), .B(n_457), .Y(n_541) );
OAI22xp5_ASAP7_75t_SL g542 ( .A1(n_488), .A2(n_437), .B1(n_478), .B2(n_452), .Y(n_542) );
AOI31xp33_ASAP7_75t_L g543 ( .A1(n_492), .A2(n_447), .A3(n_437), .B(n_458), .Y(n_543) );
AOI22x1_ASAP7_75t_L g544 ( .A1(n_488), .A2(n_498), .B1(n_508), .B2(n_493), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_486), .B(n_437), .Y(n_545) );
OAI221xp5_ASAP7_75t_L g546 ( .A1(n_516), .A2(n_460), .B1(n_434), .B2(n_478), .C(n_468), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_500), .B(n_458), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_528), .B(n_458), .C(n_461), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_520), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_500), .B(n_461), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_487), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_487), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_491), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_491), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_507), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_506), .B(n_507), .C(n_510), .Y(n_556) );
OAI211xp5_ASAP7_75t_SL g557 ( .A1(n_517), .A2(n_479), .B(n_473), .C(n_455), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_490), .B(n_469), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_508), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_498), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_510), .B(n_469), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_538), .B(n_472), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_484), .A2(n_478), .B1(n_479), .B2(n_456), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_499), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_485), .B(n_472), .Y(n_565) );
OAI221xp5_ASAP7_75t_SL g566 ( .A1(n_497), .A2(n_478), .B1(n_459), .B2(n_476), .C(n_470), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g567 ( .A1(n_530), .A2(n_466), .B1(n_459), .B2(n_470), .C(n_228), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_538), .B(n_470), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_514), .A2(n_459), .B1(n_239), .B2(n_225), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_499), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_505), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_489), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_493), .A2(n_216), .B1(n_215), .B2(n_199), .Y(n_573) );
NAND2xp33_ASAP7_75t_L g574 ( .A(n_493), .B(n_59), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_496), .Y(n_575) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_531), .B(n_60), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_496), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_513), .Y(n_578) );
OAI21xp5_ASAP7_75t_L g579 ( .A1(n_514), .A2(n_216), .B(n_215), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_551), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_552), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_556), .A2(n_503), .B1(n_497), .B2(n_501), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_541), .A2(n_503), .B1(n_501), .B2(n_495), .Y(n_583) );
AOI21xp33_ASAP7_75t_L g584 ( .A1(n_543), .A2(n_522), .B(n_536), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_544), .B(n_494), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_575), .Y(n_586) );
NAND3xp33_ASAP7_75t_SL g587 ( .A(n_539), .B(n_537), .C(n_535), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_572), .B(n_495), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_550), .B(n_504), .Y(n_589) );
OAI222xp33_ASAP7_75t_L g590 ( .A1(n_541), .A2(n_537), .B1(n_535), .B2(n_534), .C1(n_518), .C2(n_529), .Y(n_590) );
OAI21xp33_ASAP7_75t_L g591 ( .A1(n_550), .A2(n_547), .B(n_545), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_555), .B(n_502), .C(n_512), .Y(n_592) );
OAI321xp33_ASAP7_75t_L g593 ( .A1(n_542), .A2(n_534), .A3(n_529), .B1(n_526), .B2(n_518), .C(n_511), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_560), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_571), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_574), .A2(n_531), .B(n_526), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_561), .B(n_504), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_553), .Y(n_598) );
NAND4xp25_ASAP7_75t_SL g599 ( .A(n_576), .B(n_524), .C(n_511), .D(n_513), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_554), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_564), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_565), .B(n_533), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_557), .A2(n_563), .B1(n_566), .B2(n_549), .C(n_545), .Y(n_603) );
OAI322xp33_ASAP7_75t_L g604 ( .A1(n_559), .A2(n_524), .A3(n_533), .B1(n_525), .B2(n_519), .C1(n_521), .C2(n_532), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_587), .A2(n_546), .B1(n_548), .B2(n_568), .Y(n_605) );
OAI21xp33_ASAP7_75t_SL g606 ( .A1(n_585), .A2(n_540), .B(n_568), .Y(n_606) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_599), .B(n_574), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_595), .B(n_570), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_580), .Y(n_609) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_603), .A2(n_567), .B(n_573), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_603), .B(n_562), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_594), .B(n_562), .Y(n_612) );
INVx2_ASAP7_75t_SL g613 ( .A(n_594), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_581), .Y(n_614) );
INVx3_ASAP7_75t_SL g615 ( .A(n_590), .Y(n_615) );
NAND2xp33_ASAP7_75t_R g616 ( .A(n_596), .B(n_531), .Y(n_616) );
OAI322xp33_ASAP7_75t_L g617 ( .A1(n_583), .A2(n_578), .A3(n_577), .B1(n_575), .B2(n_558), .C1(n_569), .C2(n_519), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g618 ( .A1(n_582), .A2(n_584), .B1(n_591), .B2(n_592), .C(n_588), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_589), .A2(n_579), .B1(n_577), .B2(n_525), .Y(n_619) );
OAI211xp5_ASAP7_75t_SL g620 ( .A1(n_610), .A2(n_602), .B(n_601), .C(n_600), .Y(n_620) );
INVxp33_ASAP7_75t_SL g621 ( .A(n_607), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_615), .B(n_597), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_613), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_611), .B(n_598), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_606), .A2(n_593), .B1(n_604), .B2(n_599), .C(n_586), .Y(n_625) );
NAND4xp25_ASAP7_75t_SL g626 ( .A(n_606), .B(n_521), .C(n_527), .D(n_523), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_616), .A2(n_532), .B1(n_527), .B2(n_523), .Y(n_627) );
AOI221x1_ASAP7_75t_L g628 ( .A1(n_619), .A2(n_239), .B1(n_238), .B2(n_66), .C(n_67), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_623), .Y(n_629) );
NAND3x1_ASAP7_75t_SL g630 ( .A(n_625), .B(n_612), .C(n_618), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_624), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_626), .B(n_622), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_621), .B(n_605), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_630), .B(n_620), .C(n_617), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_629), .Y(n_635) );
NAND4xp25_ASAP7_75t_SL g636 ( .A(n_633), .B(n_627), .C(n_628), .D(n_608), .Y(n_636) );
OAI221xp5_ASAP7_75t_L g637 ( .A1(n_634), .A2(n_632), .B1(n_631), .B2(n_614), .C(n_609), .Y(n_637) );
AOI21xp33_ASAP7_75t_SL g638 ( .A1(n_635), .A2(n_631), .B(n_64), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_637), .A2(n_636), .B1(n_238), .B2(n_216), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_638), .Y(n_640) );
AOI222xp33_ASAP7_75t_SL g641 ( .A1(n_639), .A2(n_61), .B1(n_68), .B2(n_69), .C1(n_70), .C2(n_74), .Y(n_641) );
AOI222xp33_ASAP7_75t_L g642 ( .A1(n_641), .A2(n_640), .B1(n_199), .B2(n_215), .C1(n_75), .C2(n_238), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_642), .Y(n_643) );
AOI22xp33_ASAP7_75t_SL g644 ( .A1(n_643), .A2(n_238), .B1(n_621), .B2(n_637), .Y(n_644) );
endmodule