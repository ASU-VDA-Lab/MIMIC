module fake_jpeg_2863_n_568 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_568);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_568;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_56),
.Y(n_162)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_58),
.Y(n_132)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_59),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g144 ( 
.A(n_60),
.Y(n_144)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_62),
.B(n_64),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_53),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

CKINVDCx9p33_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_72),
.Y(n_165)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_21),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_87),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_14),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_88),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_39),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_40),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_40),
.B(n_2),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_106),
.Y(n_142)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_54),
.B(n_2),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_59),
.A2(n_54),
.B1(n_50),
.B2(n_38),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_119),
.A2(n_121),
.B1(n_34),
.B2(n_20),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_55),
.A2(n_37),
.B1(n_33),
.B2(n_50),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_56),
.A2(n_37),
.B1(n_33),
.B2(n_50),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_131),
.A2(n_45),
.B1(n_30),
.B2(n_52),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_66),
.A2(n_29),
.B1(n_23),
.B2(n_34),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_134),
.A2(n_34),
.B1(n_20),
.B2(n_18),
.Y(n_193)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_38),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_65),
.B(n_38),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_80),
.Y(n_175)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_79),
.Y(n_176)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_134),
.A2(n_61),
.B1(n_82),
.B2(n_76),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_179),
.A2(n_203),
.B1(n_44),
.B2(n_36),
.Y(n_278)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_181),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_69),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_183),
.B(n_232),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_79),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_184),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_111),
.B(n_97),
.C(n_104),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_186),
.B(n_219),
.C(n_225),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_187),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_189),
.A2(n_210),
.B1(n_221),
.B2(n_223),
.Y(n_263)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_193),
.A2(n_36),
.B1(n_30),
.B2(n_35),
.Y(n_295)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_194),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_126),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_196),
.B(n_199),
.Y(n_251)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_113),
.Y(n_197)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_126),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_200),
.Y(n_273)
);

INVx4_ASAP7_75t_SL g201 ( 
.A(n_144),
.Y(n_201)
);

INVx5_ASAP7_75t_SL g253 ( 
.A(n_201),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_130),
.A2(n_33),
.B1(n_20),
.B2(n_18),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_204),
.Y(n_284)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_137),
.Y(n_207)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_133),
.A2(n_166),
.B(n_148),
.C(n_154),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_208),
.A2(n_143),
.B(n_160),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_118),
.A2(n_23),
.B1(n_29),
.B2(n_108),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_209),
.A2(n_218),
.B1(n_235),
.B2(n_41),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_130),
.A2(n_37),
.B1(n_18),
.B2(n_77),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_141),
.Y(n_211)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_211),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_213),
.Y(n_282)
);

BUFx4f_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_214),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_129),
.B(n_77),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_123),
.A2(n_29),
.B1(n_23),
.B2(n_107),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_136),
.B(n_48),
.C(n_28),
.Y(n_219)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g223 ( 
.A1(n_152),
.A2(n_177),
.B1(n_123),
.B2(n_163),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_122),
.A2(n_169),
.B1(n_117),
.B2(n_116),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_224),
.A2(n_226),
.B1(n_233),
.B2(n_41),
.Y(n_292)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_149),
.B(n_63),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_124),
.A2(n_74),
.B1(n_67),
.B2(n_63),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_120),
.Y(n_230)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_231),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_155),
.B(n_30),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_117),
.A2(n_74),
.B1(n_67),
.B2(n_95),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_165),
.B(n_28),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_240),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_120),
.A2(n_44),
.B1(n_52),
.B2(n_51),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_143),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_237),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_159),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_238),
.B(n_239),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_159),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_170),
.B(n_52),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_150),
.Y(n_241)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_172),
.Y(n_242)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_242),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_133),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_249),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_188),
.B(n_164),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_281),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_193),
.A2(n_169),
.B1(n_122),
.B2(n_173),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_255),
.A2(n_299),
.B1(n_226),
.B2(n_214),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_256),
.A2(n_218),
.B1(n_209),
.B2(n_180),
.Y(n_321)
);

BUFx24_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_262),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_184),
.B(n_145),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_276),
.Y(n_306)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_219),
.B(n_153),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_267),
.B(n_3),
.C(n_4),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_222),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_268),
.B(n_297),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_205),
.A2(n_44),
.B(n_36),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_272),
.A2(n_279),
.B(n_301),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_212),
.B(n_51),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g342 ( 
.A1(n_278),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_225),
.B(n_51),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_186),
.B(n_48),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_228),
.B(n_48),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_285),
.B(n_290),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_208),
.A2(n_45),
.B(n_41),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_286),
.A2(n_235),
.B(n_242),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_217),
.B(n_45),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_291),
.A2(n_295),
.B1(n_300),
.B2(n_214),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_292),
.Y(n_340)
);

INVx13_ASAP7_75t_L g293 ( 
.A(n_227),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_293),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_213),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_182),
.Y(n_298)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_221),
.A2(n_110),
.B1(n_60),
.B2(n_4),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_233),
.A2(n_60),
.B1(n_3),
.B2(n_4),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_215),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_302),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_237),
.B(n_2),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_305),
.A2(n_316),
.B1(n_320),
.B2(n_323),
.Y(n_391)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_307),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_254),
.B(n_197),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_308),
.B(n_313),
.C(n_339),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_271),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_260),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_310),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_195),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_246),
.B(n_198),
.C(n_185),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_273),
.Y(n_314)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_263),
.A2(n_223),
.B1(n_190),
.B2(n_202),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_236),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_263),
.A2(n_207),
.B1(n_200),
.B2(n_187),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_342),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_244),
.A2(n_178),
.B1(n_220),
.B2(n_216),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_270),
.A2(n_191),
.B1(n_181),
.B2(n_211),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_324),
.A2(n_326),
.B1(n_346),
.B2(n_282),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_267),
.A2(n_230),
.B1(n_204),
.B2(n_206),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_325),
.A2(n_343),
.B1(n_345),
.B2(n_265),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_255),
.A2(n_206),
.B1(n_4),
.B2(n_5),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_251),
.B(n_253),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_327),
.Y(n_360)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_329),
.B(n_334),
.Y(n_392)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_261),
.Y(n_330)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_267),
.B(n_3),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_347),
.Y(n_370)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_261),
.Y(n_333)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_244),
.B(n_5),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_253),
.B(n_5),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_335),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_249),
.A2(n_5),
.B(n_6),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_336),
.A2(n_344),
.B(n_262),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_256),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_338),
.A2(n_259),
.B1(n_282),
.B2(n_289),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_257),
.B(n_7),
.C(n_8),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_280),
.Y(n_341)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_278),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_343)
);

O2A1O1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_286),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_292),
.A2(n_12),
.B1(n_13),
.B2(n_279),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_279),
.A2(n_13),
.B1(n_249),
.B2(n_299),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_272),
.B(n_264),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_287),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_348),
.B(n_349),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_260),
.B(n_275),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_350),
.B(n_353),
.Y(n_383)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_250),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_257),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_354),
.B(n_394),
.C(n_395),
.Y(n_427)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_357),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_351),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_358),
.B(n_376),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_362),
.A2(n_364),
.B1(n_368),
.B2(n_371),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_363),
.A2(n_367),
.B1(n_337),
.B2(n_339),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_340),
.A2(n_243),
.B1(n_252),
.B2(n_269),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_347),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_366),
.Y(n_415)
);

AO21x2_ASAP7_75t_SL g367 ( 
.A1(n_322),
.A2(n_295),
.B(n_262),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_319),
.A2(n_269),
.B1(n_247),
.B2(n_295),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_372),
.A2(n_314),
.B1(n_312),
.B2(n_330),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_303),
.B(n_245),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_385),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_307),
.B(n_283),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_325),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_384),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_320),
.A2(n_247),
.B1(n_295),
.B2(n_277),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_381),
.A2(n_388),
.B1(n_305),
.B2(n_326),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_306),
.B(n_277),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_308),
.B(n_245),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_316),
.A2(n_271),
.B1(n_288),
.B2(n_284),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_311),
.B(n_250),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_341),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_315),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_390),
.B(n_393),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_348),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_248),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_317),
.B(n_248),
.C(n_288),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_324),
.Y(n_396)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_396),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_400),
.A2(n_404),
.B1(n_410),
.B2(n_372),
.Y(n_434)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_397),
.Y(n_401)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_401),
.Y(n_453)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_397),
.Y(n_402)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_366),
.A2(n_323),
.B1(n_346),
.B2(n_332),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_403),
.A2(n_407),
.B1(n_411),
.B2(n_412),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_382),
.A2(n_317),
.B1(n_350),
.B2(n_309),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_391),
.A2(n_331),
.B1(n_345),
.B2(n_343),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_367),
.A2(n_344),
.B(n_336),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_408),
.A2(n_420),
.B(n_395),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_426),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_382),
.A2(n_331),
.B1(n_342),
.B2(n_304),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_365),
.A2(n_329),
.B1(n_304),
.B2(n_318),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_369),
.A2(n_352),
.B1(n_337),
.B2(n_284),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_313),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_416),
.C(n_423),
.Y(n_437)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_414),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_354),
.B(n_328),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_361),
.Y(n_417)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_417),
.Y(n_439)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_361),
.Y(n_418)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_418),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_422),
.A2(n_424),
.B1(n_430),
.B2(n_388),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_379),
.B(n_353),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_365),
.A2(n_333),
.B1(n_296),
.B2(n_289),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_355),
.B(n_296),
.Y(n_425)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_425),
.Y(n_458)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_375),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_359),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_431),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_365),
.A2(n_293),
.B1(n_367),
.B2(n_374),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_355),
.B(n_389),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_385),
.B(n_370),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_433),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_370),
.B(n_360),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_434),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_379),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_435),
.B(n_457),
.Y(n_477)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_428),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_415),
.A2(n_369),
.B1(n_367),
.B2(n_371),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_400),
.A2(n_381),
.B1(n_362),
.B2(n_383),
.Y(n_442)
);

AOI21xp33_ASAP7_75t_L g444 ( 
.A1(n_398),
.A2(n_421),
.B(n_433),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_444),
.B(n_448),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_456),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_356),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g488 ( 
.A(n_447),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_398),
.A2(n_356),
.B(n_363),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_405),
.B(n_373),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_450),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_425),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_463),
.Y(n_466)
);

INVx5_ASAP7_75t_L g454 ( 
.A(n_410),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_454),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_430),
.A2(n_364),
.B1(n_368),
.B2(n_375),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_399),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_392),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_409),
.B(n_377),
.Y(n_459)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_459),
.Y(n_478)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_414),
.Y(n_461)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_461),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_413),
.B(n_392),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_462),
.B(n_406),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_423),
.B(n_432),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_416),
.B(n_378),
.C(n_386),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_464),
.B(n_404),
.C(n_411),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_476),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_434),
.A2(n_407),
.B1(n_399),
.B2(n_406),
.Y(n_470)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_470),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_464),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_471),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_472),
.B(n_462),
.Y(n_495)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_474),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_435),
.B(n_431),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_454),
.A2(n_408),
.B1(n_424),
.B2(n_412),
.Y(n_479)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_479),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_437),
.B(n_403),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_485),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_457),
.B(n_426),
.C(n_418),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_458),
.C(n_453),
.Y(n_498)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_436),
.Y(n_483)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_483),
.Y(n_494)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_436),
.Y(n_484)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_484),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_437),
.B(n_419),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_445),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_487),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_459),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_449),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_489),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_449),
.B(n_378),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_490),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_486),
.A2(n_456),
.B(n_458),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_492),
.A2(n_468),
.B(n_466),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_495),
.B(n_476),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_498),
.B(n_509),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_477),
.B(n_451),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_502),
.B(n_503),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_441),
.Y(n_503)
);

FAx1_ASAP7_75t_SL g504 ( 
.A(n_472),
.B(n_455),
.CI(n_446),
.CON(n_504),
.SN(n_504)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_504),
.A2(n_469),
.B1(n_473),
.B2(n_487),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_442),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_485),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_473),
.A2(n_438),
.B1(n_443),
.B2(n_439),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_508),
.A2(n_478),
.B1(n_483),
.B2(n_484),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_481),
.B(n_438),
.C(n_401),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_488),
.A2(n_439),
.B1(n_443),
.B2(n_417),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_510),
.A2(n_478),
.B1(n_474),
.B2(n_482),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_512),
.B(n_514),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_499),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_515),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_465),
.C(n_469),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_516),
.B(n_520),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_491),
.B(n_509),
.C(n_501),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_521),
.Y(n_532)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_507),
.Y(n_518)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_518),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_519),
.A2(n_523),
.B1(n_526),
.B2(n_492),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_469),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_502),
.B(n_467),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_525),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_479),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_506),
.A2(n_470),
.B1(n_482),
.B2(n_475),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_507),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_527),
.B(n_500),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_530),
.B(n_535),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_528),
.A2(n_497),
.B(n_499),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_531),
.A2(n_533),
.B1(n_536),
.B2(n_402),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_526),
.A2(n_506),
.B1(n_493),
.B2(n_500),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_521),
.B(n_511),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_517),
.B(n_496),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_495),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_515),
.B(n_501),
.C(n_505),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_SL g552 ( 
.A(n_538),
.B(n_541),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_514),
.B(n_522),
.C(n_524),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_532),
.B(n_522),
.C(n_525),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_543),
.B(n_544),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_511),
.C(n_512),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_538),
.B(n_520),
.C(n_508),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_546),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_539),
.A2(n_494),
.B(n_504),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_541),
.B(n_539),
.C(n_542),
.Y(n_547)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_547),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g548 ( 
.A(n_533),
.B(n_504),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_548),
.B(n_549),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_550),
.A2(n_540),
.B1(n_534),
.B2(n_530),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_556),
.B(n_558),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_551),
.A2(n_548),
.B1(n_552),
.B2(n_460),
.Y(n_558)
);

AO21x1_ASAP7_75t_L g559 ( 
.A1(n_553),
.A2(n_534),
.B(n_387),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_559),
.B(n_560),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g560 ( 
.A1(n_555),
.A2(n_460),
.B(n_387),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_561),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_563),
.A2(n_555),
.B(n_557),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_564),
.B(n_562),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_565),
.A2(n_558),
.B(n_554),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_566),
.A2(n_461),
.B(n_386),
.Y(n_567)
);

BUFx24_ASAP7_75t_SL g568 ( 
.A(n_567),
.Y(n_568)
);


endmodule