module real_aes_7032_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_312;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_729;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g456 ( .A1(n_0), .A2(n_156), .B(n_457), .C(n_460), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_1), .B(n_451), .Y(n_461) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g154 ( .A(n_3), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_4), .B(n_157), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_5), .A2(n_446), .B(n_519), .Y(n_518) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_6), .A2(n_179), .B(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_7), .A2(n_39), .B1(n_144), .B2(n_202), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_8), .A2(n_9), .B1(n_708), .B2(n_709), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_8), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_9), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_10), .B(n_179), .Y(n_187) );
AND2x6_ASAP7_75t_L g159 ( .A(n_11), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_12), .A2(n_159), .B(n_437), .C(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_13), .B(n_40), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_13), .B(n_40), .Y(n_119) );
INVx1_ASAP7_75t_L g138 ( .A(n_14), .Y(n_138) );
INVx1_ASAP7_75t_L g135 ( .A(n_15), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_16), .B(n_140), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_17), .B(n_157), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_18), .B(n_131), .Y(n_189) );
AO32x2_ASAP7_75t_L g240 ( .A1(n_19), .A2(n_130), .A3(n_173), .B1(n_179), .B2(n_241), .Y(n_240) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_20), .A2(n_30), .B1(n_121), .B2(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_20), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_21), .B(n_144), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_22), .B(n_131), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_23), .A2(n_56), .B1(n_144), .B2(n_202), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g204 ( .A1(n_24), .A2(n_81), .B1(n_140), .B2(n_144), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_25), .B(n_144), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_26), .A2(n_173), .B(n_437), .C(n_468), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_27), .A2(n_173), .B(n_437), .C(n_530), .Y(n_529) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_29), .B(n_175), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_30), .A2(n_121), .B1(n_122), .B2(n_123), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_30), .Y(n_121) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_31), .A2(n_103), .B1(n_113), .B2(n_737), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_32), .A2(n_446), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_33), .B(n_175), .Y(n_217) );
INVx2_ASAP7_75t_L g142 ( .A(n_34), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_35), .A2(n_443), .B(n_486), .C(n_487), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_36), .B(n_144), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_37), .B(n_175), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_38), .B(n_224), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_41), .B(n_466), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_42), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_43), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_44), .B(n_157), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_45), .B(n_446), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_46), .A2(n_443), .B(n_486), .C(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_47), .B(n_144), .Y(n_182) );
INVx1_ASAP7_75t_L g458 ( .A(n_48), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_49), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_50), .A2(n_90), .B1(n_202), .B2(n_203), .Y(n_201) );
INVx1_ASAP7_75t_L g511 ( .A(n_51), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_52), .B(n_144), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_53), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_54), .B(n_446), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_55), .B(n_152), .Y(n_186) );
AOI22xp33_ASAP7_75t_SL g193 ( .A1(n_57), .A2(n_61), .B1(n_140), .B2(n_144), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_58), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_59), .B(n_144), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_60), .B(n_144), .Y(n_221) );
INVx1_ASAP7_75t_L g160 ( .A(n_62), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_63), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_64), .B(n_451), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_65), .A2(n_146), .B(n_152), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_66), .B(n_144), .Y(n_155) );
INVx1_ASAP7_75t_L g134 ( .A(n_67), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_68), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_69), .B(n_157), .Y(n_489) );
AO32x2_ASAP7_75t_L g199 ( .A1(n_70), .A2(n_173), .A3(n_179), .B1(n_200), .B2(n_205), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_71), .B(n_158), .Y(n_502) );
INVx1_ASAP7_75t_L g169 ( .A(n_72), .Y(n_169) );
INVx1_ASAP7_75t_L g212 ( .A(n_73), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_74), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_75), .B(n_470), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_76), .A2(n_437), .B(n_439), .C(n_443), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_77), .B(n_140), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_78), .Y(n_520) );
INVx1_ASAP7_75t_L g112 ( .A(n_79), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_80), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_82), .B(n_202), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_83), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_84), .B(n_140), .Y(n_216) );
INVx2_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_86), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_87), .B(n_172), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_88), .B(n_140), .Y(n_183) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_89), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g117 ( .A(n_89), .B(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g428 ( .A(n_89), .Y(n_428) );
OR2x2_ASAP7_75t_L g725 ( .A(n_89), .B(n_717), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_91), .A2(n_101), .B1(n_140), .B2(n_141), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_92), .B(n_446), .Y(n_484) );
INVx1_ASAP7_75t_L g488 ( .A(n_93), .Y(n_488) );
INVxp67_ASAP7_75t_L g523 ( .A(n_94), .Y(n_523) );
XNOR2xp5_ASAP7_75t_L g726 ( .A(n_95), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_96), .B(n_140), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_97), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g440 ( .A(n_98), .Y(n_440) );
INVx1_ASAP7_75t_L g498 ( .A(n_99), .Y(n_498) );
AND2x2_ASAP7_75t_L g513 ( .A(n_100), .B(n_175), .Y(n_513) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx12_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g738 ( .A(n_106), .Y(n_738) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g118 ( .A(n_109), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO221x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_719), .B1(n_722), .B2(n_731), .C(n_733), .Y(n_113) );
OAI222xp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_707), .B1(n_710), .B2(n_714), .C1(n_715), .C2(n_718), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B1(n_426), .B2(n_429), .Y(n_115) );
INVx2_ASAP7_75t_L g712 ( .A(n_116), .Y(n_712) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g427 ( .A(n_118), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g717 ( .A(n_118), .Y(n_717) );
OAI22xp5_ASAP7_75t_SL g711 ( .A1(n_120), .A2(n_429), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_122), .A2(n_123), .B1(n_728), .B2(n_730), .Y(n_727) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR5x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_317), .C(n_375), .D(n_411), .E(n_418), .Y(n_123) );
NAND3xp33_ASAP7_75t_SL g124 ( .A(n_125), .B(n_263), .C(n_287), .Y(n_124) );
AOI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_195), .B1(n_229), .B2(n_234), .C(n_244), .Y(n_125) );
OAI21xp5_ASAP7_75t_SL g397 ( .A1(n_126), .A2(n_398), .B(n_400), .Y(n_397) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_176), .Y(n_126) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_127), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_162), .Y(n_127) );
INVx2_ASAP7_75t_L g233 ( .A(n_128), .Y(n_233) );
AND2x2_ASAP7_75t_L g246 ( .A(n_128), .B(n_178), .Y(n_246) );
AND2x2_ASAP7_75t_L g300 ( .A(n_128), .B(n_177), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_128), .B(n_163), .Y(n_315) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_136), .B(n_161), .Y(n_128) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_129), .A2(n_164), .B(n_174), .Y(n_163) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_130), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_132), .B(n_133), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_150), .B(n_159), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_143), .C(n_146), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_139), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_139), .A2(n_531), .B(n_532), .Y(n_530) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g145 ( .A(n_142), .Y(n_145) );
INVx1_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
INVx3_ASAP7_75t_L g211 ( .A(n_144), .Y(n_211) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_144), .Y(n_442) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g202 ( .A(n_145), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
AND2x6_ASAP7_75t_L g437 ( .A(n_145), .B(n_438), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_146), .A2(n_440), .B(n_441), .C(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_147), .A2(n_215), .B(n_216), .Y(n_214) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g470 ( .A(n_148), .Y(n_470) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
INVx1_ASAP7_75t_L g224 ( .A(n_149), .Y(n_224) );
INVx1_ASAP7_75t_L g438 ( .A(n_149), .Y(n_438) );
AND2x2_ASAP7_75t_L g447 ( .A(n_149), .B(n_153), .Y(n_447) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_154), .B(n_155), .C(n_156), .Y(n_150) );
O2A1O1Ixp5_ASAP7_75t_L g168 ( .A1(n_151), .A2(n_169), .B(n_170), .C(n_171), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_151), .A2(n_469), .B(n_471), .Y(n_468) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_156), .A2(n_185), .B(n_186), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_156), .A2(n_172), .B1(n_192), .B2(n_193), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_156), .A2(n_172), .B1(n_242), .B2(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_157), .A2(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_157), .A2(n_182), .B(n_183), .Y(n_181) );
O2A1O1Ixp5_ASAP7_75t_SL g210 ( .A1(n_157), .A2(n_211), .B(n_212), .C(n_213), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_157), .B(n_523), .Y(n_522) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_158), .A2(n_172), .B1(n_201), .B2(n_204), .Y(n_200) );
BUFx3_ASAP7_75t_L g173 ( .A(n_159), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_159), .A2(n_181), .B(n_184), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_159), .A2(n_210), .B(n_214), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_159), .A2(n_220), .B(n_225), .Y(n_219) );
INVx4_ASAP7_75t_SL g444 ( .A(n_159), .Y(n_444) );
AND2x4_ASAP7_75t_L g446 ( .A(n_159), .B(n_447), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g499 ( .A(n_159), .B(n_447), .Y(n_499) );
AND2x2_ASAP7_75t_L g333 ( .A(n_162), .B(n_274), .Y(n_333) );
AND2x2_ASAP7_75t_L g366 ( .A(n_162), .B(n_178), .Y(n_366) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g273 ( .A(n_163), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g286 ( .A(n_163), .B(n_178), .Y(n_286) );
AND2x2_ASAP7_75t_L g293 ( .A(n_163), .B(n_274), .Y(n_293) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_163), .Y(n_302) );
AND2x2_ASAP7_75t_L g309 ( .A(n_163), .B(n_177), .Y(n_309) );
INVx1_ASAP7_75t_L g340 ( .A(n_163), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_173), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_171), .A2(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx4_ASAP7_75t_L g459 ( .A(n_172), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g190 ( .A(n_173), .B(n_191), .C(n_194), .Y(n_190) );
INVx2_ASAP7_75t_L g205 ( .A(n_175), .Y(n_205) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_175), .A2(n_209), .B(n_217), .Y(n_208) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_175), .A2(n_219), .B(n_228), .Y(n_218) );
INVx1_ASAP7_75t_L g476 ( .A(n_175), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_175), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_175), .A2(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g316 ( .A(n_176), .Y(n_316) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_188), .Y(n_176) );
INVx2_ASAP7_75t_L g272 ( .A(n_177), .Y(n_272) );
AND2x2_ASAP7_75t_L g294 ( .A(n_177), .B(n_233), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_177), .B(n_340), .Y(n_345) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_178), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g417 ( .A(n_178), .B(n_381), .Y(n_417) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_187), .Y(n_178) );
INVx4_ASAP7_75t_L g194 ( .A(n_179), .Y(n_194) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_179), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_179), .A2(n_528), .B(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g231 ( .A(n_188), .Y(n_231) );
INVx3_ASAP7_75t_L g332 ( .A(n_188), .Y(n_332) );
OR2x2_ASAP7_75t_L g362 ( .A(n_188), .B(n_363), .Y(n_362) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_188), .B(n_272), .Y(n_388) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
INVx1_ASAP7_75t_L g275 ( .A(n_189), .Y(n_275) );
AO21x1_ASAP7_75t_L g274 ( .A1(n_191), .A2(n_194), .B(n_275), .Y(n_274) );
AO21x2_ASAP7_75t_L g434 ( .A1(n_194), .A2(n_435), .B(n_448), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_194), .B(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g451 ( .A(n_194), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_194), .B(n_492), .Y(n_491) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_194), .A2(n_497), .B(n_504), .Y(n_496) );
AOI33xp33_ASAP7_75t_L g408 ( .A1(n_195), .A2(n_246), .A3(n_260), .B1(n_332), .B2(n_409), .B3(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_206), .Y(n_196) );
OR2x2_ASAP7_75t_L g261 ( .A(n_197), .B(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_197), .B(n_258), .Y(n_320) );
OR2x2_ASAP7_75t_L g373 ( .A(n_197), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g299 ( .A(n_198), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g324 ( .A(n_198), .B(n_206), .Y(n_324) );
AND2x2_ASAP7_75t_L g391 ( .A(n_198), .B(n_236), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_198), .A2(n_291), .B(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g238 ( .A(n_199), .Y(n_238) );
INVx1_ASAP7_75t_L g251 ( .A(n_199), .Y(n_251) );
AND2x2_ASAP7_75t_L g270 ( .A(n_199), .B(n_240), .Y(n_270) );
AND2x2_ASAP7_75t_L g319 ( .A(n_199), .B(n_239), .Y(n_319) );
INVx2_ASAP7_75t_L g460 ( .A(n_203), .Y(n_460) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_203), .Y(n_490) );
INVx1_ASAP7_75t_L g473 ( .A(n_205), .Y(n_473) );
INVx2_ASAP7_75t_SL g361 ( .A(n_206), .Y(n_361) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_218), .Y(n_206) );
INVx2_ASAP7_75t_L g281 ( .A(n_207), .Y(n_281) );
INVx1_ASAP7_75t_L g412 ( .A(n_207), .Y(n_412) );
AND2x2_ASAP7_75t_L g425 ( .A(n_207), .B(n_306), .Y(n_425) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g252 ( .A(n_208), .Y(n_252) );
OR2x2_ASAP7_75t_L g258 ( .A(n_208), .B(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_208), .Y(n_269) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_218), .Y(n_236) );
AND2x2_ASAP7_75t_L g253 ( .A(n_218), .B(n_239), .Y(n_253) );
INVx1_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
INVx1_ASAP7_75t_L g266 ( .A(n_218), .Y(n_266) );
AND2x2_ASAP7_75t_L g291 ( .A(n_218), .B(n_240), .Y(n_291) );
INVx2_ASAP7_75t_L g307 ( .A(n_218), .Y(n_307) );
AND2x2_ASAP7_75t_L g400 ( .A(n_218), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_218), .B(n_281), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g255 ( .A(n_231), .Y(n_255) );
INVx1_ASAP7_75t_L g284 ( .A(n_231), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_231), .B(n_315), .Y(n_381) );
INVx1_ASAP7_75t_SL g341 ( .A(n_232), .Y(n_341) );
INVx2_ASAP7_75t_L g262 ( .A(n_233), .Y(n_262) );
AND2x2_ASAP7_75t_L g331 ( .A(n_233), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g347 ( .A(n_233), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
INVx1_ASAP7_75t_L g409 ( .A(n_235), .Y(n_409) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g264 ( .A(n_237), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g367 ( .A(n_237), .B(n_357), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_237), .A2(n_378), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g280 ( .A(n_238), .B(n_281), .Y(n_280) );
BUFx2_ASAP7_75t_L g305 ( .A(n_238), .Y(n_305) );
INVx1_ASAP7_75t_L g329 ( .A(n_238), .Y(n_329) );
OR2x2_ASAP7_75t_L g393 ( .A(n_239), .B(n_252), .Y(n_393) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_239), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g306 ( .A(n_240), .B(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_247), .B1(n_254), .B2(n_256), .Y(n_244) );
OR2x2_ASAP7_75t_L g323 ( .A(n_245), .B(n_273), .Y(n_323) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
AOI222xp33_ASAP7_75t_L g364 ( .A1(n_246), .A2(n_365), .B1(n_367), .B2(n_368), .C1(n_369), .C2(n_372), .Y(n_364) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_253), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g311 ( .A(n_250), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x2_ASAP7_75t_SL g265 ( .A(n_252), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_252), .Y(n_336) );
AND2x2_ASAP7_75t_L g384 ( .A(n_252), .B(n_253), .Y(n_384) );
INVx1_ASAP7_75t_L g402 ( .A(n_252), .Y(n_402) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g368 ( .A(n_255), .B(n_294), .Y(n_368) );
AND2x2_ASAP7_75t_L g410 ( .A(n_255), .B(n_286), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_257), .B(n_305), .Y(n_392) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_258), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g285 ( .A(n_262), .B(n_286), .Y(n_285) );
INVx3_ASAP7_75t_L g353 ( .A(n_262), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_267), .B(n_271), .C(n_276), .Y(n_263) );
INVxp67_ASAP7_75t_L g277 ( .A(n_264), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_265), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_265), .B(n_312), .Y(n_407) );
BUFx3_ASAP7_75t_L g371 ( .A(n_266), .Y(n_371) );
INVx1_ASAP7_75t_L g278 ( .A(n_267), .Y(n_278) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g297 ( .A(n_269), .B(n_291), .Y(n_297) );
INVx1_ASAP7_75t_SL g337 ( .A(n_270), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g327 ( .A(n_272), .Y(n_327) );
AND2x2_ASAP7_75t_L g350 ( .A(n_272), .B(n_333), .Y(n_350) );
INVx1_ASAP7_75t_SL g321 ( .A(n_273), .Y(n_321) );
INVx1_ASAP7_75t_L g348 ( .A(n_274), .Y(n_348) );
AOI31xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .A3(n_279), .B(n_282), .Y(n_276) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g369 ( .A(n_280), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g343 ( .A(n_281), .Y(n_343) );
BUFx2_ASAP7_75t_L g357 ( .A(n_281), .Y(n_357) );
AND2x2_ASAP7_75t_L g385 ( .A(n_281), .B(n_306), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_SL g358 ( .A(n_285), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_286), .B(n_353), .Y(n_399) );
AND2x2_ASAP7_75t_L g406 ( .A(n_286), .B(n_332), .Y(n_406) );
AOI211xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_292), .B(n_295), .C(n_310), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_292), .A2(n_319), .B1(n_320), .B2(n_321), .C(n_322), .Y(n_318) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g326 ( .A(n_293), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g363 ( .A(n_294), .Y(n_363) );
OAI32xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_298), .A3(n_301), .B1(n_303), .B2(n_308), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_297), .A2(n_350), .B(n_351), .C(n_354), .Y(n_349) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
OAI21xp5_ASAP7_75t_SL g413 ( .A1(n_305), .A2(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g374 ( .A(n_306), .Y(n_374) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_312), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g360 ( .A(n_312), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g377 ( .A(n_314), .Y(n_377) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND4xp25_ASAP7_75t_SL g317 ( .A(n_318), .B(n_330), .C(n_349), .D(n_364), .Y(n_317) );
AND2x2_ASAP7_75t_L g356 ( .A(n_319), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g378 ( .A(n_319), .B(n_371), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_321), .B(n_353), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B1(n_325), .B2(n_328), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_323), .A2(n_374), .B1(n_405), .B2(n_407), .Y(n_404) );
O2A1O1Ixp33_ASAP7_75t_L g411 ( .A1(n_323), .A2(n_412), .B(n_413), .C(n_416), .Y(n_411) );
INVx2_ASAP7_75t_L g382 ( .A(n_324), .Y(n_382) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_326), .A2(n_360), .B1(n_377), .B2(n_378), .C1(n_379), .C2(n_382), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_334), .C(n_338), .Y(n_330) );
INVx1_ASAP7_75t_L g396 ( .A(n_331), .Y(n_396) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_335), .A2(n_339), .B1(n_342), .B2(n_344), .Y(n_338) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g365 ( .A(n_347), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g423 ( .A(n_350), .Y(n_423) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_359), .B2(n_362), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_357), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g414 ( .A(n_362), .Y(n_414) );
INVx1_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_368), .Y(n_422) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND5xp2_ASAP7_75t_L g375 ( .A(n_376), .B(n_383), .C(n_397), .D(n_403), .E(n_408), .Y(n_375) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B(n_386), .C(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI31xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .A3(n_393), .B(n_394), .Y(n_389) );
INVx1_ASAP7_75t_L g415 ( .A(n_391), .Y(n_415) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI222xp33_ASAP7_75t_L g418 ( .A1(n_405), .A2(n_407), .B1(n_419), .B2(n_422), .C1(n_423), .C2(n_424), .Y(n_418) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g713 ( .A(n_426), .Y(n_713) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NOR2x2_ASAP7_75t_L g716 ( .A(n_428), .B(n_717), .Y(n_716) );
OR3x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_615), .C(n_664), .Y(n_429) );
NAND5xp2_ASAP7_75t_L g430 ( .A(n_431), .B(n_549), .C(n_578), .D(n_586), .E(n_601), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_477), .B(n_493), .C(n_533), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_462), .Y(n_432) );
AND2x2_ASAP7_75t_L g544 ( .A(n_433), .B(n_541), .Y(n_544) );
AND2x2_ASAP7_75t_L g577 ( .A(n_433), .B(n_463), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_433), .B(n_481), .Y(n_670) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_450), .Y(n_433) );
INVx2_ASAP7_75t_L g480 ( .A(n_434), .Y(n_480) );
BUFx2_ASAP7_75t_L g644 ( .A(n_434), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_445), .Y(n_435) );
INVx5_ASAP7_75t_L g455 ( .A(n_437), .Y(n_455) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_SL g453 ( .A1(n_444), .A2(n_454), .B(n_455), .C(n_456), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_444), .A2(n_455), .B(n_520), .C(n_521), .Y(n_519) );
BUFx2_ASAP7_75t_L g466 ( .A(n_446), .Y(n_466) );
AND2x2_ASAP7_75t_L g462 ( .A(n_450), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g542 ( .A(n_450), .Y(n_542) );
AND2x2_ASAP7_75t_L g628 ( .A(n_450), .B(n_541), .Y(n_628) );
AND2x2_ASAP7_75t_L g683 ( .A(n_450), .B(n_480), .Y(n_683) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_461), .Y(n_450) );
INVx2_ASAP7_75t_L g486 ( .A(n_455), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx1_ASAP7_75t_L g600 ( .A(n_462), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_462), .B(n_481), .Y(n_647) );
INVx5_ASAP7_75t_L g541 ( .A(n_463), .Y(n_541) );
AND2x4_ASAP7_75t_L g562 ( .A(n_463), .B(n_542), .Y(n_562) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_463), .Y(n_584) );
AND2x2_ASAP7_75t_L g659 ( .A(n_463), .B(n_644), .Y(n_659) );
AND2x2_ASAP7_75t_L g662 ( .A(n_463), .B(n_482), .Y(n_662) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .Y(n_463) );
AOI21xp5_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_467), .B(n_473), .Y(n_464) );
INVx2_ASAP7_75t_L g472 ( .A(n_470), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_472), .A2(n_488), .B(n_489), .C(n_490), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_472), .A2(n_490), .B(n_511), .C(n_512), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_477), .B(n_542), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_477), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
AND2x2_ASAP7_75t_L g567 ( .A(n_479), .B(n_542), .Y(n_567) );
AND2x2_ASAP7_75t_L g585 ( .A(n_479), .B(n_482), .Y(n_585) );
INVx1_ASAP7_75t_L g605 ( .A(n_479), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_479), .B(n_541), .Y(n_650) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_479), .Y(n_692) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_480), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_481), .B(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_481), .Y(n_594) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_481), .A2(n_537), .B(n_598), .C(n_600), .Y(n_597) );
AND2x2_ASAP7_75t_L g604 ( .A(n_481), .B(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g613 ( .A(n_481), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g617 ( .A(n_481), .B(n_541), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_481), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g632 ( .A(n_481), .B(n_542), .Y(n_632) );
AND2x2_ASAP7_75t_L g682 ( .A(n_481), .B(n_683), .Y(n_682) );
INVx5_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g546 ( .A(n_482), .Y(n_546) );
AND2x2_ASAP7_75t_L g587 ( .A(n_482), .B(n_540), .Y(n_587) );
AND2x2_ASAP7_75t_L g599 ( .A(n_482), .B(n_574), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_482), .B(n_628), .Y(n_646) );
OR2x6_ASAP7_75t_L g482 ( .A(n_483), .B(n_491), .Y(n_482) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_514), .Y(n_493) );
INVx1_ASAP7_75t_L g535 ( .A(n_494), .Y(n_535) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_506), .Y(n_494) );
OR2x2_ASAP7_75t_L g537 ( .A(n_495), .B(n_506), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g543 ( .A(n_495), .B(n_544), .C(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_495), .B(n_516), .Y(n_554) );
OR2x2_ASAP7_75t_L g569 ( .A(n_495), .B(n_557), .Y(n_569) );
AND2x2_ASAP7_75t_L g575 ( .A(n_495), .B(n_525), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_495), .B(n_706), .Y(n_705) );
INVx5_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_496), .B(n_516), .Y(n_572) );
AND2x2_ASAP7_75t_L g611 ( .A(n_496), .B(n_526), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_496), .B(n_525), .Y(n_639) );
OR2x2_ASAP7_75t_L g642 ( .A(n_496), .B(n_525), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_500), .Y(n_497) );
INVx5_ASAP7_75t_SL g557 ( .A(n_506), .Y(n_557) );
OR2x2_ASAP7_75t_L g563 ( .A(n_506), .B(n_515), .Y(n_563) );
AND2x2_ASAP7_75t_L g579 ( .A(n_506), .B(n_580), .Y(n_579) );
AOI321xp33_ASAP7_75t_L g586 ( .A1(n_506), .A2(n_587), .A3(n_588), .B1(n_589), .B2(n_595), .C(n_597), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_506), .B(n_514), .Y(n_596) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_506), .Y(n_609) );
OR2x2_ASAP7_75t_L g656 ( .A(n_506), .B(n_554), .Y(n_656) );
AND2x2_ASAP7_75t_L g678 ( .A(n_506), .B(n_575), .Y(n_678) );
AND2x2_ASAP7_75t_L g697 ( .A(n_506), .B(n_516), .Y(n_697) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_513), .Y(n_506) );
INVx1_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_525), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_516), .B(n_525), .Y(n_538) );
AND2x2_ASAP7_75t_L g547 ( .A(n_516), .B(n_548), .Y(n_547) );
INVx3_ASAP7_75t_L g574 ( .A(n_516), .Y(n_574) );
AND2x2_ASAP7_75t_L g580 ( .A(n_516), .B(n_575), .Y(n_580) );
INVxp67_ASAP7_75t_L g610 ( .A(n_516), .Y(n_610) );
OR2x2_ASAP7_75t_L g652 ( .A(n_516), .B(n_557), .Y(n_652) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_524), .Y(n_516) );
OR2x2_ASAP7_75t_L g534 ( .A(n_525), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_SL g548 ( .A(n_525), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_525), .B(n_537), .Y(n_581) );
AND2x2_ASAP7_75t_L g630 ( .A(n_525), .B(n_574), .Y(n_630) );
AND2x2_ASAP7_75t_L g668 ( .A(n_525), .B(n_557), .Y(n_668) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_526), .B(n_557), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_536), .B(n_539), .C(n_543), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_534), .A2(n_536), .B1(n_661), .B2(n_663), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_536), .A2(n_559), .B1(n_614), .B2(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_SL g688 ( .A(n_537), .Y(n_688) );
INVx1_ASAP7_75t_SL g588 ( .A(n_538), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_540), .B(n_560), .Y(n_590) );
AOI222xp33_ASAP7_75t_L g601 ( .A1(n_540), .A2(n_581), .B1(n_588), .B2(n_602), .C1(n_606), .C2(n_612), .Y(n_601) );
AND2x2_ASAP7_75t_L g691 ( .A(n_540), .B(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx2_ASAP7_75t_L g566 ( .A(n_541), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_541), .B(n_561), .Y(n_636) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_541), .Y(n_673) );
AND2x2_ASAP7_75t_L g676 ( .A(n_541), .B(n_585), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_541), .B(n_692), .Y(n_702) );
INVx1_ASAP7_75t_L g593 ( .A(n_542), .Y(n_593) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_542), .Y(n_621) );
O2A1O1Ixp33_ASAP7_75t_L g684 ( .A1(n_544), .A2(n_685), .B(n_686), .C(n_689), .Y(n_684) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_546), .B(n_608), .C(n_611), .Y(n_607) );
OR2x2_ASAP7_75t_L g635 ( .A(n_546), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_546), .B(n_562), .Y(n_663) );
OR2x2_ASAP7_75t_L g568 ( .A(n_548), .B(n_569), .Y(n_568) );
AOI211xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_552), .B(n_558), .C(n_570), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_551), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g657 ( .A(n_552), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_553), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g571 ( .A(n_556), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_557), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g625 ( .A(n_557), .B(n_575), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_557), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_557), .B(n_574), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_563), .B1(n_564), .B2(n_568), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_560), .B(n_632), .Y(n_631) );
BUFx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_562), .B(n_604), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g626 ( .A1(n_563), .A2(n_627), .B1(n_629), .B2(n_631), .C(n_633), .Y(n_626) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
AND2x2_ASAP7_75t_L g681 ( .A(n_566), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g694 ( .A(n_566), .B(n_683), .Y(n_694) );
INVx1_ASAP7_75t_L g614 ( .A(n_567), .Y(n_614) );
INVx1_ASAP7_75t_L g685 ( .A(n_568), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_569), .A2(n_652), .B(n_675), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .B(n_576), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI21xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_581), .B(n_582), .Y(n_578) );
INVx1_ASAP7_75t_L g618 ( .A(n_579), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_580), .A2(n_666), .B1(n_669), .B2(n_671), .C(n_674), .Y(n_665) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_588), .A2(n_678), .B1(n_679), .B2(n_681), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g654 ( .A(n_590), .Y(n_654) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp67_ASAP7_75t_SL g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g658 ( .A(n_594), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g623 ( .A(n_599), .Y(n_623) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_604), .B(n_628), .Y(n_680) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_610), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g696 ( .A(n_611), .B(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_L g703 ( .A(n_611), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI211xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_618), .B(n_619), .C(n_653), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI211xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_622), .B(n_626), .C(n_645), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g706 ( .A(n_630), .Y(n_706) );
AND2x2_ASAP7_75t_L g643 ( .A(n_632), .B(n_644), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_637), .B1(n_641), .B2(n_643), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OR2x2_ASAP7_75t_L g651 ( .A(n_639), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g704 ( .A(n_640), .Y(n_704) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI31xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .A3(n_648), .B(n_651), .Y(n_645) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B(n_657), .C(n_660), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
CKINVDCx16_ASAP7_75t_R g661 ( .A(n_662), .Y(n_661) );
NAND5xp2_ASAP7_75t_L g664 ( .A(n_665), .B(n_677), .C(n_684), .D(n_698), .E(n_701), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_676), .A2(n_702), .B1(n_703), .B2(n_705), .Y(n_701) );
INVx1_ASAP7_75t_SL g700 ( .A(n_678), .Y(n_700) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_693), .B(n_695), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g714 ( .A(n_707), .Y(n_714) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
BUFx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_SL g732 ( .A(n_720), .Y(n_732) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
BUFx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g736 ( .A(n_725), .Y(n_736) );
INVx1_ASAP7_75t_L g730 ( .A(n_728), .Y(n_730) );
BUFx3_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
endmodule