module fake_jpeg_14423_n_297 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_297);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_19),
.B(n_18),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_27),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_56),
.Y(n_80)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_54),
.Y(n_81)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_38),
.B1(n_34),
.B2(n_36),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_34),
.B1(n_36),
.B2(n_35),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_38),
.B1(n_34),
.B2(n_36),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_34),
.B1(n_36),
.B2(n_35),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_38),
.B1(n_35),
.B2(n_39),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_68),
.A2(n_97),
.B1(n_100),
.B2(n_24),
.Y(n_134)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_39),
.B1(n_35),
.B2(n_21),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_84),
.B1(n_87),
.B2(n_89),
.Y(n_104)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_39),
.B1(n_21),
.B2(n_37),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_39),
.B1(n_40),
.B2(n_37),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_40),
.B1(n_33),
.B2(n_32),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_45),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_22),
.C(n_25),
.Y(n_108)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_47),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_20),
.B1(n_24),
.B2(n_3),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_29),
.B1(n_22),
.B2(n_25),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_22),
.B1(n_25),
.B2(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_101),
.B(n_102),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_4),
.Y(n_153)
);

NAND2x1_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_25),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_116),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_16),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_113),
.B(n_119),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_122),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_65),
.B(n_20),
.C(n_24),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_71),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_20),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_0),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_89),
.B(n_14),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_66),
.B(n_3),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_3),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_132),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_84),
.A2(n_4),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_131),
.A2(n_78),
.B(n_61),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_97),
.Y(n_132)
);

BUFx4f_ASAP7_75t_SL g133 ( 
.A(n_81),
.Y(n_133)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_67),
.B1(n_62),
.B2(n_82),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_157),
.B1(n_158),
.B2(n_139),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_163),
.Y(n_178)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_142),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_64),
.B1(n_68),
.B2(n_82),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_165),
.B1(n_129),
.B2(n_120),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_99),
.B1(n_69),
.B2(n_77),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_147),
.A2(n_153),
.B(n_161),
.Y(n_170)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_123),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_109),
.B1(n_104),
.B2(n_127),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_63),
.B1(n_96),
.B2(n_8),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_63),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_112),
.A2(n_5),
.B(n_7),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_5),
.B(n_8),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_118),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_125),
.B(n_105),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_168),
.B(n_144),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_125),
.B(n_103),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_171),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_129),
.B1(n_117),
.B2(n_121),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_172),
.A2(n_144),
.B1(n_162),
.B2(n_140),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_114),
.C(n_117),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_195),
.C(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_128),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_175),
.B(n_181),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_176),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_123),
.B1(n_11),
.B2(n_12),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_180),
.B1(n_187),
.B2(n_151),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_179),
.B(n_158),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_13),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_10),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_161),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_149),
.B(n_11),
.Y(n_186)
);

NOR2x1_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_160),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_139),
.A2(n_147),
.B1(n_135),
.B2(n_141),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_137),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_140),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_191),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_137),
.B(n_136),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_163),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_194),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_152),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_170),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_189),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_204),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_217),
.B1(n_218),
.B2(n_167),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_203),
.B(n_197),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_168),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_206),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_136),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_209),
.C(n_213),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_175),
.C(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_215),
.B(n_166),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_190),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_212),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_138),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_178),
.A2(n_164),
.B(n_150),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_178),
.A2(n_142),
.B1(n_155),
.B2(n_169),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_172),
.A2(n_171),
.B1(n_183),
.B2(n_176),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_229),
.C(n_213),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_228),
.B1(n_218),
.B2(n_202),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_186),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_176),
.B1(n_177),
.B2(n_185),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_176),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_209),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_174),
.B(n_184),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_200),
.Y(n_236)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_238),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_244),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_224),
.B(n_208),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_252),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_231),
.B(n_205),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_247),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_220),
.B(n_196),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_192),
.Y(n_250)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_202),
.B1(n_227),
.B2(n_232),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_203),
.C(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_237),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_242),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_240),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_230),
.B(n_236),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_262),
.B(n_249),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_265),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_234),
.B(n_217),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_245),
.C(n_233),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_228),
.B1(n_211),
.B2(n_216),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_249),
.B1(n_253),
.B2(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_262),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_263),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_272),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_204),
.C(n_223),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_239),
.B1(n_221),
.B2(n_166),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_279),
.Y(n_283)
);

OAI221xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.C(n_259),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_277),
.A2(n_268),
.B(n_266),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_286),
.B(n_258),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_273),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_174),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_270),
.C(n_260),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_290),
.B(n_291),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_280),
.B1(n_275),
.B2(n_258),
.Y(n_291)
);

INVxp33_ASAP7_75t_SL g293 ( 
.A(n_288),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_289),
.B(n_283),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_292),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_295),
.B(n_260),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_192),
.B1(n_193),
.B2(n_289),
.Y(n_297)
);


endmodule