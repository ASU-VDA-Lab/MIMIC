module fake_jpeg_27650_n_139 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_139);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_68),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_45),
.B1(n_50),
.B2(n_43),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_73),
.B1(n_55),
.B2(n_36),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_42),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_54),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_75),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_36),
.C(n_40),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_46),
.Y(n_90)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_38),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_44),
.B1(n_39),
.B2(n_2),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_1),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_37),
.B1(n_3),
.B2(n_4),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_94),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_82),
.B1(n_91),
.B2(n_6),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_84),
.B(n_79),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_103),
.B(n_85),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_105),
.B(n_9),
.Y(n_118)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_110),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_85),
.C(n_90),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_98),
.B1(n_102),
.B2(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_101),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_118),
.Y(n_123)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_10),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_11),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_17),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_127),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_129),
.Y(n_132)
);

OAI221xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_128),
.B1(n_123),
.B2(n_112),
.C(n_122),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_123),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_21),
.B1(n_25),
.B2(n_29),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_113),
.C(n_31),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_30),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_32),
.Y(n_139)
);


endmodule