module fake_jpeg_12071_n_484 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_484);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_484;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_58),
.B(n_60),
.Y(n_121)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_59),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_20),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_61),
.B(n_65),
.Y(n_138)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_64),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_23),
.B(n_17),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_68),
.Y(n_126)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_71),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_25),
.B(n_16),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_72),
.B(n_79),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_75),
.Y(n_173)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_77),
.Y(n_146)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

INVx2_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_90),
.Y(n_127)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_32),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_86),
.B(n_87),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_32),
.B(n_36),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_88),
.Y(n_189)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_89),
.Y(n_195)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_33),
.B(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_93),
.Y(n_139)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_36),
.B(n_38),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_95),
.Y(n_186)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx5_ASAP7_75t_SL g184 ( 
.A(n_96),
.Y(n_184)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

BUFx4f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_38),
.B(n_2),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_110),
.Y(n_136)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_105),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_43),
.B(n_4),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_19),
.Y(n_109)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_43),
.B(n_15),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_19),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_111),
.B(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_115),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_114),
.B(n_116),
.Y(n_191)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_19),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_117),
.Y(n_176)
);

INVx6_ASAP7_75t_SL g118 ( 
.A(n_48),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_118),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_44),
.B(n_4),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_5),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_39),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_56),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_67),
.A2(n_21),
.B1(n_52),
.B2(n_44),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_125),
.A2(n_131),
.B1(n_133),
.B2(n_141),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_74),
.A2(n_21),
.B1(n_52),
.B2(n_55),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_81),
.A2(n_21),
.B1(n_52),
.B2(n_55),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_91),
.A2(n_52),
.B1(n_54),
.B2(n_39),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_135),
.A2(n_140),
.B1(n_154),
.B2(n_158),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_84),
.A2(n_54),
.B1(n_39),
.B2(n_51),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_51),
.B1(n_41),
.B2(n_42),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_142),
.A2(n_183),
.B(n_196),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_35),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_145),
.B(n_148),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_59),
.B(n_50),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_62),
.A2(n_30),
.B1(n_56),
.B2(n_40),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_151),
.A2(n_152),
.B1(n_162),
.B2(n_171),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_85),
.A2(n_30),
.B1(n_40),
.B2(n_56),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_54),
.B1(n_42),
.B2(n_40),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_49),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_155),
.B(n_165),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_116),
.A2(n_42),
.B1(n_47),
.B2(n_45),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_63),
.A2(n_30),
.B1(n_42),
.B2(n_48),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_163),
.B(n_136),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_109),
.A2(n_49),
.B1(n_47),
.B2(n_45),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_164),
.A2(n_168),
.B1(n_190),
.B2(n_192),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_5),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_117),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_75),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_64),
.B(n_6),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_178),
.B(n_187),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_71),
.A2(n_15),
.B1(n_11),
.B2(n_13),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_97),
.B(n_6),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_95),
.A2(n_77),
.B1(n_120),
.B2(n_96),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_146),
.B1(n_185),
.B2(n_186),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_77),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_98),
.A2(n_13),
.B1(n_14),
.B2(n_73),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_100),
.A2(n_14),
.B1(n_107),
.B2(n_98),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_100),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_197),
.B(n_202),
.C(n_238),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_107),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_198),
.Y(n_273)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_199),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_73),
.B1(n_136),
.B2(n_172),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_200),
.A2(n_223),
.B1(n_232),
.B2(n_235),
.Y(n_272)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_145),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_203),
.B(n_208),
.Y(n_267)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_205),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_139),
.B(n_121),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_207),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_138),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_126),
.B(n_137),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_209),
.B(n_211),
.Y(n_274)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_210),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_127),
.B(n_167),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_212),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_213),
.B(n_216),
.Y(n_281)
);

NAND2x1_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_172),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_214),
.A2(n_220),
.B(n_197),
.Y(n_276)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_195),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_184),
.A2(n_172),
.B(n_136),
.C(n_189),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_224),
.Y(n_271)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_142),
.B1(n_150),
.B2(n_166),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_218),
.A2(n_229),
.B1(n_248),
.B2(n_259),
.Y(n_270)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_219),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_134),
.A2(n_173),
.B1(n_186),
.B2(n_159),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_222),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_166),
.B1(n_156),
.B2(n_150),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_225),
.B(n_231),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_124),
.B1(n_129),
.B2(n_128),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_227),
.A2(n_233),
.B1(n_258),
.B2(n_217),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_132),
.A2(n_146),
.B1(n_134),
.B2(n_173),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_159),
.B(n_174),
.Y(n_231)
);

AO21x1_ASAP7_75t_SL g232 ( 
.A1(n_196),
.A2(n_183),
.B(n_146),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_124),
.A2(n_129),
.B1(n_156),
.B2(n_128),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_174),
.B(n_147),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_234),
.B(n_236),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_170),
.B1(n_175),
.B2(n_179),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_177),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_147),
.B(n_176),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_237),
.B(n_239),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_170),
.B(n_175),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_177),
.Y(n_239)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_132),
.Y(n_240)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_123),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_241),
.B(n_246),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_179),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_244),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_130),
.Y(n_243)
);

BUFx4f_ASAP7_75t_SL g311 ( 
.A(n_243),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_153),
.B(n_130),
.Y(n_244)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_153),
.Y(n_245)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_123),
.B(n_180),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_180),
.A2(n_144),
.B1(n_181),
.B2(n_161),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_144),
.B(n_161),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_249),
.B(n_254),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_130),
.Y(n_250)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_250),
.Y(n_298)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_143),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_251),
.B(n_256),
.Y(n_303)
);

AOI32xp33_ASAP7_75t_L g252 ( 
.A1(n_148),
.A2(n_155),
.A3(n_165),
.B1(n_145),
.B2(n_137),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_221),
.Y(n_285)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_130),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_143),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_145),
.B(n_194),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_213),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_142),
.A2(n_91),
.B1(n_183),
.B2(n_135),
.Y(n_258)
);

INVx3_ASAP7_75t_SL g259 ( 
.A(n_184),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_143),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_199),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_263),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_257),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_266),
.B(n_281),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_276),
.A2(n_256),
.B(n_239),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_279),
.B(n_236),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_230),
.A2(n_247),
.B1(n_204),
.B2(n_202),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_283),
.A2(n_290),
.B1(n_306),
.B2(n_307),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_251),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_228),
.B(n_221),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_286),
.B(n_265),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g287 ( 
.A(n_202),
.B(n_214),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_287),
.B(n_294),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_230),
.A2(n_247),
.B1(n_204),
.B2(n_197),
.Y(n_290)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g294 ( 
.A(n_214),
.B(n_228),
.Y(n_294)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_232),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_299),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_238),
.B(n_261),
.C(n_255),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_304),
.C(n_309),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_218),
.B(n_244),
.C(n_205),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_218),
.B(n_215),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_308),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_218),
.A2(n_233),
.B1(n_249),
.B2(n_226),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_227),
.A2(n_224),
.B1(n_225),
.B2(n_254),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_222),
.B(n_260),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_246),
.B(n_220),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_306),
.A2(n_250),
.B1(n_243),
.B2(n_259),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_312),
.A2(n_320),
.B1(n_331),
.B2(n_336),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_313),
.B(n_347),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_316),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_207),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_338),
.C(n_343),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_271),
.A2(n_243),
.B1(n_219),
.B2(n_259),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_318),
.A2(n_325),
.B1(n_341),
.B2(n_345),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_305),
.A2(n_201),
.B1(n_253),
.B2(n_203),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_321),
.A2(n_339),
.B1(n_348),
.B2(n_336),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_286),
.B(n_210),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_323),
.B(n_329),
.Y(n_367)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_324),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_271),
.A2(n_212),
.B1(n_245),
.B2(n_240),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_295),
.Y(n_328)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_328),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_262),
.B(n_264),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_330),
.B(n_335),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_304),
.A2(n_279),
.B1(n_264),
.B2(n_272),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_332),
.B(n_340),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_293),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_337),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_267),
.B(n_289),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_270),
.A2(n_276),
.B1(n_307),
.B2(n_280),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_294),
.C(n_287),
.Y(n_338)
);

AO22x1_ASAP7_75t_SL g339 ( 
.A1(n_271),
.A2(n_296),
.B1(n_309),
.B2(n_263),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_274),
.B(n_288),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_273),
.A2(n_277),
.B1(n_303),
.B2(n_310),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_266),
.B(n_273),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_342),
.B(n_344),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_284),
.B(n_277),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_303),
.A2(n_297),
.B1(n_278),
.B2(n_298),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_278),
.B(n_265),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_282),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_298),
.A2(n_275),
.B1(n_282),
.B2(n_300),
.Y(n_348)
);

NOR2x1_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_275),
.Y(n_349)
);

AO21x1_ASAP7_75t_L g396 ( 
.A1(n_349),
.A2(n_325),
.B(n_344),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_360),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_321),
.A2(n_269),
.B(n_300),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_354),
.A2(n_361),
.B(n_364),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_346),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_355),
.B(n_368),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_348),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_370),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_323),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_316),
.A2(n_269),
.B(n_302),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_326),
.A2(n_302),
.B(n_301),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_326),
.A2(n_301),
.B(n_292),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_315),
.A2(n_292),
.B1(n_311),
.B2(n_301),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_369),
.A2(n_372),
.B1(n_328),
.B2(n_324),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_329),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_315),
.A2(n_291),
.B(n_311),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_371),
.B(n_373),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_314),
.A2(n_291),
.B1(n_311),
.B2(n_337),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_345),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_320),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_314),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_333),
.Y(n_379)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_379),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_318),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_380),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_377),
.B(n_330),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_385),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_334),
.Y(n_383)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_383),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_317),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_388),
.C(n_394),
.Y(n_418)
);

BUFx12_ASAP7_75t_L g385 ( 
.A(n_371),
.Y(n_385)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_352),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_390),
.Y(n_406)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_392),
.Y(n_416)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_395),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_313),
.Y(n_394)
);

BUFx12f_ASAP7_75t_SL g395 ( 
.A(n_364),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_387),
.Y(n_410)
);

NAND5xp2_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_322),
.C(n_319),
.D(n_339),
.E(n_338),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_398),
.A2(n_339),
.B1(n_367),
.B2(n_366),
.Y(n_415)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_358),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_399),
.B(n_400),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_366),
.A2(n_333),
.B1(n_331),
.B2(n_312),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_369),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_339),
.C(n_343),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_365),
.C(n_362),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_400),
.A2(n_356),
.B1(n_375),
.B2(n_363),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_404),
.A2(n_407),
.B1(n_408),
.B2(n_419),
.Y(n_437)
);

AOI221xp5_ASAP7_75t_L g405 ( 
.A1(n_382),
.A2(n_360),
.B1(n_373),
.B2(n_363),
.C(n_342),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_381),
.A2(n_356),
.B1(n_375),
.B2(n_355),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_379),
.A2(n_357),
.B1(n_376),
.B2(n_367),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_410),
.A2(n_415),
.B(n_380),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_368),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_414),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_365),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_383),
.A2(n_377),
.B1(n_341),
.B2(n_362),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_421),
.C(n_351),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_365),
.Y(n_421)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_423),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_386),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_432),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_411),
.A2(n_397),
.B1(n_396),
.B2(n_378),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_426),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_372),
.Y(n_427)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

AOI321xp33_ASAP7_75t_L g429 ( 
.A1(n_412),
.A2(n_398),
.A3(n_378),
.B1(n_395),
.B2(n_387),
.C(n_352),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_429),
.A2(n_435),
.B(n_436),
.Y(n_443)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_416),
.Y(n_431)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_431),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_415),
.A2(n_401),
.B1(n_396),
.B2(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_433),
.Y(n_453)
);

FAx1_ASAP7_75t_L g434 ( 
.A(n_403),
.B(n_385),
.CI(n_398),
.CON(n_434),
.SN(n_434)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_434),
.A2(n_409),
.B(n_417),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_404),
.A2(n_380),
.B1(n_385),
.B2(n_391),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_417),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_412),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_411),
.A2(n_385),
.B1(n_399),
.B2(n_349),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_446),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_414),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_444),
.C(n_447),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_421),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_413),
.C(n_418),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_420),
.C(n_409),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_407),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_450),
.C(n_437),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_435),
.Y(n_450)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_448),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_455),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_452),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_443),
.A2(n_438),
.B(n_410),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_456),
.A2(n_459),
.B1(n_461),
.B2(n_422),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_458),
.B(n_450),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_445),
.A2(n_410),
.B(n_436),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_460),
.B(n_463),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_447),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_453),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_464),
.B(n_469),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_458),
.A2(n_424),
.B1(n_449),
.B2(n_441),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_462),
.A2(n_424),
.B1(n_441),
.B2(n_419),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_459),
.A2(n_430),
.B1(n_408),
.B2(n_422),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_457),
.B(n_451),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_470),
.B(n_444),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_471),
.A2(n_456),
.B(n_457),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_472),
.A2(n_473),
.B(n_465),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_467),
.A2(n_446),
.B(n_442),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_474),
.Y(n_476)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_477),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_468),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g479 ( 
.A(n_478),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_479),
.B(n_476),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_L g483 ( 
.A(n_481),
.B(n_482),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_480),
.B(n_466),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_483),
.B(n_406),
.Y(n_484)
);


endmodule