module fake_jpeg_21320_n_286 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_182;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_265;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_60),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_31),
.B1(n_23),
.B2(n_25),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_49),
.A2(n_51),
.B1(n_32),
.B2(n_21),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_31),
.B1(n_23),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_27),
.B1(n_44),
.B2(n_29),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_23),
.B1(n_35),
.B2(n_41),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_55),
.Y(n_65)
);

BUFx2_ASAP7_75t_SL g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_62),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_35),
.B1(n_27),
.B2(n_34),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_39),
.Y(n_83)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_68),
.Y(n_126)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_70),
.B(n_71),
.Y(n_128)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_83),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_50),
.B1(n_41),
.B2(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_43),
.B1(n_19),
.B2(n_36),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_43),
.B1(n_29),
.B2(n_19),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_80),
.A2(n_101),
.B1(n_103),
.B2(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_42),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_39),
.B1(n_38),
.B2(n_2),
.Y(n_129)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_26),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_30),
.B1(n_21),
.B2(n_28),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_95),
.B1(n_98),
.B2(n_20),
.Y(n_113)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_94),
.B(n_99),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_28),
.B1(n_34),
.B2(n_32),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_100),
.B(n_45),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_18),
.B1(n_20),
.B2(n_33),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_20),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_60),
.A2(n_22),
.B1(n_18),
.B2(n_33),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_46),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_46),
.A2(n_20),
.B1(n_10),
.B2(n_15),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_0),
.B(n_1),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_112),
.B(n_117),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_0),
.B(n_2),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_70),
.B1(n_68),
.B2(n_102),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_2),
.B(n_45),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_72),
.B1(n_71),
.B2(n_88),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_39),
.C(n_38),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_132),
.C(n_94),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_39),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_86),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_118),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_38),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_67),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_38),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_136),
.B(n_137),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_143),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_78),
.B1(n_97),
.B2(n_73),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_95),
.B1(n_100),
.B2(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_82),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_145),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_106),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_148),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_149),
.A2(n_155),
.B1(n_161),
.B2(n_117),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_90),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_153),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_114),
.B(n_65),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_158),
.B(n_122),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_105),
.B1(n_84),
.B2(n_87),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_104),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_160),
.B(n_162),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_69),
.C(n_80),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_129),
.C(n_120),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_121),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_93),
.B1(n_104),
.B2(n_67),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_130),
.B(n_131),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_167),
.A2(n_174),
.B(n_154),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_171),
.B1(n_116),
.B2(n_109),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_155),
.A2(n_121),
.B1(n_119),
.B2(n_111),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_173),
.B(n_115),
.Y(n_198)
);

OR2x2_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_112),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_131),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_176),
.B(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_179),
.C(n_190),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_135),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_180),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_134),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_125),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_148),
.CI(n_150),
.CON(n_196),
.SN(n_196)
);

INVxp33_ASAP7_75t_SL g187 ( 
.A(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_122),
.C(n_116),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_180),
.A2(n_162),
.B1(n_159),
.B2(n_138),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_191),
.A2(n_192),
.B(n_201),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_160),
.B(n_144),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_209),
.B(n_212),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_149),
.B1(n_141),
.B2(n_142),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_194),
.A2(n_205),
.B1(n_213),
.B2(n_171),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_210),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_157),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_161),
.B(n_136),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_207),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_163),
.B1(n_139),
.B2(n_109),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_168),
.A2(n_133),
.B1(n_2),
.B2(n_4),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_3),
.B(n_4),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_165),
.A2(n_3),
.B(n_5),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_164),
.B(n_3),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_6),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_213)
);

OAI31xp33_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_188),
.A3(n_172),
.B(n_166),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_203),
.B1(n_204),
.B2(n_175),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_179),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_227),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_177),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_228),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_184),
.C(n_190),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_165),
.C(n_183),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_172),
.Y(n_226)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_188),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_185),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_226),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_227),
.B(n_202),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_234),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_191),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_216),
.B1(n_224),
.B2(n_218),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_192),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_231),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_239),
.C(n_244),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_183),
.C(n_196),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_196),
.C(n_201),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_194),
.B1(n_195),
.B2(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_219),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_213),
.B1(n_170),
.B2(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_230),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_231),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_256),
.Y(n_265)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_255),
.Y(n_261)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_259),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_228),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_214),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_263),
.Y(n_272)
);

A2O1A1O1Ixp25_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_239),
.B(n_234),
.C(n_221),
.D(n_217),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_238),
.C(n_233),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_256),
.C(n_236),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_229),
.B(n_217),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_250),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_268),
.B(n_273),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_254),
.C(n_248),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_270),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_260),
.A2(n_245),
.B1(n_253),
.B2(n_251),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_214),
.B1(n_212),
.B2(n_250),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_209),
.A3(n_182),
.B1(n_207),
.B2(n_237),
.C1(n_265),
.C2(n_14),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_272),
.A2(n_263),
.B(n_267),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_268),
.B(n_269),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_265),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_182),
.Y(n_280)
);

NOR2x1_ASAP7_75t_SL g281 ( 
.A(n_280),
.B(n_274),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_281),
.B(n_237),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_282),
.B(n_10),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_284),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_8),
.Y(n_286)
);


endmodule