module fake_jpeg_19057_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_77),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_18),
.C(n_40),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_69),
.C(n_67),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_61),
.B1(n_68),
.B2(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_88),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_60),
.B1(n_49),
.B2(n_53),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_69),
.C(n_65),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_73),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_59),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_63),
.B1(n_52),
.B2(n_64),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_57),
.B1(n_2),
.B2(n_3),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_64),
.C(n_65),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_81),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_1),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_0),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_101),
.Y(n_110)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_104),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_116),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_115),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_82),
.B1(n_66),
.B2(n_58),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_8),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_90),
.B1(n_98),
.B2(n_55),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_2),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_120),
.B(n_109),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_122),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_SL g120 ( 
.A1(n_116),
.A2(n_4),
.A3(n_5),
.B1(n_8),
.B2(n_11),
.C1(n_13),
.C2(n_15),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_102),
.B1(n_103),
.B2(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_20),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_129),
.A2(n_131),
.B(n_123),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_131),
.B(n_128),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_118),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_136),
.A2(n_117),
.B1(n_127),
.B2(n_121),
.Y(n_137)
);

AOI21x1_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_120),
.B(n_102),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_138),
.B(n_23),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_24),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_26),
.B1(n_28),
.B2(n_32),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_33),
.B(n_34),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_39),
.Y(n_143)
);


endmodule