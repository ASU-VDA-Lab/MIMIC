module real_jpeg_5192_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_525;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_0),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_0),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_0),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_0),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_0),
.B(n_203),
.Y(n_202)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_1),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_1),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_1),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_1),
.Y(n_319)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_1),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_1),
.Y(n_348)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_2),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_2),
.Y(n_244)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_2),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_3),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_3),
.B(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_3),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_3),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_3),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_3),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_3),
.B(n_191),
.Y(n_413)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_4),
.Y(n_533)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g398 ( 
.A(n_5),
.Y(n_398)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_6),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_7),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_7),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_7),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_7),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_7),
.B(n_209),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_7),
.B(n_111),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_7),
.B(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_8),
.Y(n_213)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_8),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_8),
.Y(n_335)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_10),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_10),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_10),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_11),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_11),
.B(n_47),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_11),
.B(n_111),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_11),
.B(n_190),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_11),
.B(n_327),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_11),
.B(n_335),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_11),
.B(n_379),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_11),
.B(n_404),
.Y(n_403)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_13),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_13),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_13),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_13),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_13),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_13),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_13),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_14),
.B(n_45),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_14),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_14),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_14),
.B(n_34),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_14),
.B(n_219),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_14),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_14),
.B(n_191),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_14),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_15),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_15),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_15),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_15),
.B(n_111),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_15),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_15),
.B(n_346),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_15),
.B(n_295),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_16),
.B(n_181),
.Y(n_180)
);

NAND2x1p5_ASAP7_75t_L g271 ( 
.A(n_16),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_16),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_16),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_16),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_16),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_16),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_17),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_17),
.B(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_17),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_17),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_17),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_17),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_17),
.B(n_370),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_17),
.B(n_406),
.Y(n_405)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_19),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_19),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_19),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_19),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_19),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_19),
.B(n_267),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_527),
.B(n_530),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_43),
.B(n_81),
.C(n_526),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_24),
.B(n_48),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_41),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.C(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_26),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_26),
.A2(n_32),
.B1(n_42),
.B2(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_30),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_32),
.B(n_52),
.C(n_60),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_35),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_77),
.C(n_79),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_49),
.B(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_64),
.C(n_66),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_50),
.B(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_60),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_52),
.A2(n_59),
.B1(n_73),
.B2(n_120),
.Y(n_124)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_57),
.Y(n_209)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_57),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_67),
.C(n_73),
.Y(n_66)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_63),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_64),
.B(n_66),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_67),
.A2(n_68),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_73),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_73),
.A2(n_115),
.B1(n_116),
.B2(n_120),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_75),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_75),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_75),
.Y(n_295)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_76),
.Y(n_339)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_76),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_76),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_79),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_131),
.B(n_525),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_128),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_83),
.B(n_128),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_125),
.C(n_126),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_84),
.A2(n_85),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_113),
.C(n_121),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_86),
.A2(n_87),
.B1(n_500),
.B2(n_502),
.Y(n_499)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_99),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_93),
.C(n_99),
.Y(n_125)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.C(n_107),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_100),
.B(n_490),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_101),
.A2(n_102),
.B1(n_107),
.B2(n_108),
.Y(n_490)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_106),
.Y(n_279)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_112),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_113),
.A2(n_121),
.B1(n_122),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_113),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.C(n_120),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_114),
.B(n_496),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_115),
.A2(n_116),
.B1(n_202),
.B2(n_205),
.Y(n_201)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_116),
.B(n_199),
.C(n_202),
.Y(n_497)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_119),
.Y(n_299)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_119),
.Y(n_406)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_125),
.B(n_126),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_519),
.B(n_524),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_483),
.B(n_516),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_301),
.B(n_482),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_252),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_135),
.B(n_252),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_196),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_136),
.B(n_197),
.C(n_231),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_170),
.C(n_178),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_137),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.C(n_158),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_138),
.B(n_467),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_143),
.C(n_146),
.Y(n_177)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_147),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_148),
.A2(n_149),
.B1(n_158),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_156),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_150),
.B(n_156),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_152),
.B(n_457),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_158),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_159),
.B(n_161),
.C(n_166),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_165),
.B1(n_166),
.B2(n_169),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_161),
.Y(n_169)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_163),
.Y(n_327)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_163),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_165),
.B(n_202),
.C(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_165),
.A2(n_166),
.B1(n_202),
.B2(n_205),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_170),
.B(n_178),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_174),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_174),
.B(n_175),
.C(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_174),
.A2(n_176),
.B1(n_241),
.B2(n_245),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_176),
.B(n_236),
.C(n_245),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_192),
.C(n_194),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_179),
.B(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_189),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_180),
.B(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_184),
.B(n_189),
.Y(n_264)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_187),
.Y(n_313)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_192),
.B(n_194),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_231),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_206),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_198),
.B(n_207),
.C(n_230),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_202),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_204),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_204),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_217),
.B1(n_229),
.B2(n_230),
.Y(n_206)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_214),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_214),
.Y(n_251)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_218),
.B(n_222),
.C(n_225),
.Y(n_498)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_246),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_233),
.B(n_235),
.C(n_246),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.C(n_250),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_250),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.C(n_259),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_254),
.B(n_257),
.Y(n_477)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_259),
.B(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_280),
.C(n_283),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_261),
.B(n_470),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.C(n_269),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_262),
.A2(n_263),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_265),
.A2(n_266),
.B(n_268),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_265),
.B(n_269),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.C(n_277),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_425)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx8_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_277),
.B(n_425),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_278),
.B(n_365),
.Y(n_364)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_279),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_283),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_296),
.C(n_300),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_285),
.B(n_459),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.C(n_293),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_286),
.B(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_289),
.A2(n_293),
.B1(n_294),
.B2(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_289),
.Y(n_438)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_292),
.Y(n_365)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_296),
.B(n_300),
.Y(n_459)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI21x1_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_475),
.B(n_481),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_462),
.B(n_474),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_444),
.B(n_461),
.Y(n_303)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_418),
.B(n_443),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_388),
.B(n_417),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_357),
.B(n_387),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_341),
.B(n_356),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_321),
.B(n_340),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_317),
.B(n_320),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_315),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_323),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_331),
.B2(n_332),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_324),
.B(n_334),
.C(n_336),
.Y(n_355)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_326),
.B(n_328),
.Y(n_349)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_336),
.B2(n_337),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_355),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_355),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_350),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_349),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_349),
.C(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_347),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_350),
.Y(n_359)
);

BUFx24_ASAP7_75t_SL g534 ( 
.A(n_350),
.Y(n_534)
);

FAx1_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.CI(n_354),
.CON(n_350),
.SN(n_350)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_375),
.C(n_376),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_353),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_360),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_373),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_361),
.B(n_374),
.C(n_377),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_362),
.B(n_364),
.C(n_366),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_369),
.B2(n_372),
.Y(n_366)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_367),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_372),
.Y(n_399)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_377),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

MAJx2_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_383),
.C(n_385),
.Y(n_415)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_385),
.B2(n_386),
.Y(n_381)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_382),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_383),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_416),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_416),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_401),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_400),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_391),
.B(n_400),
.C(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_399),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_397),
.Y(n_392)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_393),
.Y(n_432)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_397),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_432),
.C(n_433),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_401),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_408),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_410),
.C(n_414),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g537 ( 
.A(n_402),
.Y(n_537)
);

FAx1_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_405),
.CI(n_407),
.CON(n_402),
.SN(n_402)
);

MAJx2_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_405),
.C(n_407),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_410),
.B1(n_414),
.B2(n_415),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_413),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_441),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_441),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_430),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_422),
.C(n_430),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_426),
.B2(n_427),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_453),
.C(n_454),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_428),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_429),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_435),
.C(n_440),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_436),
.B1(n_439),
.B2(n_440),
.Y(n_434)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_435),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_436),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_445),
.B(n_460),
.Y(n_444)
);

NOR2xp67_ASAP7_75t_SL g461 ( 
.A(n_445),
.B(n_460),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_446),
.B(n_451),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_450),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_450),
.C(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_448),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_455),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_456),
.C(n_458),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_472),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_472),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_479),
.C(n_480),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_478),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_476),
.B(n_478),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_511),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_L g516 ( 
.A1(n_484),
.A2(n_517),
.B(n_518),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_504),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_485),
.B(n_504),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_487),
.B1(n_493),
.B2(n_503),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_486),
.B(n_494),
.C(n_499),
.Y(n_523)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.C(n_491),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_488),
.B(n_507),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_489),
.A2(n_491),
.B1(n_492),
.B2(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_489),
.Y(n_508)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_493),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_499),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_497),
.C(n_498),
.Y(n_494)
);

FAx1_ASAP7_75t_SL g509 ( 
.A(n_495),
.B(n_497),
.CI(n_498),
.CON(n_509),
.SN(n_509)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_500),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_509),
.C(n_510),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_505),
.A2(n_506),
.B1(n_509),
.B2(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_509),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_509),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_513),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_512),
.B(n_515),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_515),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_520),
.B(n_523),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_523),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g521 ( 
.A(n_522),
.Y(n_521)
);

BUFx12f_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx13_ASAP7_75t_L g532 ( 
.A(n_529),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_533),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);


endmodule