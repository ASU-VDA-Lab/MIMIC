module fake_jpeg_26523_n_123 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_123);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx13_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_29),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_9),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_14),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_22),
.C(n_23),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_48),
.C(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_29),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_50),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_27),
.A2(n_19),
.B1(n_24),
.B2(n_18),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_49),
.B1(n_54),
.B2(n_15),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_22),
.C(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_19),
.B1(n_13),
.B2(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_15),
.B1(n_18),
.B2(n_21),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_0),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_46),
.C(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_38),
.Y(n_64)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_48),
.B1(n_51),
.B2(n_46),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_51),
.B1(n_52),
.B2(n_15),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_52),
.B1(n_44),
.B2(n_51),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_78),
.B1(n_56),
.B2(n_4),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_56),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_32),
.B1(n_37),
.B2(n_34),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_3),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_0),
.B(n_1),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_2),
.B(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_2),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

AO22x1_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_55),
.B1(n_70),
.B2(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_87),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_70),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_94),
.C(n_81),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_92),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_60),
.B1(n_62),
.B2(n_57),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_103),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_88),
.C(n_94),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_72),
.B(n_83),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_89),
.B(n_79),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_109),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_108),
.Y(n_112)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_104),
.C(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_111),
.Y(n_114)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_82),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_96),
.B1(n_103),
.B2(n_86),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_118),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_115),
.A3(n_112),
.B1(n_116),
.B2(n_74),
.C1(n_76),
.C2(n_77),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_76),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_77),
.B(n_5),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_121),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_119),
.Y(n_123)
);


endmodule