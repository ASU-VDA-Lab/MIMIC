module fake_aes_5128_n_23 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_23);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_23;
wire n_20;
wire n_22;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_9), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_11), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_7), .Y(n_15) );
O2A1O1Ixp5_ASAP7_75t_SL g16 ( .A1(n_14), .A2(n_0), .B(n_1), .C(n_2), .Y(n_16) );
NOR3xp33_ASAP7_75t_SL g17 ( .A(n_16), .B(n_12), .C(n_15), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_12), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_18), .B(n_13), .Y(n_19) );
AOI322xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_0), .A3(n_2), .B1(n_3), .B2(n_4), .C1(n_5), .C2(n_6), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_20), .Y(n_21) );
INVx3_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
AOI22xp5_ASAP7_75t_SL g23 ( .A1(n_22), .A2(n_3), .B1(n_8), .B2(n_10), .Y(n_23) );
endmodule