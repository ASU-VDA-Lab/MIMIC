module fake_jpeg_3630_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_7),
.B(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_30),
.B(n_0),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_2),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_7),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_1),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_78),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_1),
.B(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_4),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_3),
.B(n_4),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_65),
.B(n_61),
.C(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_3),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_86),
.B(n_98),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_59),
.B1(n_50),
.B2(n_65),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_79),
.B1(n_53),
.B2(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_54),
.Y(n_86)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_89),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_59),
.B1(n_66),
.B2(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_5),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_66),
.B1(n_69),
.B2(n_55),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_71),
.B1(n_49),
.B2(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_79),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_9),
.B(n_10),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_101),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_68),
.A3(n_55),
.B1(n_60),
.B2(n_67),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_90),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_58),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_112),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_8),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_12),
.Y(n_139)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_27),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_9),
.B(n_10),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_117),
.B(n_88),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_84),
.C(n_85),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_123),
.C(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_122),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_28),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_115),
.C(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_25),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_136),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_29),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_24),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_11),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_31),
.C(n_44),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_35),
.Y(n_154)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_144),
.C(n_147),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_15),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_16),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_16),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_17),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_149),
.B(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_124),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_156),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_33),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_138),
.C(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_17),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_158),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_169),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_134),
.B(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_166),
.B(n_170),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_152),
.C(n_153),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_146),
.B1(n_145),
.B2(n_140),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_20),
.B1(n_21),
.B2(n_32),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_173),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_153),
.C(n_155),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_154),
.C(n_148),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_161),
.B(n_165),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_176),
.A2(n_166),
.B(n_174),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_178),
.B(n_180),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_165),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_184),
.B(n_171),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_168),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_183),
.A3(n_162),
.B1(n_169),
.B2(n_170),
.C1(n_167),
.C2(n_39),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_38),
.C(n_41),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_47),
.Y(n_188)
);


endmodule