module fake_jpeg_3799_n_157 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_157);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_27),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_52),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_17),
.B1(n_22),
.B2(n_26),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_51),
.B1(n_58),
.B2(n_11),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_18),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_67),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_22),
.B1(n_28),
.B2(n_26),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_55),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_24),
.C(n_30),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_13),
.C(n_48),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_31),
.A2(n_28),
.B1(n_20),
.B2(n_27),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_70),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_69),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_23),
.B1(n_19),
.B2(n_16),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_66),
.B1(n_71),
.B2(n_8),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_20),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_73),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_32),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_33),
.B(n_27),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_31),
.A2(n_20),
.B1(n_27),
.B2(n_10),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_4),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_3),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_4),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_8),
.Y(n_87)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_7),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_88),
.Y(n_109)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_86),
.Y(n_101)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_9),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_94),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_92),
.B1(n_53),
.B2(n_45),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_63),
.B1(n_51),
.B2(n_66),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_59),
.B(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_50),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_70),
.B(n_59),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_88),
.B(n_82),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_55),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_105),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_68),
.C(n_67),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_107),
.C(n_115),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_71),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_83),
.B(n_81),
.Y(n_125)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_97),
.B1(n_95),
.B2(n_90),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_91),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_97),
.B1(n_84),
.B2(n_86),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_125),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_120),
.B(n_113),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_96),
.B(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_87),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_83),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_98),
.B1(n_115),
.B2(n_108),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_107),
.C(n_102),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_134),
.C(n_138),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_102),
.C(n_109),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_85),
.B1(n_111),
.B2(n_108),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_124),
.B(n_121),
.C(n_129),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_116),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_137),
.A2(n_118),
.B(n_132),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_103),
.C(n_93),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_141),
.A2(n_146),
.B1(n_130),
.B2(n_132),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_123),
.C(n_127),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_144),
.C(n_134),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_128),
.C(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_121),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_152),
.A2(n_133),
.B(n_148),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_149),
.B(n_142),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_154),
.B(n_121),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_99),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_117),
.Y(n_157)
);


endmodule