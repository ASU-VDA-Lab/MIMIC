module fake_jpeg_2976_n_502 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_502);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_502;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_55),
.Y(n_105)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_52),
.Y(n_154)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_53),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_54),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_27),
.B(n_0),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_57),
.Y(n_157)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_58),
.Y(n_159)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_1),
.B(n_2),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_97),
.C(n_69),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_65),
.Y(n_133)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_82),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_78),
.Y(n_113)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_81),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_19),
.B(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_97),
.Y(n_108)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_95),
.Y(n_146)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_91),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_90),
.B(n_71),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_48),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_25),
.B(n_2),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_48),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_66),
.B1(n_92),
.B2(n_52),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_100),
.A2(n_114),
.B1(n_147),
.B2(n_93),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_111),
.B(n_138),
.C(n_63),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_59),
.A2(n_48),
.B1(n_42),
.B2(n_40),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_112),
.A2(n_126),
.B1(n_149),
.B2(n_153),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_68),
.A2(n_30),
.B1(n_42),
.B2(n_40),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_61),
.A2(n_30),
.B1(n_42),
.B2(n_40),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_115),
.A2(n_131),
.B1(n_36),
.B2(n_29),
.Y(n_175)
);

OR2x2_ASAP7_75t_SL g190 ( 
.A(n_122),
.B(n_70),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_156),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_67),
.A2(n_30),
.B1(n_42),
.B2(n_40),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g200 ( 
.A(n_127),
.Y(n_200)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_53),
.B(n_34),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_129),
.B(n_130),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_57),
.B(n_35),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_48),
.B1(n_25),
.B2(n_26),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_72),
.B(n_34),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_136),
.B(n_137),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_73),
.B(n_46),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_19),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_79),
.B(n_44),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_140),
.B(n_2),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_77),
.A2(n_33),
.B1(n_26),
.B2(n_39),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_62),
.A2(n_33),
.B1(n_26),
.B2(n_39),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_74),
.A2(n_33),
.B1(n_26),
.B2(n_39),
.Y(n_153)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_51),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_87),
.B(n_35),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_54),
.Y(n_158)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_54),
.B(n_39),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_85),
.Y(n_163)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_163),
.B(n_190),
.Y(n_247)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_164),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_160),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_165),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_108),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_166),
.B(n_177),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_168),
.B(n_199),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_112),
.A2(n_33),
.B1(n_36),
.B2(n_21),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_169),
.A2(n_175),
.B1(n_178),
.B2(n_196),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_115),
.A2(n_36),
.B1(n_21),
.B2(n_43),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_170),
.A2(n_176),
.B(n_165),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_117),
.B(n_94),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_120),
.C(n_104),
.Y(n_222)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_94),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_174),
.B(n_204),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_131),
.A2(n_36),
.B1(n_29),
.B2(n_43),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_44),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_114),
.A2(n_31),
.B1(n_75),
.B2(n_63),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_31),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_75),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_183),
.Y(n_253)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_185),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_186),
.A2(n_206),
.B1(n_217),
.B2(n_218),
.Y(n_237)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_189),
.Y(n_272)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_195),
.Y(n_241)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_147),
.A2(n_100),
.B1(n_103),
.B2(n_101),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_102),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_214),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_116),
.B(n_96),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_201),
.B(n_202),
.Y(n_265)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_116),
.B(n_3),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_143),
.B(n_3),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_205),
.B(n_210),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_127),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_121),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_207),
.B(n_209),
.Y(n_250)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_208),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_121),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_148),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_148),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_211),
.Y(n_255)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_141),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_219),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_104),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_128),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_141),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_247),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_175),
.A2(n_106),
.B1(n_110),
.B2(n_135),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_224),
.A2(n_227),
.B1(n_230),
.B2(n_235),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_119),
.C(n_120),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_225),
.B(n_236),
.C(n_256),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_170),
.A2(n_106),
.B1(n_110),
.B2(n_135),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_176),
.A2(n_151),
.B1(n_119),
.B2(n_124),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_165),
.A2(n_124),
.B(n_123),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_231),
.A2(n_270),
.B(n_179),
.Y(n_306)
);

AOI32xp33_ASAP7_75t_L g232 ( 
.A1(n_181),
.A2(n_139),
.A3(n_158),
.B1(n_150),
.B2(n_9),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_232),
.B(n_233),
.Y(n_288)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_167),
.A2(n_139),
.A3(n_150),
.B1(n_8),
.B2(n_9),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_166),
.B(n_7),
.C(n_9),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_245),
.A2(n_264),
.B1(n_237),
.B2(n_255),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_248),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_10),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_163),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_257),
.A2(n_259),
.B1(n_210),
.B2(n_161),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_177),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_163),
.A2(n_14),
.B(n_15),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_261),
.A2(n_264),
.B(n_267),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_180),
.A2(n_14),
.B(n_16),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_SL g266 ( 
.A(n_171),
.B(n_16),
.C(n_17),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_206),
.C(n_186),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_199),
.A2(n_172),
.B(n_178),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_182),
.B(n_187),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_268),
.B(n_269),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_171),
.A2(n_169),
.B(n_198),
.C(n_189),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_186),
.A2(n_219),
.B(n_216),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_273),
.B(n_223),
.Y(n_340)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_275),
.Y(n_344)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_276),
.Y(n_345)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_277),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_246),
.A2(n_186),
.B1(n_218),
.B2(n_200),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_278),
.A2(n_319),
.B1(n_257),
.B2(n_266),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_173),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_292),
.Y(n_323)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_280),
.Y(n_328)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_282),
.Y(n_357)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_283),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_223),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_284),
.B(n_285),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_265),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_214),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_287),
.B(n_298),
.C(n_304),
.Y(n_322)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_290),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_240),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_294),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_226),
.B(n_201),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_226),
.B(n_194),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_301),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_228),
.B(n_202),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_296),
.B(n_297),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_268),
.B(n_208),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_238),
.B(n_193),
.C(n_191),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_299),
.A2(n_307),
.B1(n_313),
.B2(n_314),
.Y(n_335)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_221),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_300),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_203),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_228),
.B(n_197),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_303),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_249),
.B(n_183),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_247),
.B(n_188),
.C(n_164),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_247),
.B(n_179),
.C(n_200),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_305),
.B(n_316),
.C(n_271),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_306),
.A2(n_242),
.B(n_254),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_246),
.A2(n_184),
.B1(n_185),
.B2(n_162),
.Y(n_307)
);

AND2x6_ASAP7_75t_L g308 ( 
.A(n_225),
.B(n_162),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_308),
.B(n_310),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_249),
.B(n_184),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_309),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_236),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_221),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_315),
.Y(n_355)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_267),
.A2(n_224),
.B1(n_227),
.B2(n_269),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_245),
.A2(n_230),
.B1(n_248),
.B2(n_270),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_221),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_222),
.B(n_256),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_244),
.B(n_239),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g358 ( 
.A(n_317),
.Y(n_358)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_301),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_320),
.B(n_311),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g321 ( 
.A1(n_306),
.A2(n_231),
.B(n_250),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_321),
.B(n_305),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_314),
.A2(n_241),
.B1(n_232),
.B2(n_233),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_338),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_287),
.B(n_244),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_326),
.B(n_329),
.C(n_337),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_339),
.B1(n_356),
.B2(n_295),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_261),
.C(n_235),
.Y(n_329)
);

BUFx16f_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

BUFx24_ASAP7_75t_L g359 ( 
.A(n_330),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_286),
.A2(n_255),
.B(n_258),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_331),
.A2(n_351),
.B(n_298),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_315),
.B(n_300),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_273),
.B(n_243),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_288),
.A2(n_229),
.B1(n_262),
.B2(n_240),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_278),
.A2(n_262),
.B1(n_263),
.B2(n_223),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_340),
.B(n_354),
.C(n_322),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_277),
.A2(n_263),
.B1(n_258),
.B2(n_271),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_282),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_286),
.A2(n_242),
.B(n_253),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_280),
.A2(n_253),
.B1(n_271),
.B2(n_313),
.Y(n_356)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_333),
.Y(n_360)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_327),
.A2(n_295),
.B1(n_307),
.B2(n_274),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_362),
.A2(n_376),
.B1(n_349),
.B2(n_353),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_363),
.B(n_375),
.Y(n_393)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_357),
.Y(n_364)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_364),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_310),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_380),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_366),
.A2(n_372),
.B(n_373),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_335),
.A2(n_328),
.B1(n_325),
.B2(n_356),
.Y(n_367)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_357),
.Y(n_368)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_369),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_382),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_325),
.A2(n_275),
.B1(n_276),
.B2(n_294),
.Y(n_371)
);

OAI22x1_ASAP7_75t_L g392 ( 
.A1(n_371),
.A2(n_321),
.B1(n_332),
.B2(n_323),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_355),
.A2(n_281),
.B(n_279),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_328),
.A2(n_293),
.B1(n_292),
.B2(n_308),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_377),
.A2(n_351),
.B(n_338),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_354),
.C(n_322),
.Y(n_397)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_334),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_346),
.A2(n_299),
.B(n_283),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_385),
.Y(n_410)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_336),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_326),
.B(n_289),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_330),
.Y(n_408)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_336),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_384),
.B(n_386),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_324),
.A2(n_281),
.B1(n_304),
.B2(n_289),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_346),
.A2(n_290),
.B1(n_318),
.B2(n_347),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_339),
.A2(n_352),
.B1(n_321),
.B2(n_355),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_387),
.Y(n_416)
);

NOR3xp33_ASAP7_75t_SL g388 ( 
.A(n_358),
.B(n_342),
.C(n_343),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_389),
.Y(n_405)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_390),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_330),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_391),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_392),
.A2(n_381),
.B1(n_362),
.B2(n_361),
.Y(n_433)
);

OA22x2_ASAP7_75t_L g396 ( 
.A1(n_389),
.A2(n_343),
.B1(n_331),
.B2(n_353),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_401),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_397),
.B(n_398),
.C(n_399),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_340),
.C(n_337),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_329),
.C(n_323),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_373),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_411),
.C(n_377),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_350),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_409),
.B(n_413),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_374),
.B(n_350),
.C(n_385),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_376),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_384),
.Y(n_421)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_421),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_403),
.B(n_382),
.Y(n_422)
);

OAI321xp33_ASAP7_75t_L g460 ( 
.A1(n_422),
.A2(n_424),
.A3(n_431),
.B1(n_360),
.B2(n_391),
.C(n_388),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_417),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_394),
.B(n_369),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_418),
.Y(n_425)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_425),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_418),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_426),
.A2(n_436),
.B1(n_439),
.B2(n_440),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_392),
.A2(n_366),
.B(n_377),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_427),
.A2(n_428),
.B(n_415),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_415),
.A2(n_400),
.B(n_410),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_414),
.B(n_375),
.Y(n_430)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_430),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_405),
.B(n_379),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_399),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_433),
.A2(n_434),
.B1(n_406),
.B2(n_417),
.Y(n_456)
);

AOI221xp5_ASAP7_75t_L g434 ( 
.A1(n_416),
.A2(n_361),
.B1(n_381),
.B2(n_368),
.C(n_364),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_395),
.B(n_390),
.Y(n_435)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_435),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_396),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_398),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_397),
.Y(n_448)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_438),
.Y(n_452)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_404),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_396),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_396),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_433),
.A2(n_401),
.B1(n_393),
.B2(n_407),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_442),
.A2(n_456),
.B1(n_460),
.B2(n_441),
.Y(n_462)
);

AOI221xp5_ASAP7_75t_L g443 ( 
.A1(n_422),
.A2(n_407),
.B1(n_410),
.B2(n_412),
.C(n_393),
.Y(n_443)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_443),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_431),
.B(n_409),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_451),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_455),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_449),
.A2(n_450),
.B(n_453),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_393),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_427),
.A2(n_410),
.B(n_413),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_420),
.B(n_411),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_429),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_430),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_462),
.A2(n_469),
.B1(n_446),
.B2(n_457),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_445),
.A2(n_419),
.B1(n_436),
.B2(n_421),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_464),
.A2(n_468),
.B1(n_450),
.B2(n_458),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_424),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_466),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_445),
.A2(n_419),
.B1(n_428),
.B2(n_434),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_442),
.A2(n_425),
.B1(n_423),
.B2(n_435),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_437),
.C(n_420),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_471),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_432),
.C(n_429),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_449),
.A2(n_429),
.B(n_439),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_472),
.A2(n_458),
.B(n_459),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_474),
.B(n_446),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_453),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_478),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g477 ( 
.A(n_467),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_479),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_461),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_481),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_483),
.A2(n_468),
.B1(n_464),
.B2(n_452),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_451),
.C(n_440),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_484),
.B(n_466),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_482),
.A2(n_472),
.B(n_463),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_485),
.B(n_490),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_489),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_476),
.A2(n_463),
.B(n_469),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_491),
.B(n_475),
.C(n_483),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_493),
.A2(n_494),
.B(n_486),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_484),
.Y(n_494)
);

AOI31xp33_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_497),
.A3(n_471),
.B(n_492),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_495),
.A2(n_488),
.B(n_461),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_498),
.A2(n_492),
.B(n_488),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_499),
.A2(n_491),
.B(n_452),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_500),
.A2(n_359),
.B1(n_438),
.B2(n_495),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_359),
.B(n_495),
.Y(n_502)
);


endmodule