module real_jpeg_12745_n_17 (n_5, n_4, n_8, n_0, n_12, n_250, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_250;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_1),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_184)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_4),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_5),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_81)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_58),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_58),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_58),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_60),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_60),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_60),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_44),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_10),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_69),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_69),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_69),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_14),
.B(n_54),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_139),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_14),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_14),
.B(n_26),
.C(n_40),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_14),
.B(n_63),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_14),
.A2(n_99),
.B(n_155),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_14),
.A2(n_49),
.B(n_64),
.C(n_182),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_139),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_14),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_15),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_15),
.B(n_50),
.Y(n_126)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_20),
.B(n_104),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_46),
.C(n_61),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_22),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_23),
.B(n_33),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_24),
.A2(n_28),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_24),
.A2(n_28),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_24),
.B(n_156),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_25),
.A2(n_26),
.B1(n_40),
.B2(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_25),
.B(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_28),
.B(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_31),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B1(n_43),
.B2(n_45),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_37),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_36),
.B(n_144),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_37),
.A2(n_65),
.B(n_139),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_38),
.A2(n_45),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_38),
.A2(n_43),
.B1(n_45),
.B2(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_38),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_38),
.B(n_142),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_38),
.A2(n_45),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_42),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_42),
.B(n_139),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_42),
.A2(n_152),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_45),
.B(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_46),
.B(n_61),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_57),
.B2(n_59),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_47),
.A2(n_59),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_47),
.A2(n_55),
.B(n_139),
.C(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_48),
.A2(n_57),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_48),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_71)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_49),
.A2(n_52),
.A3(n_55),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_66),
.B(n_67),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_66),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_62),
.A2(n_67),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_62),
.A2(n_90),
.B1(n_117),
.B2(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2x1_ASAP7_75t_R g70 ( 
.A(n_63),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_68),
.Y(n_118)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_85),
.B2(n_86),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_84),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_80),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_96),
.B2(n_103),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_90),
.A2(n_118),
.B(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_94),
.B(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_100),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_99),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_99),
.A2(n_100),
.B1(n_121),
.B2(n_184),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_100),
.A2(n_161),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_100),
.B(n_139),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_100),
.A2(n_169),
.B(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.C(n_109),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_105),
.B(n_107),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_109),
.B(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.C(n_119),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_110),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_237)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_119),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_120),
.A2(n_123),
.B1(n_124),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_120),
.Y(n_231)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_125),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI321xp33_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_233),
.A3(n_242),
.B1(n_247),
.B2(n_248),
.C(n_250),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_215),
.B(n_232),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_194),
.B(n_214),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_177),
.B(n_193),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_157),
.B(n_176),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_145),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_135),
.B(n_145),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_143),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_137),
.B1(n_143),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_140),
.B(n_141),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_140),
.A2(n_141),
.B(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_153),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_150),
.C(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_154),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_165),
.B(n_175),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_163),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_170),
.B(n_174),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_178),
.B(n_179),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_188),
.C(n_192),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_183),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_196),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_207),
.B2(n_208),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_210),
.C(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_202),
.C(n_206),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_217),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_228),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_229),
.C(n_230),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_227),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_224),
.C(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_240),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_240),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.C(n_239),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_235),
.A2(n_236),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_238),
.B(n_239),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);


endmodule