module fake_jpeg_30463_n_474 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_474);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_474;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_1),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_50),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_53),
.B(n_56),
.Y(n_122)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_61),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_63),
.B(n_65),
.Y(n_140)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_1),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_73),
.B(n_78),
.Y(n_147)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_18),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_89),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_82),
.B(n_85),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_27),
.Y(n_85)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_18),
.B(n_3),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_98),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_30),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_42),
.B1(n_37),
.B2(n_27),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_106),
.A2(n_130),
.B1(n_131),
.B2(n_139),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_42),
.B1(n_37),
.B2(n_27),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_114),
.A2(n_136),
.B1(n_144),
.B2(n_156),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_60),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_53),
.A2(n_49),
.B1(n_29),
.B2(n_25),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_30),
.B1(n_27),
.B2(n_37),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_20),
.B1(n_32),
.B2(n_41),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_134),
.A2(n_19),
.B1(n_45),
.B2(n_31),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_58),
.A2(n_42),
.B1(n_20),
.B2(n_41),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_63),
.B(n_34),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_50),
.A2(n_34),
.B1(n_29),
.B2(n_25),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_63),
.B(n_24),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_67),
.A2(n_41),
.B1(n_39),
.B2(n_38),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_52),
.B(n_24),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_55),
.B(n_45),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_75),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_124),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_95),
.A2(n_33),
.B1(n_39),
.B2(n_38),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_192),
.Y(n_216)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_62),
.B1(n_96),
.B2(n_94),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_162),
.A2(n_191),
.B1(n_203),
.B2(n_156),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_100),
.A2(n_51),
.B1(n_93),
.B2(n_84),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_163),
.A2(n_175),
.B1(n_188),
.B2(n_4),
.Y(n_237)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_19),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_165),
.B(n_167),
.Y(n_223)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_155),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_170),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_174),
.Y(n_235)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_107),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_178),
.B(n_179),
.Y(n_229)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_134),
.B(n_86),
.CI(n_95),
.CON(n_180),
.SN(n_180)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_180),
.B(n_200),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_181),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_33),
.B(n_39),
.C(n_38),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_L g241 ( 
.A1(n_182),
.A2(n_186),
.B(n_190),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_101),
.B(n_56),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_97),
.B1(n_69),
.B2(n_31),
.Y(n_185)
);

AO22x1_ASAP7_75t_SL g206 ( 
.A1(n_185),
.A2(n_114),
.B1(n_109),
.B2(n_137),
.Y(n_206)
);

OR2x2_ASAP7_75t_SL g186 ( 
.A(n_103),
.B(n_83),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_187),
.A2(n_197),
.B1(n_117),
.B2(n_6),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_70),
.B1(n_79),
.B2(n_76),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g224 ( 
.A(n_189),
.B(n_195),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_56),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_131),
.A2(n_33),
.B1(n_20),
.B2(n_35),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_117),
.B(n_72),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_194),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_117),
.B(n_35),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_143),
.A2(n_80),
.B1(n_35),
.B2(n_32),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_137),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_108),
.B(n_32),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_133),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_110),
.B(n_66),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_186),
.C(n_180),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_118),
.A2(n_31),
.B1(n_43),
.B2(n_17),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_121),
.B(n_3),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_121),
.B1(n_43),
.B2(n_143),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_208),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_206),
.A2(n_226),
.B(n_227),
.C(n_231),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_196),
.A2(n_154),
.B1(n_151),
.B2(n_113),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_210),
.A2(n_212),
.B1(n_217),
.B2(n_237),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_196),
.A2(n_151),
.B1(n_113),
.B2(n_116),
.Y(n_212)
);

XOR2x2_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_120),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_SL g244 ( 
.A(n_213),
.B(n_159),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_169),
.A2(n_116),
.B1(n_102),
.B2(n_148),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_202),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_169),
.A2(n_141),
.B1(n_118),
.B2(n_102),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_168),
.A2(n_141),
.B1(n_109),
.B2(n_120),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_168),
.B(n_115),
.C(n_127),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_228),
.B(n_205),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_159),
.A2(n_132),
.B1(n_115),
.B2(n_43),
.Y(n_231)
);

BUFx4f_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_161),
.A2(n_15),
.B1(n_6),
.B2(n_8),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_240),
.A2(n_191),
.B1(n_200),
.B2(n_179),
.Y(n_245)
);

AO22x1_ASAP7_75t_L g294 ( 
.A1(n_244),
.A2(n_206),
.B1(n_224),
.B2(n_217),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_245),
.A2(n_246),
.B1(n_259),
.B2(n_208),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_237),
.A2(n_185),
.B1(n_202),
.B2(n_180),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_167),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_247),
.B(n_256),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_175),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_254),
.Y(n_281)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_209),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_251),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_185),
.B1(n_188),
.B2(n_160),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_252),
.A2(n_265),
.B1(n_219),
.B2(n_215),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_204),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_223),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_241),
.A2(n_185),
.B(n_182),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_257),
.A2(n_218),
.B(n_231),
.Y(n_289)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_263),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_240),
.C(n_226),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_165),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_268),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_227),
.A2(n_176),
.B1(n_197),
.B2(n_187),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_192),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g269 ( 
.A1(n_213),
.A2(n_201),
.A3(n_164),
.B1(n_172),
.B2(n_166),
.Y(n_269)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_242),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_270),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_214),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_170),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_277),
.A2(n_303),
.B1(n_255),
.B2(n_243),
.Y(n_331)
);

NOR4xp25_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_213),
.C(n_221),
.D(n_228),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_278),
.B(n_289),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_283),
.A2(n_287),
.B1(n_296),
.B2(n_267),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_210),
.B1(n_212),
.B2(n_206),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_248),
.A2(n_267),
.B1(n_250),
.B2(n_259),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_301),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_269),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_270),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_295),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_255),
.A2(n_206),
.B1(n_236),
.B2(n_239),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_300),
.C(n_245),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_257),
.A2(n_234),
.B(n_224),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_302),
.B(n_253),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_251),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_299),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_234),
.C(n_211),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_267),
.A2(n_239),
.B1(n_236),
.B2(n_211),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_230),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_255),
.A2(n_207),
.B1(n_230),
.B2(n_195),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_267),
.A2(n_157),
.B1(n_177),
.B2(n_189),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_207),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_308),
.B(n_315),
.Y(n_342)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_256),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_312),
.B(n_318),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_313),
.A2(n_315),
.B(n_334),
.Y(n_345)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_294),
.A2(n_253),
.B(n_244),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_316),
.Y(n_346)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_317),
.B(n_322),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_264),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_319),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_320),
.B(n_324),
.C(n_289),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_287),
.A2(n_267),
.B1(n_268),
.B2(n_243),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_321),
.A2(n_328),
.B1(n_301),
.B2(n_306),
.Y(n_347)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_275),
.C(n_274),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_325),
.A2(n_329),
.B1(n_331),
.B2(n_335),
.Y(n_362)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_330),
.Y(n_340)
);

BUFx2_ASAP7_75t_SL g333 ( 
.A(n_276),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_333),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_294),
.A2(n_255),
.B(n_272),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_307),
.B(n_266),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_336),
.A2(n_295),
.B(n_276),
.Y(n_354)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_337),
.A2(n_280),
.B(n_258),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_332),
.A2(n_283),
.B1(n_304),
.B2(n_297),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_339),
.A2(n_344),
.B1(n_364),
.B2(n_334),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_349),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_332),
.A2(n_304),
.B1(n_291),
.B2(n_298),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_347),
.A2(n_335),
.B1(n_357),
.B2(n_364),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_350),
.C(n_351),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_281),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_281),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_282),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_308),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_359),
.C(n_361),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_323),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_321),
.B(n_278),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_SL g390 ( 
.A(n_356),
.B(n_319),
.Y(n_390)
);

XOR2x2_ASAP7_75t_SL g357 ( 
.A(n_312),
.B(n_282),
.Y(n_357)
);

OAI21xp33_ASAP7_75t_L g376 ( 
.A1(n_357),
.A2(n_327),
.B(n_309),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_325),
.B(n_302),
.C(n_307),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_302),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_331),
.A2(n_277),
.B1(n_290),
.B2(n_299),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_354),
.Y(n_366)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_377),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_323),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_368),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_336),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_371),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_365),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_381),
.Y(n_407)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_346),
.Y(n_374)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_374),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_376),
.B(n_319),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_362),
.A2(n_327),
.B1(n_310),
.B2(n_316),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_365),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_382),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_351),
.B(n_285),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_383),
.B(n_385),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_359),
.B(n_311),
.Y(n_384)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_386),
.C(n_387),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_322),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_350),
.B(n_317),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_344),
.B(n_314),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_360),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_388),
.A2(n_363),
.B(n_346),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_348),
.B(n_337),
.C(n_280),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_389),
.B(n_349),
.C(n_342),
.Y(n_391)
);

MAJx2_ASAP7_75t_L g392 ( 
.A(n_390),
.B(n_353),
.C(n_345),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_400),
.C(n_403),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_406),
.Y(n_424)
);

XOR2x2_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_352),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_375),
.Y(n_414)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_395),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_379),
.A2(n_345),
.B(n_356),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_396),
.A2(n_398),
.B(n_378),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_379),
.A2(n_367),
.B(n_366),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_339),
.C(n_347),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_338),
.C(n_340),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_411),
.B(n_414),
.Y(n_436)
);

BUFx24_ASAP7_75t_SL g412 ( 
.A(n_408),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_412),
.B(n_407),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_373),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_413),
.B(n_415),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_399),
.A2(n_390),
.B(n_371),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_401),
.A2(n_377),
.B1(n_380),
.B2(n_369),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_417),
.A2(n_393),
.B1(n_404),
.B2(n_260),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_380),
.C(n_374),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_419),
.C(n_396),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_388),
.C(n_383),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_399),
.A2(n_382),
.B(n_330),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_395),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_397),
.B(n_290),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_421),
.B(n_422),
.Y(n_439)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_405),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_286),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_406),
.Y(n_426)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_425),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_427),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_430),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_391),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_437),
.C(n_158),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_410),
.A2(n_401),
.B1(n_402),
.B2(n_409),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_418),
.B(n_416),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_434),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_416),
.B(n_392),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_415),
.A2(n_402),
.B1(n_404),
.B2(n_398),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_435),
.B(n_438),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_431),
.A2(n_424),
.B(n_420),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_442),
.A2(n_15),
.B(n_6),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_437),
.B(n_419),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_444),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_432),
.A2(n_424),
.B1(n_417),
.B2(n_249),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_434),
.B(n_235),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_447),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_439),
.B(n_235),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_436),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_449),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_427),
.A2(n_233),
.B1(n_174),
.B2(n_173),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_10),
.Y(n_460)
);

NOR2x1_ASAP7_75t_L g452 ( 
.A(n_444),
.B(n_436),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_452),
.A2(n_440),
.B(n_442),
.C(n_441),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_451),
.B(n_429),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_453),
.A2(n_455),
.B(n_457),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_445),
.A2(n_5),
.B(n_6),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_448),
.B(n_8),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_10),
.B(n_11),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_11),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_462),
.B(n_465),
.C(n_452),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_463),
.B(n_464),
.Y(n_469)
);

A2O1A1O1Ixp25_ASAP7_75t_L g464 ( 
.A1(n_456),
.A2(n_450),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_459),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_466),
.A2(n_454),
.B(n_460),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_468),
.Y(n_471)
);

OAI321xp33_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_461),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_470),
.B(n_11),
.C(n_12),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_472),
.A2(n_471),
.B(n_13),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_473),
.B(n_14),
.Y(n_474)
);


endmodule