module fake_netlist_5_955_n_36 (n_8, n_10, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_11, n_6, n_1, n_36);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_11;
input n_6;
input n_1;

output n_36;

wire n_29;
wire n_16;
wire n_12;
wire n_25;
wire n_18;
wire n_27;
wire n_22;
wire n_24;
wire n_28;
wire n_21;
wire n_34;
wire n_32;
wire n_35;
wire n_17;
wire n_19;
wire n_15;
wire n_26;
wire n_30;
wire n_33;
wire n_14;
wire n_31;
wire n_23;
wire n_13;
wire n_20;

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_6),
.B(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx8_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2x1p5_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_1),
.Y(n_20)
);

OA21x2_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_0),
.B(n_2),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_20),
.A2(n_18),
.B1(n_12),
.B2(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_18),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_16),
.A2(n_12),
.B(n_17),
.Y(n_24)
);

NOR2x1_ASAP7_75t_SL g25 ( 
.A(n_15),
.B(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_17),
.B1(n_21),
.B2(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_21),
.B(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_32),
.Y(n_33)
);

OAI211xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_29),
.B(n_28),
.C(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_34),
.B(n_30),
.Y(n_36)
);


endmodule