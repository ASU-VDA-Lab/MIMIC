module fake_jpeg_5840_n_101 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_64),
.Y(n_67)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_49),
.B1(n_39),
.B2(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_70),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_54),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_50),
.B1(n_57),
.B2(n_51),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_49),
.B(n_43),
.C(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_75),
.B(n_76),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_0),
.C(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_41),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_65),
.C(n_55),
.Y(n_82)
);

FAx1_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_58),
.CI(n_44),
.CON(n_85),
.SN(n_85)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_20),
.B1(n_2),
.B2(n_4),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_84),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_77),
.B(n_83),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

AO221x1_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.C(n_13),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_9),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_91),
.B1(n_11),
.B2(n_16),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_10),
.B1(n_17),
.B2(n_18),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_19),
.C(n_22),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_23),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_24),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_26),
.Y(n_101)
);


endmodule