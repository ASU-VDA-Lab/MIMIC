module fake_jpeg_7033_n_99 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_0),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.Y(n_67)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_43),
.B1(n_51),
.B2(n_47),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_52),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_53),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_57),
.B1(n_46),
.B2(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_58),
.B1(n_55),
.B2(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_76),
.B(n_1),
.Y(n_79)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_79),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_75),
.A2(n_68),
.B1(n_71),
.B2(n_59),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_82),
.B1(n_84),
.B2(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_2),
.B1(n_4),
.B2(n_8),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_81),
.A2(n_54),
.B(n_48),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_10),
.B(n_11),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_12),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_14),
.B(n_15),
.C(n_17),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_20),
.Y(n_96)
);

AOI322xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_21),
.A3(n_23),
.B1(n_27),
.B2(n_29),
.C1(n_31),
.C2(n_32),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_35),
.B(n_37),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_39),
.C(n_40),
.Y(n_99)
);


endmodule