module real_aes_8948_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_884;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_316;
wire n_532;
wire n_746;
wire n_656;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_754;
wire n_607;
wire n_449;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_0), .A2(n_190), .B1(n_466), .B2(n_468), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_1), .A2(n_87), .B1(n_535), .B2(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_2), .A2(n_51), .B1(n_520), .B2(n_521), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_3), .A2(n_272), .B1(n_362), .B2(n_451), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_4), .A2(n_844), .B1(n_866), .B2(n_867), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_4), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_5), .A2(n_255), .B1(n_451), .B2(n_646), .Y(n_890) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_6), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g761 ( .A1(n_7), .A2(n_279), .B1(n_604), .B2(n_605), .Y(n_761) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_8), .A2(n_33), .B1(n_135), .B2(n_329), .C1(n_442), .C2(n_443), .Y(n_441) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_9), .A2(n_112), .B1(n_489), .B2(n_575), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_10), .A2(n_91), .B1(n_365), .B2(n_390), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_11), .A2(n_138), .B1(n_520), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_12), .A2(n_269), .B1(n_509), .B2(n_731), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_13), .A2(n_114), .B1(n_509), .B2(n_510), .Y(n_856) );
AOI22xp33_ASAP7_75t_SL g864 ( .A1(n_14), .A2(n_241), .B1(n_516), .B2(n_815), .Y(n_864) );
INVx1_ASAP7_75t_L g849 ( .A(n_15), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_16), .A2(n_126), .B1(n_466), .B2(n_505), .Y(n_887) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_17), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_18), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_19), .A2(n_236), .B1(n_535), .B2(n_537), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_20), .A2(n_143), .B1(n_730), .B2(n_731), .C(n_732), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_21), .A2(n_43), .B1(n_521), .B2(n_568), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_22), .A2(n_159), .B1(n_505), .B2(n_851), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_23), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_24), .A2(n_165), .B1(n_472), .B2(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_25), .A2(n_149), .B1(n_444), .B2(n_617), .Y(n_807) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_26), .A2(n_49), .B1(n_426), .B2(n_430), .C(n_432), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_27), .A2(n_234), .B1(n_401), .B2(n_404), .C(n_405), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_28), .A2(n_146), .B1(n_362), .B2(n_365), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_29), .A2(n_278), .B1(n_528), .B2(n_529), .Y(n_527) );
AO22x2_ASAP7_75t_L g311 ( .A1(n_30), .A2(n_102), .B1(n_312), .B2(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g840 ( .A(n_30), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_31), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_32), .A2(n_56), .B1(n_770), .B2(n_771), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_34), .A2(n_253), .B1(n_520), .B2(n_521), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_35), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_36), .A2(n_89), .B1(n_380), .B2(n_413), .C(n_417), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_37), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_38), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_39), .A2(n_225), .B1(n_860), .B2(n_861), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_40), .A2(n_247), .B1(n_390), .B2(n_646), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_41), .A2(n_274), .B1(n_575), .B2(n_669), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_42), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_44), .A2(n_151), .B1(n_607), .B2(n_609), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_45), .A2(n_53), .B1(n_364), .B2(n_372), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_46), .A2(n_140), .B1(n_382), .B2(n_894), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_47), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_48), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_50), .A2(n_181), .B1(n_383), .B2(n_579), .Y(n_629) );
AO22x2_ASAP7_75t_L g315 ( .A1(n_52), .A2(n_105), .B1(n_312), .B2(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g841 ( .A(n_52), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_54), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_55), .Y(n_497) );
AOI22xp33_ASAP7_75t_SL g854 ( .A1(n_57), .A2(n_232), .B1(n_528), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_58), .A2(n_220), .B1(n_364), .B2(n_574), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_59), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_60), .B(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_61), .A2(n_206), .B1(n_533), .B2(n_535), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_62), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_63), .A2(n_222), .B1(n_578), .B2(n_609), .Y(n_666) );
AOI222xp33_ASAP7_75t_L g470 ( .A1(n_64), .A2(n_167), .B1(n_178), .B2(n_331), .C1(n_471), .C2(n_472), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_65), .A2(n_101), .B1(n_392), .B2(n_533), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_66), .A2(n_107), .B1(n_459), .B2(n_716), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_67), .A2(n_119), .B1(n_386), .B2(n_403), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_68), .A2(n_170), .B1(n_442), .B2(n_504), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_69), .A2(n_90), .B1(n_577), .B2(n_579), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_70), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_71), .A2(n_240), .B1(n_349), .B2(n_468), .Y(n_592) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_72), .A2(n_245), .B1(n_604), .B2(n_605), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_73), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_74), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_75), .A2(n_192), .B1(n_501), .B2(n_529), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_76), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_77), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_78), .A2(n_133), .B1(n_337), .B2(n_343), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_79), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_80), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_81), .A2(n_145), .B1(n_390), .B2(n_392), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_82), .A2(n_152), .B1(n_337), .B2(n_444), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_83), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_84), .Y(n_721) );
XNOR2x2_ASAP7_75t_L g447 ( .A(n_85), .B(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_86), .A2(n_212), .B1(n_370), .B2(n_375), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_88), .A2(n_271), .B1(n_442), .B2(n_443), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_92), .Y(n_679) );
AOI222xp33_ASAP7_75t_L g538 ( .A1(n_93), .A2(n_179), .B1(n_188), .B2(n_329), .C1(n_443), .C2(n_468), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_94), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_95), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_96), .A2(n_130), .B1(n_404), .B2(n_570), .Y(n_569) );
AOI222xp33_ASAP7_75t_L g647 ( .A1(n_97), .A2(n_104), .B1(n_141), .B2(n_331), .C1(n_507), .C2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_98), .A2(n_202), .B1(n_535), .B2(n_671), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_99), .A2(n_173), .B1(n_776), .B2(n_777), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_100), .A2(n_168), .B1(n_344), .B2(n_507), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_103), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_106), .A2(n_399), .B1(n_445), .B2(n_446), .Y(n_398) );
INVx1_ASAP7_75t_L g445 ( .A(n_106), .Y(n_445) );
INVx1_ASAP7_75t_L g294 ( .A(n_108), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_109), .A2(n_205), .B1(n_411), .B2(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g877 ( .A(n_110), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_110), .A2(n_877), .B1(n_880), .B2(n_897), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_111), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_113), .A2(n_282), .B1(n_607), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_115), .A2(n_283), .B1(n_579), .B2(n_607), .Y(n_639) );
INVx1_ASAP7_75t_L g290 ( .A(n_116), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_117), .A2(n_254), .B1(n_456), .B2(n_457), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_118), .A2(n_191), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_120), .A2(n_127), .B1(n_520), .B2(n_521), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_121), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_122), .A2(n_203), .B1(n_456), .B2(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_123), .A2(n_256), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_124), .A2(n_249), .B1(n_664), .B2(n_665), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_125), .A2(n_276), .B1(n_350), .B2(n_617), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_128), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_129), .A2(n_175), .B1(n_577), .B2(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_131), .A2(n_136), .B1(n_529), .B2(n_617), .Y(n_693) );
OA22x2_ASAP7_75t_L g681 ( .A1(n_132), .A2(n_682), .B1(n_683), .B2(n_701), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_132), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_134), .B(n_430), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_137), .B(n_464), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_139), .A2(n_144), .B1(n_516), .B2(n_517), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_142), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_147), .A2(n_154), .B1(n_509), .B2(n_510), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_148), .A2(n_180), .B1(n_365), .B2(n_570), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_150), .A2(n_264), .B1(n_411), .B2(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_153), .A2(n_189), .B1(n_390), .B2(n_483), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_155), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_156), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_157), .B(n_427), .Y(n_619) );
XNOR2x2_ASAP7_75t_L g478 ( .A(n_158), .B(n_479), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_160), .A2(n_182), .B1(n_566), .B2(n_567), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_161), .Y(n_714) );
AND2x2_ASAP7_75t_L g293 ( .A(n_162), .B(n_294), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_163), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_164), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_166), .A2(n_171), .B1(n_386), .B2(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_169), .B(n_690), .Y(n_689) );
AOI222xp33_ASAP7_75t_L g735 ( .A1(n_172), .A2(n_230), .B1(n_263), .B2(n_329), .C1(n_499), .C2(n_559), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_174), .Y(n_791) );
AND2x6_ASAP7_75t_L g289 ( .A(n_176), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_176), .Y(n_834) );
AO22x2_ASAP7_75t_L g321 ( .A1(n_177), .A2(n_235), .B1(n_312), .B2(n_316), .Y(n_321) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_183), .A2(n_250), .B1(n_504), .B2(n_505), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_184), .B(n_510), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_185), .Y(n_557) );
INVx1_ASAP7_75t_L g562 ( .A(n_186), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_187), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_193), .A2(n_201), .B1(n_344), .B2(n_471), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_194), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g700 ( .A1(n_195), .A2(n_270), .B1(n_383), .B2(n_671), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_196), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_197), .A2(n_217), .B1(n_364), .B2(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_198), .A2(n_259), .B1(n_362), .B2(n_665), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_199), .A2(n_285), .B1(n_365), .B2(n_600), .Y(n_599) );
AO22x2_ASAP7_75t_L g319 ( .A1(n_200), .A2(n_257), .B1(n_312), .B2(n_313), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_204), .B(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_207), .A2(n_238), .B1(n_372), .B2(n_579), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_208), .A2(n_219), .B1(n_485), .B2(n_516), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_209), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_210), .A2(n_258), .B1(n_444), .B2(n_471), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_211), .A2(n_262), .B1(n_380), .B2(n_384), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_213), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_214), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_215), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_216), .A2(n_237), .B1(n_444), .B2(n_617), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_218), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_221), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_223), .Y(n_804) );
INVx1_ASAP7_75t_L g461 ( .A(n_224), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_226), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_227), .B(n_526), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_228), .A2(n_706), .B1(n_736), .B2(n_737), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_228), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_229), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_231), .B(n_472), .Y(n_787) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_233), .A2(n_287), .B(n_295), .C(n_842), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_235), .B(n_839), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_239), .Y(n_789) );
INVx1_ASAP7_75t_L g660 ( .A(n_242), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_243), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_244), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g763 ( .A(n_246), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_248), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_251), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_252), .Y(n_406) );
INVx1_ASAP7_75t_L g837 ( .A(n_257), .Y(n_837) );
XNOR2x2_ASAP7_75t_L g635 ( .A(n_260), .B(n_636), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_261), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_265), .Y(n_782) );
OA22x2_ASAP7_75t_SL g542 ( .A1(n_266), .A2(n_543), .B1(n_544), .B2(n_580), .Y(n_542) );
INVx1_ASAP7_75t_L g580 ( .A(n_266), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_267), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_268), .A2(n_766), .B1(n_792), .B2(n_793), .Y(n_765) );
INVx1_ASAP7_75t_L g792 ( .A(n_268), .Y(n_792) );
INVx1_ASAP7_75t_L g312 ( .A(n_273), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_273), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g615 ( .A(n_275), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_277), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_280), .Y(n_786) );
OA22x2_ASAP7_75t_L g796 ( .A1(n_281), .A2(n_797), .B1(n_798), .B2(n_799), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_281), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_284), .Y(n_753) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_290), .Y(n_833) );
OAI21xp5_ASAP7_75t_L g875 ( .A1(n_291), .A2(n_832), .B(n_876), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_652), .B1(n_653), .B2(n_828), .C(n_829), .Y(n_295) );
INVx1_ASAP7_75t_L g828 ( .A(n_296), .Y(n_828) );
XNOR2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_541), .Y(n_296) );
XNOR2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_394), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
XNOR2x1_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_360), .Y(n_301) );
NOR3xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_327), .C(n_347), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B1(n_322), .B2(n_323), .Y(n_303) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_307), .A2(n_524), .B1(n_782), .B2(n_783), .Y(n_781) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g549 ( .A(n_308), .Y(n_549) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_308), .A2(n_553), .B1(n_673), .B2(n_674), .C(n_675), .Y(n_672) );
BUFx3_ASAP7_75t_L g747 ( .A(n_308), .Y(n_747) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_317), .Y(n_308) );
INVx2_ASAP7_75t_L g393 ( .A(n_309), .Y(n_393) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_315), .Y(n_309) );
AND2x2_ASAP7_75t_L g326 ( .A(n_310), .B(n_315), .Y(n_326) );
AND2x2_ASAP7_75t_L g368 ( .A(n_310), .B(n_341), .Y(n_368) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g332 ( .A(n_311), .B(n_315), .Y(n_332) );
AND2x2_ASAP7_75t_L g342 ( .A(n_311), .B(n_321), .Y(n_342) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g316 ( .A(n_314), .Y(n_316) );
INVx2_ASAP7_75t_L g341 ( .A(n_315), .Y(n_341) );
INVx1_ASAP7_75t_L g346 ( .A(n_315), .Y(n_346) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_318), .B(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g383 ( .A(n_318), .B(n_368), .Y(n_383) );
AND2x4_ASAP7_75t_L g429 ( .A(n_318), .B(n_393), .Y(n_429) );
AND2x6_ASAP7_75t_L g431 ( .A(n_318), .B(n_326), .Y(n_431) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g334 ( .A(n_319), .Y(n_334) );
INVx1_ASAP7_75t_L g340 ( .A(n_319), .Y(n_340) );
INVx1_ASAP7_75t_L g358 ( .A(n_319), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_319), .B(n_321), .Y(n_378) );
AND2x2_ASAP7_75t_L g333 ( .A(n_320), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g367 ( .A(n_321), .B(n_358), .Y(n_367) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g462 ( .A(n_324), .Y(n_462) );
INVx1_ASAP7_75t_SL g524 ( .A(n_324), .Y(n_524) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g553 ( .A(n_325), .Y(n_553) );
AND2x4_ASAP7_75t_L g364 ( .A(n_326), .B(n_333), .Y(n_364) );
AND2x2_ASAP7_75t_L g374 ( .A(n_326), .B(n_367), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_326), .B(n_367), .Y(n_408) );
OAI21xp33_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_335), .B(n_336), .Y(n_327) );
OAI221xp5_ASAP7_75t_L g554 ( .A1(n_328), .A2(n_555), .B1(n_556), .B2(n_557), .C(n_558), .Y(n_554) );
OAI221xp5_ASAP7_75t_L g784 ( .A1(n_328), .A2(n_556), .B1(n_785), .B2(n_786), .C(n_787), .Y(n_784) );
OAI21xp5_ASAP7_75t_SL g848 ( .A1(n_328), .A2(n_849), .B(n_850), .Y(n_848) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI21xp5_ASAP7_75t_SL g749 ( .A1(n_330), .A2(n_750), .B(n_751), .Y(n_749) );
INVx4_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g496 ( .A(n_331), .Y(n_496) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_331), .Y(n_591) );
BUFx3_ASAP7_75t_L g678 ( .A(n_331), .Y(n_678) );
AND2x6_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g355 ( .A(n_332), .Y(n_355) );
AND2x4_ASAP7_75t_L g469 ( .A(n_332), .B(n_357), .Y(n_469) );
AND2x2_ASAP7_75t_L g391 ( .A(n_333), .B(n_368), .Y(n_391) );
AND2x6_ASAP7_75t_L g392 ( .A(n_333), .B(n_393), .Y(n_392) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_337), .Y(n_442) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx4f_ASAP7_75t_SL g471 ( .A(n_338), .Y(n_471) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_338), .Y(n_501) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_338), .Y(n_528) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_342), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g351 ( .A(n_340), .Y(n_351) );
INVx1_ASAP7_75t_L g437 ( .A(n_341), .Y(n_437) );
AND2x4_ASAP7_75t_L g344 ( .A(n_342), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g350 ( .A(n_342), .B(n_351), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_342), .B(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g467 ( .A(n_344), .Y(n_467) );
BUFx3_ASAP7_75t_L g529 ( .A(n_344), .Y(n_529) );
BUFx2_ASAP7_75t_L g855 ( .A(n_344), .Y(n_855) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x6_ASAP7_75t_L g377 ( .A(n_346), .B(n_378), .Y(n_377) );
OAI22xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_352), .B1(n_353), .B2(n_359), .Y(n_347) );
INVx1_ASAP7_75t_L g648 ( .A(n_348), .Y(n_648) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g559 ( .A(n_349), .Y(n_559) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx12f_ASAP7_75t_L g444 ( .A(n_350), .Y(n_444) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_350), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_353), .A2(n_434), .B1(n_561), .B2(n_562), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_353), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_788) );
BUFx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g440 ( .A(n_354), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_354), .A2(n_436), .B1(n_733), .B2(n_734), .Y(n_732) );
OR2x6_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND4x1_ASAP7_75t_L g360 ( .A(n_361), .B(n_369), .C(n_379), .D(n_389), .Y(n_360) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_363), .A2(n_422), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g516 ( .A(n_363), .Y(n_516) );
INVx2_ASAP7_75t_L g604 ( .A(n_363), .Y(n_604) );
INVx2_ASAP7_75t_L g894 ( .A(n_363), .Y(n_894) );
INVx6_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g420 ( .A(n_364), .Y(n_420) );
BUFx3_ASAP7_75t_L g669 ( .A(n_364), .Y(n_669) );
INVx1_ASAP7_75t_L g778 ( .A(n_365), .Y(n_778) );
BUFx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx3_ASAP7_75t_L g457 ( .A(n_366), .Y(n_457) );
BUFx3_ASAP7_75t_L g533 ( .A(n_366), .Y(n_533) );
BUFx3_ASAP7_75t_L g575 ( .A(n_366), .Y(n_575) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_367), .B(n_368), .Y(n_424) );
AND2x4_ASAP7_75t_L g387 ( .A(n_368), .B(n_388), .Y(n_387) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_372), .Y(n_485) );
INVx4_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g459 ( .A(n_373), .Y(n_459) );
BUFx3_ASAP7_75t_L g518 ( .A(n_373), .Y(n_518) );
INVx5_ASAP7_75t_L g578 ( .A(n_373), .Y(n_578) );
INVx3_ASAP7_75t_L g605 ( .A(n_373), .Y(n_605) );
INVx1_ASAP7_75t_L g815 ( .A(n_373), .Y(n_815) );
INVx8_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
BUFx2_ASAP7_75t_L g521 ( .A(n_376), .Y(n_521) );
BUFx2_ASAP7_75t_L g716 ( .A(n_376), .Y(n_716) );
INVx6_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g579 ( .A(n_377), .Y(n_579) );
INVx1_ASAP7_75t_SL g896 ( .A(n_377), .Y(n_896) );
INVx1_ASAP7_75t_L g388 ( .A(n_378), .Y(n_388) );
INVx4_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g453 ( .A(n_381), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_381), .A2(n_487), .B1(n_488), .B2(n_490), .Y(n_486) );
INVx4_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g520 ( .A(n_383), .Y(n_520) );
BUFx3_ASAP7_75t_L g568 ( .A(n_383), .Y(n_568) );
INVx2_ASAP7_75t_L g608 ( .A(n_383), .Y(n_608) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_385), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_708) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g404 ( .A(n_387), .Y(n_404) );
BUFx2_ASAP7_75t_SL g483 ( .A(n_387), .Y(n_483) );
BUFx3_ASAP7_75t_L g537 ( .A(n_387), .Y(n_537) );
BUFx3_ASAP7_75t_L g626 ( .A(n_387), .Y(n_626) );
BUFx2_ASAP7_75t_SL g646 ( .A(n_387), .Y(n_646) );
BUFx2_ASAP7_75t_L g671 ( .A(n_387), .Y(n_671) );
AND2x2_ASAP7_75t_L g609 ( .A(n_388), .B(n_437), .Y(n_609) );
BUFx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_391), .Y(n_403) );
INVx2_ASAP7_75t_L g536 ( .A(n_391), .Y(n_536) );
BUFx2_ASAP7_75t_SL g820 ( .A(n_391), .Y(n_820) );
INVx11_ASAP7_75t_L g416 ( .A(n_392), .Y(n_416) );
INVx11_ASAP7_75t_L g571 ( .A(n_392), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_475), .B2(n_476), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI22xp5_ASAP7_75t_SL g396 ( .A1(n_397), .A2(n_398), .B1(n_447), .B2(n_474), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g446 ( .A(n_399), .Y(n_446) );
AND4x1_ASAP7_75t_L g399 ( .A(n_400), .B(n_412), .C(n_425), .D(n_441), .Y(n_399) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_403), .Y(n_456) );
BUFx3_ASAP7_75t_L g566 ( .A(n_403), .Y(n_566) );
BUFx3_ASAP7_75t_L g770 ( .A(n_403), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B1(n_409), .B2(n_410), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_407), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
BUFx2_ASAP7_75t_R g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g451 ( .A(n_416), .Y(n_451) );
INVx5_ASAP7_75t_SL g489 ( .A(n_416), .Y(n_489) );
INVx1_ASAP7_75t_L g532 ( .A(n_416), .Y(n_532) );
INVx4_ASAP7_75t_L g600 ( .A(n_416), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_421), .B2(n_422), .Y(n_417) );
INVx2_ASAP7_75t_L g776 ( .A(n_419), .Y(n_776) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_422), .A2(n_824), .B1(n_825), .B2(n_826), .Y(n_823) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g722 ( .A(n_423), .Y(n_722) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx5_ASAP7_75t_L g464 ( .A(n_428), .Y(n_464) );
INVx2_ASAP7_75t_L g509 ( .A(n_428), .Y(n_509) );
INVx2_ASAP7_75t_L g526 ( .A(n_428), .Y(n_526) );
INVx4_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx4f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g510 ( .A(n_431), .Y(n_510) );
INVx1_ASAP7_75t_SL g691 ( .A(n_431), .Y(n_691) );
BUFx2_ASAP7_75t_L g731 ( .A(n_431), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_438), .B2(n_439), .Y(n_432) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_436), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_752) );
BUFx3_ASAP7_75t_L g790 ( .A(n_436), .Y(n_790) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g754 ( .A(n_442), .Y(n_754) );
BUFx4f_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g852 ( .A(n_444), .Y(n_852) );
INVx1_ASAP7_75t_L g474 ( .A(n_447), .Y(n_474) );
NAND4xp75_ASAP7_75t_L g448 ( .A(n_449), .B(n_454), .C(n_460), .D(n_470), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_458), .Y(n_454) );
BUFx4f_ASAP7_75t_SL g861 ( .A(n_457), .Y(n_861) );
OA211x2_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_463), .C(n_465), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_462), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_745) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_464), .Y(n_730) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g504 ( .A(n_467), .Y(n_504) );
BUFx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_469), .Y(n_507) );
BUFx2_ASAP7_75t_SL g617 ( .A(n_469), .Y(n_617) );
BUFx4f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B1(n_511), .B2(n_540), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_480), .B(n_494), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_486), .C(n_491), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
INVx2_ASAP7_75t_L g771 ( .A(n_488), .Y(n_771) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_489), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_502), .Y(n_494) );
OAI21xp5_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_497), .B(n_498), .Y(n_495) );
OAI21xp5_ASAP7_75t_SL g614 ( .A1(n_496), .A2(n_615), .B(n_616), .Y(n_614) );
OAI21xp5_ASAP7_75t_SL g882 ( .A1(n_496), .A2(n_883), .B(n_884), .Y(n_882) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g556 ( .A(n_501), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_508), .Y(n_502) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g540 ( .A(n_511), .Y(n_540) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
XOR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_539), .Y(n_512) );
NAND4xp75_ASAP7_75t_L g513 ( .A(n_514), .B(n_522), .C(n_530), .D(n_538), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OA211x2_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_525), .C(n_527), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_528), .Y(n_810) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_534), .Y(n_530) );
INVx2_ASAP7_75t_L g824 ( .A(n_532), .Y(n_824) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx3_ASAP7_75t_L g664 ( .A(n_536), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_581), .B1(n_650), .B2(n_651), .Y(n_541) );
INVx2_ASAP7_75t_L g650 ( .A(n_542), .Y(n_650) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_SL g544 ( .A(n_545), .B(n_563), .Y(n_544) );
NOR3xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_554), .C(n_560), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_550), .B2(n_551), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g802 ( .A(n_549), .Y(n_802) );
OAI22xp5_ASAP7_75t_SL g801 ( .A1(n_551), .A2(n_802), .B1(n_803), .B2(n_804), .Y(n_801) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_572), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_565), .B(n_569), .Y(n_564) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g728 ( .A(n_568), .Y(n_728) );
INVx4_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx4_ASAP7_75t_L g665 ( .A(n_571), .Y(n_665) );
INVx3_ASAP7_75t_L g860 ( .A(n_571), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g651 ( .A(n_581), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B1(n_632), .B2(n_633), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI22x1_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B1(n_611), .B2(n_631), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_584), .A2(n_585), .B1(n_635), .B2(n_649), .Y(n_634) );
INVx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
XOR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_610), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_587), .B(n_597), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_593), .Y(n_587) );
OAI21xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_592), .Y(n_588) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .C(n_596), .Y(n_593) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_602), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .Y(n_602) );
INVxp67_ASAP7_75t_L g720 ( .A(n_604), .Y(n_720) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx3_ASAP7_75t_L g631 ( .A(n_611), .Y(n_631) );
XOR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_630), .Y(n_611) );
NAND2x1_ASAP7_75t_SL g612 ( .A(n_613), .B(n_622), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_618), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .C(n_621), .Y(n_618) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_623), .B(n_627), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
BUFx2_ASAP7_75t_L g773 ( .A(n_626), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g649 ( .A(n_635), .Y(n_649) );
NAND4xp75_ASAP7_75t_L g636 ( .A(n_637), .B(n_640), .C(n_643), .D(n_647), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_641), .B(n_642), .Y(n_640) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_SL g822 ( .A(n_646), .Y(n_822) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
XNOR2xp5_ASAP7_75t_SL g653 ( .A(n_654), .B(n_738), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_658), .B1(n_704), .B2(n_705), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_681), .B1(n_702), .B2(n_703), .Y(n_658) );
INVx2_ASAP7_75t_SL g702 ( .A(n_659), .Y(n_702) );
XNOR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NOR4xp75_ASAP7_75t_L g661 ( .A(n_662), .B(n_667), .C(n_672), .D(n_676), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVxp67_ASAP7_75t_L g710 ( .A(n_664), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_668), .B(n_670), .Y(n_667) );
OAI21xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_679), .B(n_680), .Y(n_676) );
OAI21xp5_ASAP7_75t_SL g685 ( .A1(n_677), .A2(n_686), .B(n_687), .Y(n_685) );
OAI21xp33_ASAP7_75t_L g805 ( .A1(n_677), .A2(n_806), .B(n_807), .Y(n_805) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g703 ( .A(n_681), .Y(n_703) );
INVx1_ASAP7_75t_L g701 ( .A(n_683), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_694), .Y(n_683) );
NOR2xp67_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_692), .C(n_693), .Y(n_688) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
NOR2x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g737 ( .A(n_706), .Y(n_737) );
AND4x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_717), .C(n_729), .D(n_735), .Y(n_706) );
NOR2xp33_ASAP7_75t_SL g707 ( .A(n_708), .B(n_712), .Y(n_707) );
INVxp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_723), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_727), .B2(n_728), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B1(n_794), .B2(n_795), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_742), .B1(n_764), .B2(n_765), .Y(n_740) );
OAI22xp5_ASAP7_75t_SL g795 ( .A1(n_741), .A2(n_742), .B1(n_796), .B2(n_827), .Y(n_795) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
XOR2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_763), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_756), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_749), .C(n_752), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_760), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g793 ( .A(n_766), .Y(n_793) );
AND2x2_ASAP7_75t_SL g766 ( .A(n_767), .B(n_780), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_774), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_772), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_779), .Y(n_774) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NOR3xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_784), .C(n_788), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g808 ( .A1(n_790), .A2(n_809), .B1(n_810), .B2(n_811), .Y(n_808) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g827 ( .A(n_796), .Y(n_827) );
INVx2_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_812), .Y(n_799) );
NOR3xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_805), .C(n_808), .Y(n_800) );
NOR3xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_817), .C(n_823), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_819), .B1(n_821), .B2(n_822), .Y(n_817) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_SL g829 ( .A(n_830), .Y(n_829) );
NOR2x1_ASAP7_75t_L g830 ( .A(n_831), .B(n_835), .Y(n_830) );
OR2x2_ASAP7_75t_SL g900 ( .A(n_831), .B(n_836), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_832), .B(n_834), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_832), .Y(n_869) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_833), .B(n_873), .Y(n_876) );
CKINVDCx16_ASAP7_75t_R g873 ( .A(n_834), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .Y(n_839) );
OAI322xp33_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_868), .A3(n_870), .B1(n_874), .B2(n_877), .C1(n_878), .C2(n_898), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_844), .Y(n_867) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_SL g845 ( .A(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_SL g846 ( .A(n_847), .B(n_857), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_848), .B(n_853), .Y(n_847) );
INVx3_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_856), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_858), .B(n_863), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_862), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
BUFx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
BUFx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_875), .Y(n_874) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx2_ASAP7_75t_SL g897 ( .A(n_880), .Y(n_897) );
AND2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_888), .Y(n_880) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_885), .Y(n_881) );
NAND2xp5_ASAP7_75t_SL g885 ( .A(n_886), .B(n_887), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_892), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_893), .B(n_895), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_899), .Y(n_898) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_900), .Y(n_899) );
endmodule