module real_aes_10274_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1584;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1280;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_0), .A2(n_149), .B1(n_374), .B2(n_461), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_0), .A2(n_149), .B1(n_526), .B2(n_597), .Y(n_967) );
AO221x1_ASAP7_75t_L g1310 ( .A1(n_1), .A2(n_127), .B1(n_1274), .B2(n_1311), .C(n_1313), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_2), .A2(n_75), .B1(n_541), .B2(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g620 ( .A(n_2), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g1502 ( .A(n_3), .Y(n_1502) );
AOI22xp5_ASAP7_75t_L g1298 ( .A1(n_4), .A2(n_112), .B1(n_1274), .B2(n_1280), .Y(n_1298) );
INVx1_ASAP7_75t_L g899 ( .A(n_5), .Y(n_899) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_6), .A2(n_15), .B1(n_651), .B2(n_653), .Y(n_650) );
INVxp67_ASAP7_75t_SL g702 ( .A(n_6), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_7), .A2(n_160), .B1(n_464), .B2(n_465), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_7), .A2(n_160), .B1(n_851), .B2(n_855), .Y(n_1073) );
INVx1_ASAP7_75t_L g586 ( .A(n_8), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_8), .A2(n_233), .B1(n_531), .B2(n_600), .Y(n_599) );
INVxp33_ASAP7_75t_SL g640 ( .A(n_9), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_9), .A2(n_281), .B1(n_673), .B2(n_675), .Y(n_672) );
INVxp33_ASAP7_75t_SL g1189 ( .A(n_10), .Y(n_1189) );
AOI22xp5_ASAP7_75t_SL g1215 ( .A1(n_10), .A2(n_252), .B1(n_653), .B2(n_1216), .Y(n_1215) );
INVx1_ASAP7_75t_L g509 ( .A(n_11), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_11), .A2(n_60), .B1(n_447), .B2(n_536), .Y(n_535) );
AO22x1_ASAP7_75t_L g1171 ( .A1(n_12), .A2(n_1172), .B1(n_1173), .B2(n_1218), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_12), .Y(n_1172) );
AOI22xp33_ASAP7_75t_SL g964 ( .A1(n_13), .A2(n_263), .B1(n_464), .B2(n_965), .Y(n_964) );
INVxp67_ASAP7_75t_L g974 ( .A(n_13), .Y(n_974) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_14), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_14), .A2(n_203), .B1(n_410), .B2(n_413), .Y(n_698) );
INVxp67_ASAP7_75t_SL g703 ( .A(n_15), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g1197 ( .A1(n_16), .A2(n_209), .B1(n_1022), .B2(n_1198), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_16), .A2(n_209), .B1(n_1211), .B2(n_1214), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_17), .A2(n_202), .B1(n_795), .B2(n_1238), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_17), .A2(n_202), .B1(n_1164), .B2(n_1244), .Y(n_1243) );
INVx1_ASAP7_75t_L g1314 ( .A(n_18), .Y(n_1314) );
INVx1_ASAP7_75t_L g1232 ( .A(n_19), .Y(n_1232) );
OAI22xp5_ASAP7_75t_L g1256 ( .A1(n_19), .A2(n_220), .B1(n_618), .B2(n_759), .Y(n_1256) );
INVx1_ASAP7_75t_L g1099 ( .A(n_20), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_20), .A2(n_284), .B1(n_828), .B2(n_833), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_21), .A2(n_307), .B1(n_374), .B2(n_461), .Y(n_609) );
INVx1_ASAP7_75t_L g615 ( .A(n_21), .Y(n_615) );
XOR2x2_ASAP7_75t_L g627 ( .A(n_22), .B(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_23), .A2(n_67), .B1(n_728), .B2(n_1014), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_23), .A2(n_67), .B1(n_1026), .B2(n_1028), .Y(n_1025) );
INVxp67_ASAP7_75t_SL g912 ( .A(n_24), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_24), .A2(n_199), .B1(n_653), .B2(n_664), .Y(n_937) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_25), .A2(n_229), .B1(n_440), .B2(n_441), .Y(n_524) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_25), .A2(n_229), .B1(n_541), .B2(n_542), .Y(n_540) );
OAI211xp5_ASAP7_75t_L g835 ( .A1(n_26), .A2(n_573), .B(n_836), .C(n_839), .Y(n_835) );
INVx1_ASAP7_75t_L g862 ( .A(n_26), .Y(n_862) );
INVx1_ASAP7_75t_L g997 ( .A(n_27), .Y(n_997) );
INVx1_ASAP7_75t_L g434 ( .A(n_28), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_28), .A2(n_183), .B1(n_464), .B2(n_475), .Y(n_474) );
OAI222xp33_ASAP7_75t_L g1496 ( .A1(n_29), .A2(n_61), .B1(n_130), .B2(n_384), .C1(n_1497), .C2(n_1498), .Y(n_1496) );
INVx1_ASAP7_75t_L g1512 ( .A(n_29), .Y(n_1512) );
INVx1_ASAP7_75t_L g949 ( .A(n_30), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_30), .A2(n_33), .B1(n_618), .B2(n_759), .Y(n_971) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_31), .A2(n_80), .B1(n_795), .B2(n_796), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_31), .A2(n_80), .B1(n_664), .B2(n_816), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_32), .Y(n_874) );
INVx1_ASAP7_75t_L g950 ( .A(n_33), .Y(n_950) );
INVx1_ASAP7_75t_L g487 ( .A(n_34), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_34), .A2(n_147), .B1(n_464), .B2(n_475), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_35), .A2(n_303), .B1(n_1250), .B2(n_1251), .Y(n_1249) );
INVxp67_ASAP7_75t_SL g1259 ( .A(n_35), .Y(n_1259) );
INVx1_ASAP7_75t_L g318 ( .A(n_36), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g1050 ( .A1(n_37), .A2(n_214), .B1(n_734), .B2(n_795), .C(n_1051), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_37), .A2(n_214), .B1(n_464), .B2(n_475), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1574 ( .A1(n_38), .A2(n_54), .B1(n_327), .B2(n_429), .Y(n_1574) );
OAI22xp33_ASAP7_75t_L g1583 ( .A1(n_38), .A2(n_298), .B1(n_828), .B2(n_833), .Y(n_1583) );
INVx1_ASAP7_75t_L g1183 ( .A(n_39), .Y(n_1183) );
INVx1_ASAP7_75t_L g952 ( .A(n_40), .Y(n_952) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_41), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_41), .A2(n_176), .B1(n_531), .B2(n_918), .Y(n_1158) );
AOI22xp5_ASAP7_75t_L g1324 ( .A1(n_42), .A2(n_132), .B1(n_1274), .B2(n_1280), .Y(n_1324) );
AOI22xp33_ASAP7_75t_SL g1236 ( .A1(n_43), .A2(n_171), .B1(n_724), .B2(n_725), .Y(n_1236) );
AOI22xp33_ASAP7_75t_SL g1246 ( .A1(n_43), .A2(n_171), .B1(n_589), .B2(n_1247), .Y(n_1246) );
INVxp33_ASAP7_75t_L g791 ( .A(n_44), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_44), .A2(n_253), .B1(n_539), .B2(n_813), .Y(n_819) );
INVxp33_ASAP7_75t_SL g1194 ( .A(n_45), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_45), .A2(n_250), .B1(n_947), .B2(n_1211), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_46), .A2(n_273), .B1(n_440), .B2(n_1552), .Y(n_1551) );
AOI22xp33_ASAP7_75t_L g1560 ( .A1(n_46), .A2(n_273), .B1(n_542), .B2(n_652), .Y(n_1560) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_47), .A2(n_179), .B1(n_443), .B2(n_447), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_47), .A2(n_179), .B1(n_374), .B2(n_461), .Y(n_460) );
INVxp33_ASAP7_75t_SL g900 ( .A(n_48), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_48), .A2(n_181), .B1(n_531), .B2(n_918), .Y(n_917) );
INVxp33_ASAP7_75t_SL g914 ( .A(n_49), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_49), .A2(n_65), .B1(n_747), .B2(n_932), .Y(n_936) );
AO221x2_ASAP7_75t_L g1357 ( .A1(n_50), .A2(n_241), .B1(n_1311), .B2(n_1358), .C(n_1360), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_51), .A2(n_73), .B1(n_851), .B2(n_855), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_51), .A2(n_73), .B1(n_652), .B2(n_1164), .Y(n_1167) );
INVxp67_ASAP7_75t_SL g993 ( .A(n_52), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_52), .A2(n_63), .B1(n_475), .B2(n_1033), .Y(n_1032) );
INVxp67_ASAP7_75t_SL g713 ( .A(n_53), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_53), .A2(n_197), .B1(n_733), .B2(n_734), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g1563 ( .A1(n_54), .A2(n_167), .B1(n_963), .B2(n_1564), .Y(n_1563) );
INVx1_ASAP7_75t_L g1064 ( .A(n_55), .Y(n_1064) );
OAI211xp5_ASAP7_75t_L g1043 ( .A1(n_56), .A2(n_573), .B(n_1044), .C(n_1045), .Y(n_1043) );
INVx1_ASAP7_75t_L g1058 ( .A(n_56), .Y(n_1058) );
INVx1_ASAP7_75t_L g1515 ( .A(n_57), .Y(n_1515) );
AOI22xp33_ASAP7_75t_SL g1532 ( .A1(n_57), .A2(n_98), .B1(n_813), .B2(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g490 ( .A(n_58), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_58), .A2(n_162), .B1(n_546), .B2(n_548), .Y(n_545) );
OAI211xp5_ASAP7_75t_L g555 ( .A1(n_58), .A2(n_504), .B(n_556), .C(n_561), .Y(n_555) );
XNOR2xp5_ASAP7_75t_L g577 ( .A(n_59), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g513 ( .A(n_60), .Y(n_513) );
OAI211xp5_ASAP7_75t_L g567 ( .A1(n_60), .A2(n_568), .B(n_573), .C(n_574), .Y(n_567) );
AOI22xp33_ASAP7_75t_SL g1518 ( .A1(n_61), .A2(n_261), .B1(n_802), .B2(n_920), .Y(n_1518) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_62), .A2(n_262), .B1(n_1274), .B2(n_1280), .Y(n_1336) );
INVxp67_ASAP7_75t_SL g1000 ( .A(n_63), .Y(n_1000) );
AOI22xp5_ASAP7_75t_L g1292 ( .A1(n_64), .A2(n_293), .B1(n_1293), .B2(n_1296), .Y(n_1292) );
INVxp67_ASAP7_75t_SL g908 ( .A(n_65), .Y(n_908) );
INVx1_ASAP7_75t_L g510 ( .A(n_66), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_66), .A2(n_287), .B1(n_531), .B2(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g1572 ( .A(n_68), .Y(n_1572) );
CKINVDCx5p33_ASAP7_75t_R g1120 ( .A(n_69), .Y(n_1120) );
AO22x1_ASAP7_75t_L g1319 ( .A1(n_70), .A2(n_225), .B1(n_1280), .B2(n_1320), .Y(n_1319) );
AO22x1_ASAP7_75t_L g1321 ( .A1(n_71), .A2(n_224), .B1(n_1293), .B2(n_1296), .Y(n_1321) );
INVx1_ASAP7_75t_L g1182 ( .A(n_72), .Y(n_1182) );
AOI22xp33_ASAP7_75t_SL g1204 ( .A1(n_72), .A2(n_108), .B1(n_725), .B2(n_1198), .Y(n_1204) );
AOI221xp5_ASAP7_75t_L g867 ( .A1(n_74), .A2(n_234), .B1(n_868), .B2(n_869), .C(n_871), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_74), .A2(n_234), .B1(n_475), .B2(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g622 ( .A(n_75), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_76), .A2(n_86), .B1(n_927), .B2(n_929), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_76), .A2(n_86), .B1(n_747), .B2(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g1179 ( .A(n_77), .Y(n_1179) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_78), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_79), .A2(n_221), .B1(n_851), .B2(n_855), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_79), .A2(n_221), .B1(n_465), .B2(n_884), .Y(n_889) );
BUFx2_ASAP7_75t_L g394 ( .A(n_81), .Y(n_394) );
BUFx2_ASAP7_75t_L g436 ( .A(n_81), .Y(n_436) );
INVx1_ASAP7_75t_L g683 ( .A(n_81), .Y(n_683) );
INVx1_ASAP7_75t_L g1230 ( .A(n_82), .Y(n_1230) );
AOI22xp33_ASAP7_75t_SL g1241 ( .A1(n_82), .A2(n_177), .B1(n_724), .B2(n_736), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_83), .A2(n_223), .B1(n_645), .B2(n_648), .Y(n_644) );
INVxp67_ASAP7_75t_SL g697 ( .A(n_83), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_84), .A2(n_300), .B1(n_664), .B2(n_666), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_84), .A2(n_300), .B1(n_673), .B2(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g902 ( .A(n_85), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_85), .A2(n_105), .B1(n_491), .B2(n_920), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1553 ( .A1(n_87), .A2(n_283), .B1(n_443), .B2(n_491), .Y(n_1553) );
AOI22xp33_ASAP7_75t_L g1559 ( .A1(n_87), .A2(n_283), .B1(n_374), .B2(n_962), .Y(n_1559) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_88), .A2(n_247), .B1(n_648), .B2(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_88), .A2(n_247), .B1(n_616), .B2(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g361 ( .A(n_89), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_89), .A2(n_305), .B1(n_441), .B2(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_90), .A2(n_246), .B1(n_531), .B2(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_90), .A2(n_246), .B1(n_607), .B2(n_934), .Y(n_933) );
XNOR2xp5_ASAP7_75t_L g1131 ( .A(n_91), .B(n_1132), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_92), .A2(n_274), .B1(n_491), .B2(n_724), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_92), .A2(n_274), .B1(n_749), .B2(n_963), .Y(n_1024) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_93), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_94), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_95), .A2(n_304), .B1(n_962), .B2(n_963), .Y(n_961) );
INVxp33_ASAP7_75t_L g976 ( .A(n_95), .Y(n_976) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_96), .A2(n_222), .B1(n_831), .B2(n_834), .Y(n_1048) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_96), .A2(n_222), .B1(n_728), .B2(n_1019), .C(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1509 ( .A(n_97), .Y(n_1509) );
AOI22xp33_ASAP7_75t_L g1534 ( .A1(n_97), .A2(n_192), .B1(n_822), .B2(n_934), .Y(n_1534) );
INVx1_ASAP7_75t_L g1511 ( .A(n_98), .Y(n_1511) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_99), .A2(n_106), .B1(n_379), .B2(n_384), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_99), .A2(n_106), .B1(n_410), .B2(n_413), .Y(n_409) );
AO221x1_ASAP7_75t_L g1273 ( .A1(n_100), .A2(n_114), .B1(n_1274), .B2(n_1280), .C(n_1281), .Y(n_1273) );
INVx1_ASAP7_75t_L g1186 ( .A(n_101), .Y(n_1186) );
AO221x1_ASAP7_75t_L g1303 ( .A1(n_102), .A2(n_279), .B1(n_1274), .B2(n_1280), .C(n_1304), .Y(n_1303) );
AO22x2_ASAP7_75t_L g1491 ( .A1(n_102), .A2(n_1492), .B1(n_1493), .B2(n_1537), .Y(n_1491) );
INVxp67_ASAP7_75t_SL g1492 ( .A(n_102), .Y(n_1492) );
AOI22xp5_ASAP7_75t_L g1543 ( .A1(n_102), .A2(n_1544), .B1(n_1585), .B2(n_1589), .Y(n_1543) );
INVx1_ASAP7_75t_L g1306 ( .A(n_103), .Y(n_1306) );
INVx1_ASAP7_75t_L g1052 ( .A(n_104), .Y(n_1052) );
INVxp33_ASAP7_75t_SL g896 ( .A(n_105), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_107), .A2(n_139), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_107), .A2(n_139), .B1(n_472), .B2(n_539), .Y(n_538) );
INVxp33_ASAP7_75t_SL g1176 ( .A(n_108), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1523 ( .A1(n_109), .A2(n_184), .B1(n_920), .B2(n_1524), .Y(n_1523) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_109), .A2(n_184), .B1(n_813), .B2(n_1528), .Y(n_1527) );
CKINVDCx5p33_ASAP7_75t_R g872 ( .A(n_110), .Y(n_872) );
AO22x2_ASAP7_75t_L g939 ( .A1(n_111), .A2(n_940), .B1(n_977), .B2(n_978), .Y(n_939) );
INVx1_ASAP7_75t_L g977 ( .A(n_111), .Y(n_977) );
INVx1_ASAP7_75t_L g1047 ( .A(n_113), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g1323 ( .A1(n_115), .A2(n_138), .B1(n_1293), .B2(n_1296), .Y(n_1323) );
INVxp33_ASAP7_75t_SL g788 ( .A(n_116), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_116), .A2(n_200), .B1(n_821), .B2(n_822), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_117), .A2(n_227), .B1(n_648), .B2(n_749), .Y(n_748) );
INVxp67_ASAP7_75t_SL g757 ( .A(n_117), .Y(n_757) );
XOR2xp5_ASAP7_75t_L g1080 ( .A(n_118), .B(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_119), .A2(n_271), .B1(n_475), .B2(n_884), .Y(n_956) );
AOI22xp33_ASAP7_75t_SL g966 ( .A1(n_119), .A2(n_271), .B1(n_440), .B2(n_441), .Y(n_966) );
INVx1_ASAP7_75t_L g1361 ( .A(n_120), .Y(n_1361) );
INVx1_ASAP7_75t_L g585 ( .A(n_121), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_121), .A2(n_235), .B1(n_491), .B2(n_536), .Y(n_601) );
INVx1_ASAP7_75t_L g717 ( .A(n_122), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_122), .A2(n_264), .B1(n_618), .B2(n_759), .Y(n_758) );
INVxp33_ASAP7_75t_L g1003 ( .A(n_123), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_123), .A2(n_169), .B1(n_724), .B2(n_1022), .Y(n_1021) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_124), .A2(n_259), .B1(n_800), .B2(n_802), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_124), .A2(n_259), .B1(n_645), .B2(n_813), .Y(n_812) );
INVxp33_ASAP7_75t_SL g775 ( .A(n_125), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_125), .A2(n_296), .B1(n_805), .B2(n_807), .Y(n_804) );
INVxp67_ASAP7_75t_SL g946 ( .A(n_126), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_126), .A2(n_196), .B1(n_443), .B2(n_597), .Y(n_959) );
INVx1_ASAP7_75t_L g992 ( .A(n_128), .Y(n_992) );
INVx1_ASAP7_75t_L g1097 ( .A(n_129), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_129), .A2(n_254), .B1(n_831), .B2(n_834), .Y(n_1122) );
INVx1_ASAP7_75t_L g1513 ( .A(n_130), .Y(n_1513) );
INVxp33_ASAP7_75t_SL g944 ( .A(n_131), .Y(n_944) );
AOI22xp33_ASAP7_75t_SL g958 ( .A1(n_131), .A2(n_278), .B1(n_440), .B2(n_441), .Y(n_958) );
INVx1_ASAP7_75t_L g1279 ( .A(n_133), .Y(n_1279) );
OAI211xp5_ASAP7_75t_L g1147 ( .A1(n_134), .A2(n_504), .B(n_1126), .C(n_1148), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_134), .A2(n_232), .B1(n_461), .B2(n_1162), .Y(n_1166) );
INVxp33_ASAP7_75t_SL g709 ( .A(n_135), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_135), .A2(n_172), .B1(n_724), .B2(n_736), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_136), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_137), .A2(n_210), .B1(n_1153), .B2(n_1154), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_137), .A2(n_210), .B1(n_652), .B2(n_1164), .Y(n_1163) );
XOR2x2_ASAP7_75t_L g1220 ( .A(n_138), .B(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1305 ( .A(n_140), .Y(n_1305) );
CKINVDCx20_ASAP7_75t_R g995 ( .A(n_141), .Y(n_995) );
INVx1_ASAP7_75t_L g781 ( .A(n_142), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_142), .A2(n_249), .B1(n_495), .B2(n_618), .Y(n_786) );
AO22x2_ASAP7_75t_SL g704 ( .A1(n_143), .A2(n_705), .B1(n_706), .B2(n_765), .Y(n_704) );
CKINVDCx16_ASAP7_75t_R g705 ( .A(n_143), .Y(n_705) );
INVx1_ASAP7_75t_L g1111 ( .A(n_144), .Y(n_1111) );
OAI22xp33_ASAP7_75t_SL g1129 ( .A1(n_144), .A2(n_157), .B1(n_327), .B2(n_851), .Y(n_1129) );
INVxp33_ASAP7_75t_SL g631 ( .A(n_145), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_145), .A2(n_155), .B1(n_616), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_146), .A2(n_256), .B1(n_532), .B2(n_728), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_146), .A2(n_256), .B1(n_1207), .B2(n_1208), .Y(n_1206) );
INVx1_ASAP7_75t_L g488 ( .A(n_147), .Y(n_488) );
INVx1_ASAP7_75t_L g1277 ( .A(n_148), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_148), .B(n_1287), .Y(n_1289) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_150), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_151), .A2(n_206), .B1(n_526), .B2(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_151), .A2(n_206), .B1(n_374), .B2(n_461), .Y(n_603) );
INVxp33_ASAP7_75t_SL g1177 ( .A(n_152), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_152), .A2(n_217), .B1(n_728), .B2(n_1202), .Y(n_1201) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_153), .A2(n_163), .B1(n_828), .B2(n_831), .Y(n_827) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_153), .A2(n_267), .B1(n_728), .B2(n_730), .C(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g330 ( .A(n_154), .Y(n_330) );
INVxp67_ASAP7_75t_SL g634 ( .A(n_155), .Y(n_634) );
INVxp33_ASAP7_75t_L g774 ( .A(n_156), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_156), .A2(n_289), .B1(n_597), .B2(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_157), .A2(n_248), .B1(n_465), .B2(n_652), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1521 ( .A1(n_158), .A2(n_236), .B1(n_795), .B2(n_1522), .Y(n_1521) );
AOI22xp33_ASAP7_75t_L g1529 ( .A1(n_158), .A2(n_236), .B1(n_822), .B2(n_1530), .Y(n_1529) );
AOI22xp33_ASAP7_75t_SL g1248 ( .A1(n_159), .A2(n_269), .B1(n_747), .B2(n_749), .Y(n_1248) );
INVxp33_ASAP7_75t_SL g1261 ( .A(n_159), .Y(n_1261) );
BUFx3_ASAP7_75t_L g353 ( .A(n_161), .Y(n_353) );
INVx1_ASAP7_75t_L g371 ( .A(n_161), .Y(n_371) );
INVx1_ASAP7_75t_L g501 ( .A(n_162), .Y(n_501) );
INVx1_ASAP7_75t_L g859 ( .A(n_163), .Y(n_859) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_164), .A2(n_216), .B1(n_440), .B2(n_441), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_164), .A2(n_216), .B1(n_464), .B2(n_465), .Y(n_463) );
INVx1_ASAP7_75t_L g344 ( .A(n_165), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_165), .A2(n_270), .B1(n_443), .B2(n_447), .Y(n_454) );
INVxp33_ASAP7_75t_L g999 ( .A(n_166), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_166), .A2(n_219), .B1(n_749), .B2(n_1036), .Y(n_1035) );
OAI211xp5_ASAP7_75t_SL g1567 ( .A1(n_167), .A2(n_504), .B(n_1568), .C(n_1571), .Y(n_1567) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_168), .A2(n_212), .B1(n_728), .B2(n_730), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_168), .A2(n_212), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g1008 ( .A(n_169), .Y(n_1008) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_170), .A2(n_306), .B1(n_724), .B2(n_725), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_170), .A2(n_306), .B1(n_746), .B2(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g715 ( .A(n_172), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g1557 ( .A1(n_173), .A2(n_298), .B1(n_491), .B2(n_526), .Y(n_1557) );
INVx1_ASAP7_75t_L g1578 ( .A(n_173), .Y(n_1578) );
INVx1_ASAP7_75t_L g1315 ( .A(n_174), .Y(n_1315) );
INVx1_ASAP7_75t_L g1140 ( .A(n_175), .Y(n_1140) );
INVx1_ASAP7_75t_L g1143 ( .A(n_176), .Y(n_1143) );
INVxp33_ASAP7_75t_SL g1224 ( .A(n_177), .Y(n_1224) );
XNOR2xp5_ASAP7_75t_L g824 ( .A(n_178), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g1363 ( .A(n_180), .Y(n_1363) );
INVxp33_ASAP7_75t_SL g897 ( .A(n_181), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_182), .A2(n_251), .B1(n_828), .B2(n_833), .Y(n_1042) );
INVx1_ASAP7_75t_L g1072 ( .A(n_182), .Y(n_1072) );
INVx1_ASAP7_75t_L g426 ( .A(n_183), .Y(n_426) );
INVx1_ASAP7_75t_L g392 ( .A(n_185), .Y(n_392) );
INVx1_ASAP7_75t_L g1573 ( .A(n_186), .Y(n_1573) );
INVx1_ASAP7_75t_L g592 ( .A(n_187), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g617 ( .A1(n_187), .A2(n_285), .B1(n_495), .B2(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_SL g1093 ( .A(n_188), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_188), .A2(n_290), .B1(n_465), .B2(n_541), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_189), .A2(n_301), .B1(n_440), .B2(n_441), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_189), .A2(n_301), .B1(n_605), .B2(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g1282 ( .A(n_190), .Y(n_1282) );
AOI22xp5_ASAP7_75t_L g1337 ( .A1(n_191), .A2(n_311), .B1(n_1293), .B2(n_1296), .Y(n_1337) );
INVx1_ASAP7_75t_L g1508 ( .A(n_192), .Y(n_1508) );
CKINVDCx14_ASAP7_75t_R g1039 ( .A(n_193), .Y(n_1039) );
INVx1_ASAP7_75t_L g1046 ( .A(n_194), .Y(n_1046) );
INVx1_ASAP7_75t_L g1227 ( .A(n_195), .Y(n_1227) );
INVxp33_ASAP7_75t_SL g943 ( .A(n_196), .Y(n_943) );
INVxp33_ASAP7_75t_SL g710 ( .A(n_197), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g1562 ( .A1(n_198), .A2(n_260), .B1(n_541), .B2(n_607), .Y(n_1562) );
OAI22xp5_ASAP7_75t_L g1566 ( .A1(n_198), .A2(n_260), .B1(n_851), .B2(n_855), .Y(n_1566) );
INVxp33_ASAP7_75t_L g911 ( .A(n_199), .Y(n_911) );
INVxp67_ASAP7_75t_SL g789 ( .A(n_200), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_201), .A2(n_267), .B1(n_833), .B2(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g849 ( .A(n_201), .Y(n_849) );
INVxp67_ASAP7_75t_SL g637 ( .A(n_203), .Y(n_637) );
INVx1_ASAP7_75t_L g712 ( .A(n_204), .Y(n_712) );
INVx1_ASAP7_75t_L g1088 ( .A(n_205), .Y(n_1088) );
INVx1_ASAP7_75t_L g639 ( .A(n_207), .Y(n_639) );
INVx1_ASAP7_75t_L g1139 ( .A(n_208), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1545 ( .A1(n_211), .A2(n_1546), .B1(n_1547), .B2(n_1584), .Y(n_1545) );
CKINVDCx5p33_ASAP7_75t_R g1546 ( .A(n_211), .Y(n_1546) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_213), .A2(n_238), .B1(n_491), .B2(n_526), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_213), .A2(n_238), .B1(n_539), .B2(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1054 ( .A(n_215), .Y(n_1054) );
INVxp33_ASAP7_75t_SL g1180 ( .A(n_217), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1555 ( .A1(n_218), .A2(n_243), .B1(n_440), .B2(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1582 ( .A(n_218), .Y(n_1582) );
INVxp67_ASAP7_75t_SL g996 ( .A(n_219), .Y(n_996) );
INVx1_ASAP7_75t_L g1233 ( .A(n_220), .Y(n_1233) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_223), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_226), .Y(n_845) );
INVxp33_ASAP7_75t_L g764 ( .A(n_227), .Y(n_764) );
BUFx3_ASAP7_75t_L g355 ( .A(n_228), .Y(n_355) );
INVx1_ASAP7_75t_L g366 ( .A(n_228), .Y(n_366) );
INVx1_ASAP7_75t_L g1065 ( .A(n_230), .Y(n_1065) );
INVxp67_ASAP7_75t_SL g1228 ( .A(n_231), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_231), .A2(n_239), .B1(n_728), .B2(n_734), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_232), .A2(n_286), .B1(n_327), .B2(n_429), .Y(n_1149) );
INVx1_ASAP7_75t_L g582 ( .A(n_233), .Y(n_582) );
INVx1_ASAP7_75t_L g588 ( .A(n_235), .Y(n_588) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_237), .Y(n_326) );
INVx1_ASAP7_75t_L g458 ( .A(n_237), .Y(n_458) );
INVxp33_ASAP7_75t_SL g1225 ( .A(n_239), .Y(n_1225) );
CKINVDCx5p33_ASAP7_75t_R g1121 ( .A(n_240), .Y(n_1121) );
INVx2_ASAP7_75t_L g348 ( .A(n_242), .Y(n_348) );
INVxp67_ASAP7_75t_SL g1581 ( .A(n_243), .Y(n_1581) );
INVx1_ASAP7_75t_L g777 ( .A(n_244), .Y(n_777) );
INVx1_ASAP7_75t_L g904 ( .A(n_245), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_245), .A2(n_276), .B1(n_413), .B2(n_759), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_248), .A2(n_284), .B1(n_429), .B2(n_855), .Y(n_1124) );
INVx1_ASAP7_75t_L g782 ( .A(n_249), .Y(n_782) );
INVx1_ASAP7_75t_L g1192 ( .A(n_250), .Y(n_1192) );
INVx1_ASAP7_75t_L g1057 ( .A(n_251), .Y(n_1057) );
INVxp33_ASAP7_75t_SL g1190 ( .A(n_252), .Y(n_1190) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_253), .Y(n_785) );
INVx1_ASAP7_75t_L g1095 ( .A(n_254), .Y(n_1095) );
INVx1_ASAP7_75t_L g1505 ( .A(n_255), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g1519 ( .A1(n_255), .A2(n_266), .B1(n_805), .B2(n_1154), .Y(n_1519) );
AO22x2_ASAP7_75t_L g483 ( .A1(n_257), .A2(n_484), .B1(n_551), .B2(n_552), .Y(n_483) );
INVxp67_ASAP7_75t_L g551 ( .A(n_257), .Y(n_551) );
INVx1_ASAP7_75t_L g1112 ( .A(n_258), .Y(n_1112) );
OAI211xp5_ASAP7_75t_SL g1125 ( .A1(n_258), .A2(n_504), .B(n_1126), .C(n_1128), .Y(n_1125) );
INVx1_ASAP7_75t_L g1501 ( .A(n_261), .Y(n_1501) );
INVxp33_ASAP7_75t_L g973 ( .A(n_263), .Y(n_973) );
INVx1_ASAP7_75t_L g718 ( .A(n_264), .Y(n_718) );
INVx1_ASAP7_75t_L g418 ( .A(n_265), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_265), .A2(n_295), .B1(n_461), .B2(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g1504 ( .A(n_266), .Y(n_1504) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_268), .Y(n_502) );
INVxp67_ASAP7_75t_SL g1255 ( .A(n_269), .Y(n_1255) );
INVx1_ASAP7_75t_L g377 ( .A(n_270), .Y(n_377) );
INVx1_ASAP7_75t_L g988 ( .A(n_272), .Y(n_988) );
OAI22xp33_ASAP7_75t_L g1144 ( .A1(n_275), .A2(n_286), .B1(n_828), .B2(n_833), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_275), .A2(n_297), .B1(n_536), .B2(n_929), .Y(n_1159) );
INVx1_ASAP7_75t_L g903 ( .A(n_276), .Y(n_903) );
INVxp67_ASAP7_75t_SL g1004 ( .A(n_277), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_277), .A2(n_294), .B1(n_733), .B2(n_1019), .Y(n_1018) );
INVxp33_ASAP7_75t_SL g953 ( .A(n_278), .Y(n_953) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_280), .Y(n_320) );
AND3x2_ASAP7_75t_L g1278 ( .A(n_280), .B(n_318), .C(n_1279), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_280), .B(n_318), .Y(n_1285) );
INVxp33_ASAP7_75t_SL g632 ( .A(n_281), .Y(n_632) );
INVx2_ASAP7_75t_L g331 ( .A(n_282), .Y(n_331) );
INVx1_ASAP7_75t_L g590 ( .A(n_285), .Y(n_590) );
INVx1_ASAP7_75t_L g518 ( .A(n_287), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g840 ( .A(n_288), .Y(n_840) );
INVxp67_ASAP7_75t_SL g780 ( .A(n_289), .Y(n_780) );
INVxp67_ASAP7_75t_SL g1090 ( .A(n_290), .Y(n_1090) );
INVx1_ASAP7_75t_L g1087 ( .A(n_291), .Y(n_1087) );
INVx1_ASAP7_75t_L g333 ( .A(n_292), .Y(n_333) );
INVx2_ASAP7_75t_L g408 ( .A(n_292), .Y(n_408) );
XNOR2xp5_ASAP7_75t_L g340 ( .A(n_293), .B(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_SL g1006 ( .A(n_294), .Y(n_1006) );
INVx1_ASAP7_75t_L g397 ( .A(n_295), .Y(n_397) );
INVxp33_ASAP7_75t_L g778 ( .A(n_296), .Y(n_778) );
INVx1_ASAP7_75t_L g1136 ( .A(n_297), .Y(n_1136) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_299), .Y(n_841) );
XOR2x2_ASAP7_75t_L g892 ( .A(n_302), .B(n_893), .Y(n_892) );
INVxp33_ASAP7_75t_SL g1258 ( .A(n_303), .Y(n_1258) );
INVxp67_ASAP7_75t_SL g970 ( .A(n_304), .Y(n_970) );
INVx1_ASAP7_75t_L g367 ( .A(n_305), .Y(n_367) );
INVx1_ASAP7_75t_L g624 ( .A(n_307), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_308), .A2(n_310), .B1(n_752), .B2(n_753), .Y(n_751) );
INVxp33_ASAP7_75t_L g761 ( .A(n_308), .Y(n_761) );
INVx1_ASAP7_75t_L g1101 ( .A(n_309), .Y(n_1101) );
INVxp67_ASAP7_75t_SL g762 ( .A(n_310), .Y(n_762) );
AO22x1_ASAP7_75t_L g769 ( .A1(n_311), .A2(n_770), .B1(n_771), .B2(n_823), .Y(n_769) );
INVxp67_ASAP7_75t_L g770 ( .A(n_311), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_334), .B(n_1263), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_321), .Y(n_315) );
AND2x4_ASAP7_75t_L g1542 ( .A(n_316), .B(n_322), .Y(n_1542) );
NOR2xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_SL g1588 ( .A(n_317), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1594 ( .A(n_317), .B(n_319), .Y(n_1594) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_319), .B(n_1588), .Y(n_1587) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g435 ( .A(n_324), .B(n_436), .Y(n_435) );
OR2x6_ASAP7_75t_L g506 ( .A(n_324), .B(n_436), .Y(n_506) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g450 ( .A(n_325), .B(n_333), .Y(n_450) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g1085 ( .A(n_326), .B(n_421), .Y(n_1085) );
INVx8_ASAP7_75t_L g417 ( .A(n_327), .Y(n_417) );
OR2x6_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .Y(n_327) );
OR2x6_ASAP7_75t_L g429 ( .A(n_328), .B(n_420), .Y(n_429) );
INVx2_ASAP7_75t_SL g861 ( .A(n_328), .Y(n_861) );
BUFx6f_ASAP7_75t_L g873 ( .A(n_328), .Y(n_873) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_328), .Y(n_1053) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g402 ( .A(n_330), .Y(n_402) );
INVx1_ASAP7_75t_L g415 ( .A(n_330), .Y(n_415) );
INVx2_ASAP7_75t_L g423 ( .A(n_330), .Y(n_423) );
AND2x4_ASAP7_75t_L g433 ( .A(n_330), .B(n_403), .Y(n_433) );
AND2x2_ASAP7_75t_L g446 ( .A(n_330), .B(n_331), .Y(n_446) );
INVx2_ASAP7_75t_L g403 ( .A(n_331), .Y(n_403) );
INVx1_ASAP7_75t_L g412 ( .A(n_331), .Y(n_412) );
INVx1_ASAP7_75t_L g425 ( .A(n_331), .Y(n_425) );
INVx1_ASAP7_75t_L g560 ( .A(n_331), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_331), .B(n_423), .Y(n_854) );
AND2x4_ASAP7_75t_L g411 ( .A(n_332), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g413 ( .A(n_333), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g618 ( .A(n_333), .B(n_414), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B1(n_983), .B2(n_1262), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
XNOR2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_479), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_390), .B(n_395), .C(n_437), .Y(n_341) );
NAND4xp25_ASAP7_75t_L g342 ( .A(n_343), .B(n_360), .C(n_372), .D(n_387), .Y(n_342) );
AOI22xp5_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_345), .B1(n_356), .B2(n_357), .Y(n_343) );
AOI22xp5_ASAP7_75t_SL g508 ( .A1(n_345), .A2(n_362), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_345), .A2(n_362), .B1(n_774), .B2(n_775), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_345), .A2(n_362), .B1(n_1224), .B2(n_1225), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1500 ( .A1(n_345), .A2(n_357), .B1(n_1501), .B2(n_1502), .Y(n_1500) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
AND2x6_ASAP7_75t_L g368 ( .A(n_346), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g584 ( .A(n_346), .B(n_349), .Y(n_584) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g380 ( .A(n_347), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_348), .Y(n_359) );
INVx1_ASAP7_75t_L g364 ( .A(n_348), .Y(n_364) );
AND2x2_ASAP7_75t_L g469 ( .A(n_348), .B(n_392), .Y(n_469) );
INVx2_ASAP7_75t_L g478 ( .A(n_348), .Y(n_478) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_350), .Y(n_547) );
INVx2_ASAP7_75t_SL g647 ( .A(n_350), .Y(n_647) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_350), .Y(n_662) );
INVx2_ASAP7_75t_L g750 ( .A(n_350), .Y(n_750) );
INVx2_ASAP7_75t_L g1213 ( .A(n_350), .Y(n_1213) );
INVx1_ASAP7_75t_L g1533 ( .A(n_350), .Y(n_1533) );
INVx1_ASAP7_75t_L g1564 ( .A(n_350), .Y(n_1564) );
INVx6_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g357 ( .A(n_351), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g462 ( .A(n_351), .Y(n_462) );
BUFx2_ASAP7_75t_L g539 ( .A(n_351), .Y(n_539) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g386 ( .A(n_352), .Y(n_386) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g365 ( .A(n_353), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g376 ( .A(n_353), .B(n_355), .Y(n_376) );
INVx1_ASAP7_75t_L g383 ( .A(n_354), .Y(n_383) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g370 ( .A(n_355), .B(n_371), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_356), .A2(n_428), .B1(n_430), .B2(n_434), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_357), .A2(n_368), .B1(n_502), .B2(n_518), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_357), .A2(n_368), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_357), .A2(n_368), .B1(n_639), .B2(n_640), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_357), .A2(n_368), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_357), .A2(n_368), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx4_ASAP7_75t_L g833 ( .A(n_357), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_357), .A2(n_368), .B1(n_899), .B2(n_900), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_357), .A2(n_368), .B1(n_952), .B2(n_953), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_357), .A2(n_368), .B1(n_992), .B2(n_1006), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_357), .A2(n_368), .B1(n_1179), .B2(n_1180), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_357), .A2(n_368), .B1(n_1227), .B2(n_1228), .Y(n_1226) );
AND2x4_ASAP7_75t_L g515 ( .A(n_358), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_358), .B(n_516), .Y(n_591) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B1(n_367), .B2(n_368), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_362), .A2(n_584), .B1(n_585), .B2(n_586), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_362), .A2(n_388), .B1(n_584), .B2(n_631), .C(n_632), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_362), .A2(n_584), .B1(n_709), .B2(n_710), .Y(n_708) );
CKINVDCx6p67_ASAP7_75t_R g831 ( .A(n_362), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_362), .A2(n_584), .B1(n_896), .B2(n_897), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_362), .A2(n_584), .B1(n_943), .B2(n_944), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_362), .A2(n_584), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_362), .A2(n_368), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_362), .A2(n_584), .B1(n_1176), .B2(n_1177), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_362), .A2(n_368), .B1(n_1504), .B2(n_1505), .Y(n_1503) );
AOI22xp5_ASAP7_75t_L g1580 ( .A1(n_362), .A2(n_368), .B1(n_1581), .B2(n_1582), .Y(n_1580) );
AND2x6_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
AND2x2_ASAP7_75t_L g373 ( .A(n_363), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g389 ( .A(n_363), .Y(n_389) );
INVx1_ASAP7_75t_L g829 ( .A(n_363), .Y(n_829) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x6_ASAP7_75t_L g385 ( .A(n_364), .B(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g464 ( .A(n_365), .Y(n_464) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_365), .Y(n_541) );
INVx2_ASAP7_75t_SL g606 ( .A(n_365), .Y(n_606) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_365), .Y(n_652) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_365), .Y(n_665) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_365), .Y(n_742) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_365), .Y(n_821) );
BUFx6f_ASAP7_75t_L g884 ( .A(n_365), .Y(n_884) );
BUFx2_ASAP7_75t_L g934 ( .A(n_365), .Y(n_934) );
BUFx2_ASAP7_75t_L g1530 ( .A(n_365), .Y(n_1530) );
INVx1_ASAP7_75t_L g572 ( .A(n_366), .Y(n_572) );
INVx4_ASAP7_75t_L g834 ( .A(n_368), .Y(n_834) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_369), .Y(n_475) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_369), .Y(n_607) );
INVx1_ASAP7_75t_L g612 ( .A(n_369), .Y(n_612) );
INVx1_ASAP7_75t_L g667 ( .A(n_369), .Y(n_667) );
INVx1_ASAP7_75t_L g817 ( .A(n_369), .Y(n_817) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_370), .Y(n_465) );
INVx1_ASAP7_75t_L g543 ( .A(n_370), .Y(n_543) );
INVx2_ASAP7_75t_L g656 ( .A(n_370), .Y(n_656) );
INVx1_ASAP7_75t_L g744 ( .A(n_370), .Y(n_744) );
INVx1_ASAP7_75t_L g571 ( .A(n_371), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_377), .B(n_378), .Y(n_372) );
INVx1_ASAP7_75t_L g1044 ( .A(n_373), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_374), .Y(n_512) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_374), .Y(n_716) );
HB1xp67_ASAP7_75t_L g1231 ( .A(n_374), .Y(n_1231) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g388 ( .A(n_375), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g549 ( .A(n_375), .Y(n_549) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_375), .Y(n_649) );
INVx2_ASAP7_75t_L g814 ( .A(n_375), .Y(n_814) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_376), .Y(n_473) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI222xp33_ASAP7_75t_L g1117 ( .A1(n_380), .A2(n_385), .B1(n_1101), .B2(n_1118), .C1(n_1120), .C2(n_1121), .Y(n_1117) );
INVx2_ASAP7_75t_L g1497 ( .A(n_380), .Y(n_1497) );
AOI222xp33_ASAP7_75t_L g1577 ( .A1(n_380), .A2(n_385), .B1(n_1572), .B2(n_1573), .C1(n_1578), .C2(n_1579), .Y(n_1577) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g516 ( .A(n_382), .Y(n_516) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI222xp33_ASAP7_75t_L g511 ( .A1(n_385), .A2(n_493), .B1(n_496), .B2(n_512), .C1(n_513), .C2(n_514), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_385), .A2(n_493), .B1(n_496), .B2(n_515), .Y(n_574) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_385), .A2(n_588), .B1(n_589), .B2(n_590), .C1(n_591), .C2(n_592), .Y(n_587) );
AOI222xp33_ASAP7_75t_L g633 ( .A1(n_385), .A2(n_591), .B1(n_634), .B2(n_635), .C1(n_636), .C2(n_637), .Y(n_633) );
AOI222xp33_ASAP7_75t_L g714 ( .A1(n_385), .A2(n_514), .B1(n_715), .B2(n_716), .C1(n_717), .C2(n_718), .Y(n_714) );
AOI222xp33_ASAP7_75t_L g779 ( .A1(n_385), .A2(n_472), .B1(n_591), .B2(n_780), .C1(n_781), .C2(n_782), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_385), .A2(n_515), .B1(n_840), .B2(n_841), .Y(n_839) );
AOI222xp33_ASAP7_75t_L g901 ( .A1(n_385), .A2(n_591), .B1(n_648), .B2(n_902), .C1(n_903), .C2(n_904), .Y(n_901) );
AOI222xp33_ASAP7_75t_L g945 ( .A1(n_385), .A2(n_591), .B1(n_946), .B2(n_947), .C1(n_949), .C2(n_950), .Y(n_945) );
AOI222xp33_ASAP7_75t_L g1007 ( .A1(n_385), .A2(n_514), .B1(n_995), .B2(n_997), .C1(n_1008), .C2(n_1009), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_385), .A2(n_515), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
AOI222xp33_ASAP7_75t_L g1135 ( .A1(n_385), .A2(n_591), .B1(n_1136), .B2(n_1137), .C1(n_1139), .C2(n_1140), .Y(n_1135) );
AOI222xp33_ASAP7_75t_L g1181 ( .A1(n_385), .A2(n_589), .B1(n_1182), .B2(n_1183), .C1(n_1184), .C2(n_1186), .Y(n_1181) );
AOI222xp33_ASAP7_75t_L g1229 ( .A1(n_385), .A2(n_514), .B1(n_1230), .B2(n_1231), .C1(n_1232), .C2(n_1233), .Y(n_1229) );
NAND4xp25_ASAP7_75t_L g507 ( .A(n_387), .B(n_508), .C(n_511), .D(n_517), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g579 ( .A(n_387), .B(n_580), .C(n_583), .D(n_587), .Y(n_579) );
NAND4xp25_ASAP7_75t_SL g707 ( .A(n_387), .B(n_708), .C(n_711), .D(n_714), .Y(n_707) );
NAND4xp25_ASAP7_75t_SL g772 ( .A(n_387), .B(n_773), .C(n_776), .D(n_779), .Y(n_772) );
NAND4xp25_ASAP7_75t_L g1001 ( .A(n_387), .B(n_1002), .C(n_1005), .D(n_1007), .Y(n_1001) );
NAND4xp25_ASAP7_75t_L g1174 ( .A(n_387), .B(n_1175), .C(n_1178), .D(n_1181), .Y(n_1174) );
NAND4xp25_ASAP7_75t_SL g1222 ( .A(n_387), .B(n_1223), .C(n_1226), .D(n_1229), .Y(n_1222) );
INVx5_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
CKINVDCx8_ASAP7_75t_R g573 ( .A(n_388), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g1495 ( .A(n_388), .B(n_1496), .Y(n_1495) );
AOI211xp5_ASAP7_75t_L g578 ( .A1(n_390), .A2(n_579), .B(n_593), .C(n_613), .Y(n_578) );
OAI31xp33_ASAP7_75t_SL g826 ( .A1(n_390), .A2(n_827), .A3(n_832), .B(n_835), .Y(n_826) );
AOI211x1_ASAP7_75t_L g940 ( .A1(n_390), .A2(n_941), .B(n_954), .C(n_968), .Y(n_940) );
OAI31xp33_ASAP7_75t_L g1041 ( .A1(n_390), .A2(n_1042), .A3(n_1043), .B(n_1048), .Y(n_1041) );
OAI31xp33_ASAP7_75t_SL g1114 ( .A1(n_390), .A2(n_1115), .A3(n_1116), .B(n_1122), .Y(n_1114) );
OAI21xp5_ASAP7_75t_L g1133 ( .A1(n_390), .A2(n_1134), .B(n_1144), .Y(n_1133) );
OAI21xp5_ASAP7_75t_SL g1575 ( .A1(n_390), .A2(n_1576), .B(n_1583), .Y(n_1575) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
AND2x4_ASAP7_75t_L g520 ( .A(n_391), .B(n_393), .Y(n_520) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g477 ( .A(n_392), .B(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g449 ( .A(n_394), .Y(n_449) );
OR2x6_ASAP7_75t_L g1084 ( .A(n_394), .B(n_1085), .Y(n_1084) );
AOI31xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_416), .A3(n_427), .B(n_435), .Y(n_395) );
AOI211xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_404), .C(n_409), .Y(n_396) );
AOI222xp33_ASAP7_75t_L g1191 ( .A1(n_398), .A2(n_411), .B1(n_563), .B2(n_1183), .C1(n_1186), .C2(n_1192), .Y(n_1191) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g929 ( .A(n_399), .Y(n_929) );
INVx2_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_400), .Y(n_802) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x4_ASAP7_75t_L g404 ( .A(n_401), .B(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g447 ( .A(n_401), .Y(n_447) );
BUFx3_ASAP7_75t_L g492 ( .A(n_401), .Y(n_492) );
INVx1_ASAP7_75t_L g528 ( .A(n_401), .Y(n_528) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_401), .Y(n_597) );
BUFx2_ASAP7_75t_L g738 ( .A(n_401), .Y(n_738) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
CKINVDCx11_ASAP7_75t_R g504 ( .A(n_404), .Y(n_504) );
AOI211xp5_ASAP7_75t_L g614 ( .A1(n_404), .A2(n_615), .B(n_616), .C(n_617), .Y(n_614) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_404), .A2(n_491), .B(n_697), .C(n_698), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g756 ( .A1(n_404), .A2(n_491), .B(n_757), .C(n_758), .Y(n_756) );
AOI211xp5_ASAP7_75t_L g784 ( .A1(n_404), .A2(n_616), .B(n_785), .C(n_786), .Y(n_784) );
AOI211xp5_ASAP7_75t_L g906 ( .A1(n_404), .A2(n_907), .B(n_908), .C(n_909), .Y(n_906) );
AOI211xp5_ASAP7_75t_L g969 ( .A1(n_404), .A2(n_616), .B(n_970), .C(n_971), .Y(n_969) );
AOI211xp5_ASAP7_75t_SL g1254 ( .A1(n_404), .A2(n_527), .B(n_1255), .C(n_1256), .Y(n_1254) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g499 ( .A(n_406), .Y(n_499) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2x1p5_ASAP7_75t_L g457 ( .A(n_407), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g421 ( .A(n_408), .Y(n_421) );
INVx1_ASAP7_75t_L g562 ( .A(n_410), .Y(n_562) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g495 ( .A(n_411), .Y(n_495) );
INVx2_ASAP7_75t_L g759 ( .A(n_411), .Y(n_759) );
AOI222xp33_ASAP7_75t_SL g844 ( .A1(n_411), .A2(n_497), .B1(n_840), .B2(n_841), .C1(n_845), .C2(n_846), .Y(n_844) );
AOI222xp33_ASAP7_75t_L g1069 ( .A1(n_411), .A2(n_563), .B1(n_1046), .B2(n_1047), .C1(n_1065), .C2(n_1070), .Y(n_1069) );
AOI22xp5_ASAP7_75t_L g1128 ( .A1(n_411), .A2(n_563), .B1(n_1120), .B2(n_1121), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1571 ( .A1(n_411), .A2(n_563), .B1(n_1572), .B2(n_1573), .Y(n_1571) );
INVx1_ASAP7_75t_L g498 ( .A(n_414), .Y(n_498) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g559 ( .A(n_415), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_415), .B(n_560), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_419), .B2(n_426), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_417), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_417), .A2(n_503), .B1(n_581), .B2(n_624), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_417), .A2(n_503), .B1(n_639), .B2(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_417), .A2(n_428), .B1(n_712), .B2(n_764), .Y(n_763) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_417), .A2(n_428), .B1(n_777), .B2(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_417), .A2(n_503), .B1(n_848), .B2(n_849), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_417), .A2(n_428), .B1(n_899), .B2(n_914), .Y(n_913) );
AOI22xp33_ASAP7_75t_SL g975 ( .A1(n_417), .A2(n_428), .B1(n_952), .B2(n_976), .Y(n_975) );
AOI22xp33_ASAP7_75t_SL g998 ( .A1(n_417), .A2(n_621), .B1(n_999), .B2(n_1000), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_417), .A2(n_503), .B1(n_1064), .B2(n_1072), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_417), .A2(n_428), .B1(n_1179), .B2(n_1194), .Y(n_1193) );
AOI22xp33_ASAP7_75t_SL g1260 ( .A1(n_417), .A2(n_503), .B1(n_1227), .B2(n_1261), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g1514 ( .A1(n_417), .A2(n_428), .B1(n_1502), .B2(n_1515), .Y(n_1514) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_419), .A2(n_430), .B1(n_487), .B2(n_488), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_419), .A2(n_620), .B1(n_621), .B2(n_622), .Y(n_619) );
AOI22xp5_ASAP7_75t_SL g701 ( .A1(n_419), .A2(n_621), .B1(n_702), .B2(n_703), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_419), .A2(n_430), .B1(n_761), .B2(n_762), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_419), .A2(n_621), .B1(n_788), .B2(n_789), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_419), .A2(n_621), .B1(n_911), .B2(n_912), .Y(n_910) );
AOI22xp33_ASAP7_75t_SL g972 ( .A1(n_419), .A2(n_621), .B1(n_973), .B2(n_974), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g991 ( .A1(n_419), .A2(n_503), .B1(n_992), .B2(n_993), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_419), .A2(n_430), .B1(n_1189), .B2(n_1190), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_419), .A2(n_430), .B1(n_1258), .B2(n_1259), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1507 ( .A1(n_419), .A2(n_621), .B1(n_1508), .B2(n_1509), .Y(n_1507) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
AND2x4_ASAP7_75t_L g430 ( .A(n_420), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g621 ( .A(n_420), .B(n_431), .Y(n_621) );
INVx1_ASAP7_75t_L g852 ( .A(n_420), .Y(n_852) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_422), .Y(n_440) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_422), .Y(n_453) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_422), .Y(n_531) );
INVx1_ASAP7_75t_L g674 ( .A(n_422), .Y(n_674) );
BUFx2_ASAP7_75t_L g733 ( .A(n_422), .Y(n_733) );
BUFx2_ASAP7_75t_L g795 ( .A(n_422), .Y(n_795) );
INVx1_ASAP7_75t_L g806 ( .A(n_422), .Y(n_806) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx5_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx4_ASAP7_75t_L g503 ( .A(n_429), .Y(n_503) );
INVx5_ASAP7_75t_SL g855 ( .A(n_430), .Y(n_855) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g1203 ( .A(n_432), .Y(n_1203) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_433), .Y(n_441) );
INVx3_ASAP7_75t_L g534 ( .A(n_433), .Y(n_534) );
INVx1_ASAP7_75t_L g689 ( .A(n_433), .Y(n_689) );
AOI31xp33_ASAP7_75t_L g968 ( .A1(n_435), .A2(n_969), .A3(n_972), .B(n_975), .Y(n_968) );
AND2x4_ASAP7_75t_L g476 ( .A(n_436), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g658 ( .A(n_436), .B(n_477), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g437 ( .A(n_438), .B(n_451), .C(n_459), .D(n_470), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .C(n_448), .Y(n_438) );
INVx2_ASAP7_75t_SL g731 ( .A(n_441), .Y(n_731) );
BUFx3_ASAP7_75t_L g734 ( .A(n_441), .Y(n_734) );
INVx2_ASAP7_75t_SL g1020 ( .A(n_441), .Y(n_1020) );
INVx2_ASAP7_75t_SL g1239 ( .A(n_441), .Y(n_1239) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g526 ( .A(n_444), .Y(n_526) );
INVx2_ASAP7_75t_L g920 ( .A(n_444), .Y(n_920) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g536 ( .A(n_445), .Y(n_536) );
BUFx6f_ASAP7_75t_L g1199 ( .A(n_445), .Y(n_1199) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx3_ASAP7_75t_L g679 ( .A(n_446), .Y(n_679) );
BUFx2_ASAP7_75t_L g1070 ( .A(n_447), .Y(n_1070) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_448), .B(n_524), .C(n_525), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_448), .B(n_595), .C(n_596), .Y(n_594) );
INVx2_ASAP7_75t_L g722 ( .A(n_448), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g793 ( .A(n_448), .B(n_794), .C(n_799), .Y(n_793) );
BUFx3_ASAP7_75t_L g875 ( .A(n_448), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g921 ( .A(n_448), .B(n_922), .C(n_926), .Y(n_921) );
AOI33xp33_ASAP7_75t_L g960 ( .A1(n_448), .A2(n_476), .A3(n_961), .B1(n_964), .B2(n_966), .B3(n_967), .Y(n_960) );
NAND3xp33_ASAP7_75t_L g1151 ( .A(n_448), .B(n_1152), .C(n_1156), .Y(n_1151) );
NAND3xp33_ASAP7_75t_L g1550 ( .A(n_448), .B(n_1551), .C(n_1553), .Y(n_1550) );
AND2x4_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
AND2x2_ASAP7_75t_L g455 ( .A(n_449), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g467 ( .A(n_449), .B(n_468), .Y(n_467) );
OR2x6_ASAP7_75t_L g669 ( .A(n_449), .B(n_670), .Y(n_669) );
AND2x4_ASAP7_75t_L g694 ( .A(n_449), .B(n_450), .Y(n_694) );
OR2x2_ASAP7_75t_L g877 ( .A(n_449), .B(n_670), .Y(n_877) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .C(n_455), .Y(n_451) );
INVx2_ASAP7_75t_SL g729 ( .A(n_453), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_455), .B(n_530), .C(n_535), .Y(n_529) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_455), .B(n_599), .C(n_601), .Y(n_598) );
AOI33xp33_ASAP7_75t_L g955 ( .A1(n_455), .A2(n_466), .A3(n_956), .B1(n_957), .B2(n_958), .B3(n_959), .Y(n_955) );
INVx1_ASAP7_75t_L g1102 ( .A(n_455), .Y(n_1102) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x6_ASAP7_75t_L g681 ( .A(n_457), .B(n_682), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_463), .C(n_466), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g962 ( .A(n_462), .Y(n_962) );
INVx2_ASAP7_75t_SL g1034 ( .A(n_464), .Y(n_1034) );
BUFx3_ASAP7_75t_L g1207 ( .A(n_464), .Y(n_1207) );
BUFx6f_ASAP7_75t_L g1164 ( .A(n_465), .Y(n_1164) );
INVx1_ASAP7_75t_L g1252 ( .A(n_465), .Y(n_1252) );
NAND3xp33_ASAP7_75t_L g537 ( .A(n_466), .B(n_538), .C(n_540), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_466), .B(n_603), .C(n_604), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g811 ( .A(n_466), .B(n_812), .C(n_815), .Y(n_811) );
NAND3xp33_ASAP7_75t_L g930 ( .A(n_466), .B(n_931), .C(n_933), .Y(n_930) );
NAND3xp33_ASAP7_75t_L g1160 ( .A(n_466), .B(n_1161), .C(n_1163), .Y(n_1160) );
NAND3xp33_ASAP7_75t_L g1526 ( .A(n_466), .B(n_1527), .C(n_1529), .Y(n_1526) );
NAND3xp33_ASAP7_75t_L g1558 ( .A(n_466), .B(n_1559), .C(n_1560), .Y(n_1558) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_SL g1103 ( .A1(n_467), .A2(n_885), .B1(n_1104), .B2(n_1110), .Y(n_1103) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g670 ( .A(n_469), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_474), .C(n_476), .Y(n_470) );
BUFx2_ASAP7_75t_SL g635 ( .A(n_472), .Y(n_635) );
INVx1_ASAP7_75t_L g1037 ( .A(n_472), .Y(n_1037) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g589 ( .A(n_473), .Y(n_589) );
BUFx4f_ASAP7_75t_L g747 ( .A(n_473), .Y(n_747) );
INVx1_ASAP7_75t_L g948 ( .A(n_473), .Y(n_948) );
INVx2_ASAP7_75t_SL g1119 ( .A(n_473), .Y(n_1119) );
INVx1_ASAP7_75t_L g1138 ( .A(n_473), .Y(n_1138) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_476), .B(n_545), .C(n_550), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_476), .B(n_609), .C(n_610), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g818 ( .A(n_476), .B(n_819), .C(n_820), .Y(n_818) );
NAND3xp33_ASAP7_75t_L g935 ( .A(n_476), .B(n_936), .C(n_937), .Y(n_935) );
NAND3xp33_ASAP7_75t_L g1165 ( .A(n_476), .B(n_1166), .C(n_1167), .Y(n_1165) );
INVx1_ASAP7_75t_L g1536 ( .A(n_476), .Y(n_1536) );
NAND3xp33_ASAP7_75t_L g1561 ( .A(n_476), .B(n_1562), .C(n_1563), .Y(n_1561) );
AO22x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_767), .B1(n_981), .B2(n_982), .Y(n_479) );
INVx1_ASAP7_75t_L g981 ( .A(n_480), .Y(n_981) );
XNOR2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_625), .Y(n_480) );
AO22x2_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B1(n_576), .B2(n_577), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI221x1_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_505), .B1(n_507), .B2(n_519), .C(n_521), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_486), .B(n_489), .C(n_500), .D(n_504), .Y(n_485) );
INVx1_ASAP7_75t_L g564 ( .A(n_486), .Y(n_564) );
AOI222xp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_493), .B2(n_494), .C1(n_496), .C2(n_497), .Y(n_489) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_491), .Y(n_907) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g1525 ( .A(n_492), .Y(n_1525) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_493), .A2(n_496), .B1(n_562), .B2(n_563), .Y(n_561) );
AOI222xp33_ASAP7_75t_L g994 ( .A1(n_494), .A2(n_563), .B1(n_616), .B2(n_995), .C1(n_996), .C2(n_997), .Y(n_994) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AOI222xp33_ASAP7_75t_L g1510 ( .A1(n_497), .A2(n_562), .B1(n_1022), .B2(n_1511), .C1(n_1512), .C2(n_1513), .Y(n_1510) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
AND2x4_ASAP7_75t_L g563 ( .A(n_498), .B(n_499), .Y(n_563) );
INVx1_ASAP7_75t_L g554 ( .A(n_500), .Y(n_554) );
NAND3xp33_ASAP7_75t_SL g843 ( .A(n_504), .B(n_844), .C(n_847), .Y(n_843) );
NAND4xp25_ASAP7_75t_L g990 ( .A(n_504), .B(n_991), .C(n_994), .D(n_998), .Y(n_990) );
NAND3xp33_ASAP7_75t_L g1068 ( .A(n_504), .B(n_1069), .C(n_1071), .Y(n_1068) );
NAND4xp25_ASAP7_75t_SL g1187 ( .A(n_504), .B(n_1188), .C(n_1191), .D(n_1193), .Y(n_1187) );
NAND4xp25_ASAP7_75t_SL g1506 ( .A(n_504), .B(n_1507), .C(n_1510), .D(n_1514), .Y(n_1506) );
OAI31xp33_ASAP7_75t_L g553 ( .A1(n_505), .A2(n_554), .A3(n_555), .B(n_564), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g842 ( .A1(n_505), .A2(n_843), .B(n_850), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g893 ( .A1(n_505), .A2(n_520), .B1(n_894), .B2(n_905), .C(n_915), .Y(n_893) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_505), .A2(n_990), .B1(n_1001), .B2(n_1010), .C(n_1011), .Y(n_989) );
OAI21xp5_ASAP7_75t_L g1067 ( .A1(n_505), .A2(n_1068), .B(n_1073), .Y(n_1067) );
OAI31xp33_ASAP7_75t_SL g1123 ( .A1(n_505), .A2(n_1124), .A3(n_1125), .B(n_1129), .Y(n_1123) );
OAI31xp33_ASAP7_75t_L g1145 ( .A1(n_505), .A2(n_1146), .A3(n_1147), .B(n_1149), .Y(n_1145) );
AOI221xp5_ASAP7_75t_L g1173 ( .A1(n_505), .A2(n_520), .B1(n_1174), .B2(n_1187), .C(n_1195), .Y(n_1173) );
AOI221x1_ASAP7_75t_L g1493 ( .A1(n_505), .A2(n_519), .B1(n_1494), .B2(n_1506), .C(n_1516), .Y(n_1493) );
OAI31xp33_ASAP7_75t_SL g1565 ( .A1(n_505), .A2(n_1566), .A3(n_1567), .B(n_1574), .Y(n_1565) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
AOI31xp33_ASAP7_75t_L g613 ( .A1(n_506), .A2(n_614), .A3(n_619), .B(n_623), .Y(n_613) );
AOI31xp33_ASAP7_75t_SL g695 ( .A1(n_506), .A2(n_696), .A3(n_699), .B(n_701), .Y(n_695) );
AOI31xp33_ASAP7_75t_L g755 ( .A1(n_506), .A2(n_756), .A3(n_760), .B(n_763), .Y(n_755) );
AOI31xp33_ASAP7_75t_L g783 ( .A1(n_506), .A2(n_784), .A3(n_787), .B(n_790), .Y(n_783) );
AOI31xp33_ASAP7_75t_L g1253 ( .A1(n_506), .A2(n_1254), .A3(n_1257), .B(n_1260), .Y(n_1253) );
INVxp67_ASAP7_75t_L g566 ( .A(n_508), .Y(n_566) );
BUFx4f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g1185 ( .A(n_515), .Y(n_1185) );
INVxp67_ASAP7_75t_L g575 ( .A(n_517), .Y(n_575) );
OAI31xp33_ASAP7_75t_L g565 ( .A1(n_519), .A2(n_566), .A3(n_567), .B(n_575), .Y(n_565) );
AOI211x1_ASAP7_75t_SL g706 ( .A1(n_519), .A2(n_707), .B(n_719), .C(n_755), .Y(n_706) );
AOI211xp5_ASAP7_75t_L g771 ( .A1(n_519), .A2(n_772), .B(n_783), .C(n_792), .Y(n_771) );
AOI211xp5_ASAP7_75t_SL g1221 ( .A1(n_519), .A2(n_1222), .B(n_1234), .C(n_1253), .Y(n_1221) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g641 ( .A(n_520), .Y(n_641) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_522), .B(n_553), .C(n_565), .Y(n_552) );
AND4x1_ASAP7_75t_L g522 ( .A(n_523), .B(n_529), .C(n_537), .D(n_544), .Y(n_522) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_SL g600 ( .A(n_533), .Y(n_600) );
INVx2_ASAP7_75t_L g918 ( .A(n_533), .Y(n_918) );
INVx2_ASAP7_75t_L g1552 ( .A(n_533), .Y(n_1552) );
INVx2_ASAP7_75t_L g1556 ( .A(n_533), .Y(n_1556) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g676 ( .A(n_534), .Y(n_676) );
INVx3_ASAP7_75t_L g798 ( .A(n_534), .Y(n_798) );
BUFx3_ASAP7_75t_L g752 ( .A(n_541), .Y(n_752) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g746 ( .A(n_547), .Y(n_746) );
INVx2_ASAP7_75t_L g932 ( .A(n_547), .Y(n_932) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_558), .A2(n_872), .B1(n_873), .B2(n_874), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_558), .A2(n_1052), .B1(n_1053), .B2(n_1054), .Y(n_1051) );
OAI22xp33_ASAP7_75t_SL g1056 ( .A1(n_558), .A2(n_860), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g1100 ( .A(n_559), .Y(n_1100) );
BUFx2_ASAP7_75t_L g1127 ( .A(n_559), .Y(n_1127) );
INVx2_ASAP7_75t_L g1570 ( .A(n_559), .Y(n_1570) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_562), .A2(n_563), .B1(n_1139), .B2(n_1140), .Y(n_1148) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g1499 ( .A(n_569), .Y(n_1499) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx2_ASAP7_75t_L g838 ( .A(n_570), .Y(n_838) );
INVx2_ASAP7_75t_L g882 ( .A(n_570), .Y(n_882) );
BUFx4f_ASAP7_75t_L g888 ( .A(n_570), .Y(n_888) );
INVx1_ASAP7_75t_L g1108 ( .A(n_570), .Y(n_1108) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
OR2x2_ASAP7_75t_L g830 ( .A(n_571), .B(n_572), .Y(n_830) );
NAND4xp25_ASAP7_75t_L g894 ( .A(n_573), .B(n_895), .C(n_898), .D(n_901), .Y(n_894) );
NAND4xp25_ASAP7_75t_L g941 ( .A(n_573), .B(n_942), .C(n_945), .D(n_951), .Y(n_941) );
NAND2xp5_ASAP7_75t_SL g1116 ( .A(n_573), .B(n_1117), .Y(n_1116) );
NAND3xp33_ASAP7_75t_SL g1134 ( .A(n_573), .B(n_1135), .C(n_1141), .Y(n_1134) );
NAND3xp33_ASAP7_75t_SL g1576 ( .A(n_573), .B(n_1577), .C(n_1580), .Y(n_1576) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_594), .B(n_598), .C(n_602), .D(n_608), .Y(n_593) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_597), .Y(n_616) );
INVx2_ASAP7_75t_SL g726 ( .A(n_597), .Y(n_726) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_SL g1216 ( .A(n_606), .Y(n_1216) );
INVx1_ASAP7_75t_L g1209 ( .A(n_607), .Y(n_1209) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_704), .B2(n_766), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_642), .C(n_695), .Y(n_628) );
AOI31xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_633), .A3(n_638), .B(n_641), .Y(n_629) );
INVx1_ASAP7_75t_L g1010 ( .A(n_641), .Y(n_1010) );
NAND4xp25_ASAP7_75t_L g642 ( .A(n_643), .B(n_659), .C(n_671), .D(n_684), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_650), .C(n_657), .Y(n_643) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g1245 ( .A(n_652), .Y(n_1245) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g822 ( .A(n_654), .Y(n_822) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
BUFx2_ASAP7_75t_L g965 ( .A(n_655), .Y(n_965) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g753 ( .A(n_656), .Y(n_753) );
BUFx4f_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx4f_ASAP7_75t_L g754 ( .A(n_658), .Y(n_754) );
INVx4_ASAP7_75t_L g885 ( .A(n_658), .Y(n_885) );
AOI33xp33_ASAP7_75t_L g1205 ( .A1(n_658), .A2(n_668), .A3(n_1206), .B1(n_1210), .B2(n_1215), .B3(n_1217), .Y(n_1205) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .C(n_668), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g1247 ( .A(n_662), .Y(n_1247) );
BUFx4f_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI33xp33_ASAP7_75t_L g740 ( .A1(n_668), .A2(n_741), .A3(n_745), .B1(n_748), .B2(n_751), .B3(n_754), .Y(n_740) );
AOI33xp33_ASAP7_75t_L g1242 ( .A1(n_668), .A2(n_754), .A3(n_1243), .B1(n_1246), .B2(n_1248), .B3(n_1249), .Y(n_1242) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_669), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_669), .Y(n_1029) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_677), .C(n_680), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g868 ( .A(n_674), .Y(n_868) );
INVx1_ASAP7_75t_L g1153 ( .A(n_674), .Y(n_1153) );
BUFx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g1015 ( .A(n_676), .Y(n_1015) );
INVx2_ASAP7_75t_L g1096 ( .A(n_676), .Y(n_1096) );
BUFx3_ASAP7_75t_L g724 ( .A(n_678), .Y(n_724) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g693 ( .A(n_679), .Y(n_693) );
INVx2_ASAP7_75t_SL g801 ( .A(n_679), .Y(n_801) );
NAND3xp33_ASAP7_75t_L g803 ( .A(n_680), .B(n_804), .C(n_809), .Y(n_803) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_680), .B(n_917), .C(n_919), .Y(n_916) );
NAND3xp33_ASAP7_75t_L g1017 ( .A(n_680), .B(n_1018), .C(n_1021), .Y(n_1017) );
NAND3xp33_ASAP7_75t_L g1157 ( .A(n_680), .B(n_1158), .C(n_1159), .Y(n_1157) );
NAND3xp33_ASAP7_75t_L g1517 ( .A(n_680), .B(n_1518), .C(n_1519), .Y(n_1517) );
INVx5_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx6_ASAP7_75t_L g739 ( .A(n_681), .Y(n_739) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_690), .C(n_694), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g925 ( .A(n_689), .Y(n_925) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
BUFx2_ASAP7_75t_L g810 ( .A(n_693), .Y(n_810) );
INVx1_ASAP7_75t_L g928 ( .A(n_693), .Y(n_928) );
AOI33xp33_ASAP7_75t_L g1235 ( .A1(n_694), .A2(n_739), .A3(n_1236), .B1(n_1237), .B2(n_1240), .B3(n_1241), .Y(n_1235) );
NAND3xp33_ASAP7_75t_L g1520 ( .A(n_694), .B(n_1521), .C(n_1523), .Y(n_1520) );
INVx1_ASAP7_75t_L g766 ( .A(n_704), .Y(n_766) );
INVx1_ASAP7_75t_L g765 ( .A(n_706), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_740), .Y(n_719) );
AOI33xp33_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_723), .A3(n_727), .B1(n_732), .B2(n_735), .B3(n_739), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g1012 ( .A(n_721), .B(n_1013), .C(n_1016), .Y(n_1012) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g1022 ( .A(n_726), .Y(n_1022) );
INVx3_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g846 ( .A(n_737), .Y(n_846) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_739), .A2(n_857), .B1(n_867), .B2(n_875), .C(n_876), .Y(n_856) );
AOI221xp5_ASAP7_75t_L g1049 ( .A1(n_739), .A2(n_875), .B1(n_1050), .B2(n_1055), .C(n_1059), .Y(n_1049) );
AOI33xp33_ASAP7_75t_L g1196 ( .A1(n_739), .A2(n_875), .A3(n_1197), .B1(n_1200), .B2(n_1201), .B3(n_1204), .Y(n_1196) );
NAND3xp33_ASAP7_75t_L g1554 ( .A(n_739), .B(n_1555), .C(n_1557), .Y(n_1554) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g1028 ( .A(n_744), .Y(n_1028) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_747), .Y(n_1009) );
BUFx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g982 ( .A(n_767), .Y(n_982) );
AO22x2_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_890), .B1(n_891), .B2(n_980), .Y(n_767) );
INVx1_ASAP7_75t_L g980 ( .A(n_768), .Y(n_980) );
XNOR2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_824), .Y(n_768) );
INVx1_ASAP7_75t_L g823 ( .A(n_771), .Y(n_823) );
NAND4xp25_ASAP7_75t_L g792 ( .A(n_793), .B(n_803), .C(n_811), .D(n_818), .Y(n_792) );
INVx2_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g808 ( .A(n_798), .Y(n_808) );
INVx1_ASAP7_75t_L g870 ( .A(n_798), .Y(n_870) );
INVx2_ASAP7_75t_L g1155 ( .A(n_798), .Y(n_1155) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx3_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g963 ( .A(n_814), .Y(n_963) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND3x1_ASAP7_75t_L g825 ( .A(n_826), .B(n_842), .C(n_856), .Y(n_825) );
OR2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
INVx2_ASAP7_75t_L g880 ( .A(n_830), .Y(n_880) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
OAI221xp5_ASAP7_75t_L g1110 ( .A1(n_837), .A2(n_879), .B1(n_1111), .B2(n_1112), .C(n_1113), .Y(n_1110) );
INVx2_ASAP7_75t_SL g837 ( .A(n_838), .Y(n_837) );
OAI221xp5_ASAP7_75t_L g886 ( .A1(n_845), .A2(n_848), .B1(n_879), .B2(n_887), .C(n_889), .Y(n_886) );
OR2x2_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
BUFx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g1092 ( .A(n_854), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .B1(n_862), .B2(n_863), .Y(n_858) );
INVx3_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g1086 ( .A1(n_865), .A2(n_873), .B1(n_1087), .B2(n_1088), .Y(n_1086) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
OAI22xp33_ASAP7_75t_SL g1089 ( .A1(n_870), .A2(n_1090), .B1(n_1091), .B2(n_1093), .Y(n_1089) );
OAI221xp5_ASAP7_75t_L g878 ( .A1(n_872), .A2(n_874), .B1(n_879), .B2(n_881), .C(n_883), .Y(n_878) );
OAI22xp5_ASAP7_75t_SL g876 ( .A1(n_877), .A2(n_878), .B1(n_885), .B2(n_886), .Y(n_876) );
OAI22xp5_ASAP7_75t_SL g1059 ( .A1(n_877), .A2(n_885), .B1(n_1060), .B2(n_1063), .Y(n_1059) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g1061 ( .A(n_880), .Y(n_1061) );
INVx2_ASAP7_75t_L g1105 ( .A(n_880), .Y(n_1105) );
OAI221xp5_ASAP7_75t_L g1060 ( .A1(n_881), .A2(n_1052), .B1(n_1054), .B2(n_1061), .C(n_1062), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_881), .A2(n_1061), .B1(n_1064), .B2(n_1065), .C(n_1066), .Y(n_1063) );
BUFx3_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g1027 ( .A(n_884), .Y(n_1027) );
INVx1_ASAP7_75t_L g1031 ( .A(n_885), .Y(n_1031) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVxp67_ASAP7_75t_SL g890 ( .A(n_891), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_938), .B1(n_939), .B2(n_979), .Y(n_891) );
INVx1_ASAP7_75t_L g979 ( .A(n_892), .Y(n_979) );
NAND3xp33_ASAP7_75t_L g905 ( .A(n_906), .B(n_910), .C(n_913), .Y(n_905) );
NAND4xp25_ASAP7_75t_L g915 ( .A(n_916), .B(n_921), .C(n_930), .D(n_935), .Y(n_915) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g978 ( .A(n_940), .Y(n_978) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_960), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g1281 ( .A1(n_977), .A2(n_1282), .B1(n_1283), .B2(n_1288), .Y(n_1281) );
INVxp67_ASAP7_75t_SL g1262 ( .A(n_983), .Y(n_1262) );
AOI22xp5_ASAP7_75t_L g983 ( .A1(n_984), .A2(n_985), .B1(n_1074), .B2(n_1075), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
XNOR2x2_ASAP7_75t_L g986 ( .A(n_987), .B(n_1038), .Y(n_986) );
XNOR2xp5_ASAP7_75t_L g987 ( .A(n_988), .B(n_989), .Y(n_987) );
NAND4xp25_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1017), .C(n_1023), .D(n_1030), .Y(n_1011) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVxp67_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
NAND3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .C(n_1029), .Y(n_1023) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
NAND3xp33_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1032), .C(n_1035), .Y(n_1030) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1037), .Y(n_1214) );
XNOR2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1040), .Y(n_1038) );
NAND3x1_ASAP7_75t_SL g1040 ( .A(n_1041), .B(n_1049), .C(n_1067), .Y(n_1040) );
OAI22xp33_ASAP7_75t_L g1098 ( .A1(n_1053), .A2(n_1099), .B1(n_1100), .B2(n_1101), .Y(n_1098) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
XNOR2xp5_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1169), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1078), .B1(n_1130), .B2(n_1168), .Y(n_1076) );
INVx2_ASAP7_75t_SL g1077 ( .A(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
NAND3xp33_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1114), .C(n_1123), .Y(n_1081) );
NOR2xp33_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1103), .Y(n_1082) );
OAI33xp33_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1086), .A3(n_1089), .B1(n_1094), .B2(n_1098), .B3(n_1102), .Y(n_1083) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_1087), .A2(n_1088), .B1(n_1105), .B2(n_1106), .C(n_1109), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_1091), .A2(n_1095), .B1(n_1096), .B2(n_1097), .Y(n_1094) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1096), .Y(n_1522) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1119), .Y(n_1162) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1130), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
NAND3x1_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1145), .C(n_1150), .Y(n_1132) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1138), .Y(n_1579) );
AND4x1_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1157), .C(n_1160), .D(n_1165), .Y(n_1150) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1171), .B1(n_1219), .B2(n_1220), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1173), .Y(n_1218) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1205), .Y(n_1195) );
HB1xp67_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx2_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
BUFx6f_ASAP7_75t_L g1528 ( .A(n_1213), .Y(n_1528) );
INVx2_ASAP7_75t_SL g1219 ( .A(n_1220), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1242), .Y(n_1234) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx2_ASAP7_75t_SL g1250 ( .A(n_1245), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
OAI221xp5_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1487), .B1(n_1490), .B2(n_1538), .C(n_1543), .Y(n_1263) );
NOR3xp33_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1448), .C(n_1470), .Y(n_1264) );
AOI22xp5_ASAP7_75t_L g1265 ( .A1(n_1266), .A2(n_1343), .B1(n_1410), .B2(n_1422), .Y(n_1265) );
AOI311xp33_ASAP7_75t_L g1266 ( .A1(n_1267), .A2(n_1307), .A3(n_1322), .B(n_1325), .C(n_1338), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
NOR2xp33_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1299), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1269), .B(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
OAI22xp33_ASAP7_75t_L g1345 ( .A1(n_1270), .A2(n_1318), .B1(n_1346), .B2(n_1349), .Y(n_1345) );
NOR2xp33_ASAP7_75t_L g1428 ( .A(n_1270), .B(n_1378), .Y(n_1428) );
OAI21xp33_ASAP7_75t_SL g1435 ( .A1(n_1270), .A2(n_1377), .B(n_1436), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1290), .Y(n_1270) );
INVx2_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1272), .B(n_1303), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1272), .B(n_1290), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1272), .B(n_1329), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g1404 ( .A(n_1272), .B(n_1290), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1272), .B(n_1353), .Y(n_1441) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1273), .B(n_1329), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1273), .B(n_1303), .Y(n_1387) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1274), .Y(n_1359) );
BUFx3_ASAP7_75t_L g1489 ( .A(n_1274), .Y(n_1489) );
AND2x4_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1278), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1275), .B(n_1278), .Y(n_1320) );
HB1xp67_ASAP7_75t_L g1593 ( .A(n_1275), .Y(n_1593) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
AND2x4_ASAP7_75t_L g1280 ( .A(n_1276), .B(n_1278), .Y(n_1280) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1277), .B(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1279), .Y(n_1287) );
INVx2_ASAP7_75t_L g1312 ( .A(n_1280), .Y(n_1312) );
OAI22xp33_ASAP7_75t_L g1304 ( .A1(n_1283), .A2(n_1288), .B1(n_1305), .B2(n_1306), .Y(n_1304) );
OAI22xp33_ASAP7_75t_L g1313 ( .A1(n_1283), .A2(n_1314), .B1(n_1315), .B2(n_1316), .Y(n_1313) );
BUFx3_ASAP7_75t_L g1362 ( .A(n_1283), .Y(n_1362) );
BUFx6f_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1286), .Y(n_1284) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_1285), .B(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1285), .Y(n_1295) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1286), .Y(n_1294) );
HB1xp67_ASAP7_75t_L g1592 ( .A(n_1287), .Y(n_1592) );
HB1xp67_ASAP7_75t_L g1316 ( .A(n_1288), .Y(n_1316) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1288), .Y(n_1365) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1289), .Y(n_1297) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1290), .B(n_1301), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1290), .B(n_1322), .Y(n_1330) );
OR2x2_ASAP7_75t_L g1425 ( .A(n_1290), .B(n_1352), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1290), .B(n_1433), .Y(n_1468) );
BUFx3_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1291), .B(n_1328), .Y(n_1339) );
INVx2_ASAP7_75t_L g1353 ( .A(n_1291), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1374 ( .A(n_1291), .B(n_1375), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1291), .B(n_1372), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1291), .B(n_1387), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1291), .B(n_1302), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1291), .B(n_1352), .Y(n_1453) );
O2A1O1Ixp33_ASAP7_75t_L g1462 ( .A1(n_1291), .A2(n_1463), .B(n_1467), .C(n_1469), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1298), .Y(n_1291) );
AND2x4_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1295), .Y(n_1293) );
AND2x4_ASAP7_75t_L g1296 ( .A(n_1295), .B(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
AOI21xp5_ASAP7_75t_L g1373 ( .A1(n_1301), .A2(n_1374), .B(n_1376), .Y(n_1373) );
AOI32xp33_ASAP7_75t_L g1426 ( .A1(n_1301), .A2(n_1326), .A3(n_1380), .B1(n_1427), .B2(n_1428), .Y(n_1426) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1302), .B(n_1378), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1302), .B(n_1330), .Y(n_1452) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1303), .Y(n_1329) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1303), .Y(n_1352) );
NAND2xp5_ASAP7_75t_L g1389 ( .A(n_1307), .B(n_1390), .Y(n_1389) );
AOI22xp33_ASAP7_75t_SL g1451 ( .A1(n_1307), .A2(n_1408), .B1(n_1452), .B2(n_1453), .Y(n_1451) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1317), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1309), .B(n_1318), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1309), .B(n_1384), .Y(n_1445) );
AND2x4_ASAP7_75t_SL g1461 ( .A(n_1309), .B(n_1317), .Y(n_1461) );
INVx2_ASAP7_75t_SL g1309 ( .A(n_1310), .Y(n_1309) );
INVx2_ASAP7_75t_L g1341 ( .A(n_1310), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1383 ( .A(n_1310), .B(n_1384), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1310), .B(n_1317), .Y(n_1486) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1317), .B(n_1332), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1317), .B(n_1335), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1317), .B(n_1380), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1317), .B(n_1419), .Y(n_1442) );
CKINVDCx6p67_ASAP7_75t_R g1317 ( .A(n_1318), .Y(n_1317) );
CKINVDCx5p33_ASAP7_75t_R g1326 ( .A(n_1318), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1318), .B(n_1335), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1318), .B(n_1370), .Y(n_1369) );
AOI221xp5_ASAP7_75t_L g1477 ( .A1(n_1318), .A2(n_1412), .B1(n_1478), .B2(n_1482), .C(n_1483), .Y(n_1477) );
OR2x6_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1321), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1322), .B(n_1335), .Y(n_1334) );
INVx4_ASAP7_75t_L g1347 ( .A(n_1322), .Y(n_1347) );
INVx3_ASAP7_75t_L g1378 ( .A(n_1322), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1322), .B(n_1372), .Y(n_1436) );
NOR2xp67_ASAP7_75t_SL g1458 ( .A(n_1322), .B(n_1333), .Y(n_1458) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_1322), .B(n_1335), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1322), .B(n_1369), .Y(n_1482) );
AND2x4_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1324), .Y(n_1322) );
OAI21xp33_ASAP7_75t_L g1325 ( .A1(n_1326), .A2(n_1327), .B(n_1331), .Y(n_1325) );
A2O1A1Ixp33_ASAP7_75t_L g1417 ( .A1(n_1326), .A2(n_1384), .B(n_1418), .C(n_1420), .Y(n_1417) );
OAI211xp5_ASAP7_75t_SL g1423 ( .A1(n_1327), .A2(n_1368), .B(n_1424), .C(n_1426), .Y(n_1423) );
OR2x2_ASAP7_75t_L g1471 ( .A(n_1327), .B(n_1384), .Y(n_1471) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1327), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1330), .Y(n_1327) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1328), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1328), .B(n_1347), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1328), .B(n_1427), .Y(n_1450) );
INVxp67_ASAP7_75t_L g1484 ( .A(n_1332), .Y(n_1484) );
NOR2xp33_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1334), .Y(n_1332) );
INVx1_ASAP7_75t_SL g1370 ( .A(n_1335), .Y(n_1370) );
CKINVDCx5p33_ASAP7_75t_R g1380 ( .A(n_1335), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1335), .B(n_1347), .Y(n_1395) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1335), .Y(n_1409) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1335), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1335), .B(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1335), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1337), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1340), .Y(n_1338) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1339), .Y(n_1446) );
OAI21xp33_ASAP7_75t_L g1411 ( .A1(n_1340), .A2(n_1412), .B(n_1413), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1342), .Y(n_1340) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1341), .Y(n_1354) );
INVx2_ASAP7_75t_L g1399 ( .A(n_1341), .Y(n_1399) );
OAI211xp5_ASAP7_75t_SL g1470 ( .A1(n_1341), .A2(n_1471), .B(n_1472), .C(n_1477), .Y(n_1470) );
NOR2xp33_ASAP7_75t_L g1473 ( .A(n_1341), .B(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1342), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1381), .Y(n_1343) );
AOI211xp5_ASAP7_75t_L g1344 ( .A1(n_1345), .A2(n_1354), .B(n_1355), .C(n_1373), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1347), .B(n_1348), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1347), .B(n_1351), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1347), .B(n_1386), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1347), .B(n_1369), .Y(n_1416) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1347), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1347), .B(n_1353), .Y(n_1427) );
AOI22xp5_ASAP7_75t_L g1440 ( .A1(n_1348), .A2(n_1351), .B1(n_1441), .B2(n_1442), .Y(n_1440) );
AOI31xp33_ASAP7_75t_L g1456 ( .A1(n_1349), .A2(n_1374), .A3(n_1434), .B(n_1457), .Y(n_1456) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
NOR2x1_ASAP7_75t_L g1351 ( .A(n_1352), .B(n_1353), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1353), .B(n_1372), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1353), .B(n_1387), .Y(n_1386) );
OR2x2_ASAP7_75t_L g1421 ( .A(n_1353), .B(n_1401), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1354), .B(n_1397), .Y(n_1396) );
OAI21xp33_ASAP7_75t_L g1402 ( .A1(n_1354), .A2(n_1403), .B(n_1405), .Y(n_1402) );
AOI211xp5_ASAP7_75t_L g1422 ( .A1(n_1354), .A2(n_1423), .B(n_1429), .C(n_1439), .Y(n_1422) );
OAI221xp5_ASAP7_75t_L g1448 ( .A1(n_1354), .A2(n_1449), .B1(n_1451), .B2(n_1454), .C(n_1455), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1366), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
BUFx3_ASAP7_75t_L g1438 ( .A(n_1357), .Y(n_1438) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
OAI22xp33_ASAP7_75t_L g1360 ( .A1(n_1361), .A2(n_1362), .B1(n_1363), .B2(n_1364), .Y(n_1360) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
NOR2xp33_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1371), .Y(n_1367) );
OAI21xp33_ASAP7_75t_L g1429 ( .A1(n_1368), .A2(n_1430), .B(n_1432), .Y(n_1429) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1371), .Y(n_1412) );
OR2x2_ASAP7_75t_L g1460 ( .A(n_1371), .B(n_1378), .Y(n_1460) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1372), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1475 ( .A(n_1374), .B(n_1476), .Y(n_1475) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1379), .Y(n_1376) );
OR2x2_ASAP7_75t_L g1424 ( .A(n_1377), .B(n_1425), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1377), .B(n_1386), .Y(n_1431) );
INVx2_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1378), .B(n_1392), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1378), .B(n_1404), .Y(n_1413) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1379), .Y(n_1447) );
INVx3_ASAP7_75t_L g1384 ( .A(n_1380), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_1380), .B(n_1461), .Y(n_1469) );
AOI211xp5_ASAP7_75t_SL g1381 ( .A1(n_1382), .A2(n_1385), .B(n_1388), .C(n_1393), .Y(n_1381) );
AOI221xp5_ASAP7_75t_L g1432 ( .A1(n_1382), .A2(n_1433), .B1(n_1434), .B2(n_1435), .C(n_1437), .Y(n_1432) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1387), .Y(n_1466) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1392), .Y(n_1476) );
OAI21xp5_ASAP7_75t_SL g1393 ( .A1(n_1394), .A2(n_1396), .B(n_1398), .Y(n_1393) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
OAI211xp5_ASAP7_75t_L g1398 ( .A1(n_1399), .A2(n_1400), .B(n_1402), .C(n_1406), .Y(n_1398) );
OAI222xp33_ASAP7_75t_L g1439 ( .A1(n_1399), .A2(n_1440), .B1(n_1443), .B2(n_1445), .C1(n_1446), .C2(n_1447), .Y(n_1439) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVxp33_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1404), .B(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1408), .B(n_1409), .Y(n_1407) );
AND3x1_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1414), .C(n_1417), .Y(n_1410) );
OAI21xp33_ASAP7_75t_L g1472 ( .A1(n_1415), .A2(n_1473), .B(n_1475), .Y(n_1472) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1434), .Y(n_1454) );
INVx2_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
AOI21xp5_ASAP7_75t_L g1483 ( .A1(n_1443), .A2(n_1484), .B(n_1485), .Y(n_1483) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
O2A1O1Ixp33_ASAP7_75t_L g1455 ( .A1(n_1456), .A2(n_1459), .B(n_1461), .C(n_1462), .Y(n_1455) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
NAND2xp5_ASAP7_75t_L g1464 ( .A(n_1465), .B(n_1466), .Y(n_1464) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1481), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
HB1xp67_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1493), .Y(n_1537) );
NAND3xp33_ASAP7_75t_L g1494 ( .A(n_1495), .B(n_1500), .C(n_1503), .Y(n_1494) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
NAND4xp25_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1520), .C(n_1526), .D(n_1531), .Y(n_1516) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
NAND3xp33_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1534), .C(n_1535), .Y(n_1531) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
CKINVDCx5p33_ASAP7_75t_R g1538 ( .A(n_1539), .Y(n_1538) );
BUFx2_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
INVxp33_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1547), .Y(n_1584) );
INVxp33_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
NAND3xp33_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1565), .C(n_1575), .Y(n_1548) );
AND4x1_ASAP7_75t_L g1549 ( .A(n_1550), .B(n_1554), .C(n_1558), .D(n_1561), .Y(n_1549) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
CKINVDCx5p33_ASAP7_75t_R g1586 ( .A(n_1587), .Y(n_1586) );
A2O1A1Ixp33_ASAP7_75t_L g1590 ( .A1(n_1588), .A2(n_1591), .B(n_1593), .C(n_1594), .Y(n_1590) );
HB1xp67_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
endmodule