module fake_jpeg_12292_n_156 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_8),
.B(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_72),
.Y(n_82)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_19),
.B1(n_41),
.B2(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_73),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_0),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_83),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_87),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_62),
.B1(n_54),
.B2(n_46),
.Y(n_81)
);

OAI22x1_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_45),
.B1(n_49),
.B2(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_1),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_62),
.B1(n_64),
.B2(n_54),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_93),
.B1(n_5),
.B2(n_6),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_65),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_95),
.C(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_100),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_80),
.B(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_50),
.B1(n_45),
.B2(n_3),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_10),
.B(n_11),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_2),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_1),
.B(n_2),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_110),
.Y(n_120)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_114),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_4),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_4),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_116),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_7),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_7),
.C(n_8),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_93),
.C(n_24),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_129),
.B1(n_124),
.B2(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_12),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_13),
.Y(n_127)
);

NOR4xp25_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_128),
.C(n_23),
.D(n_26),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_14),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_138),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_42),
.C(n_25),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_141),
.B1(n_121),
.B2(n_130),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_118),
.B1(n_115),
.B2(n_129),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_146),
.A2(n_27),
.B1(n_30),
.B2(n_32),
.Y(n_151)
);

OAI321xp33_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_131),
.A3(n_133),
.B1(n_137),
.B2(n_138),
.C(n_111),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_147),
.A2(n_135),
.B1(n_133),
.B2(n_142),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_149),
.A2(n_150),
.B(n_151),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_143),
.B(n_144),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_143),
.B(n_145),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_149),
.Y(n_156)
);


endmodule