module fake_netlist_6_1845_n_1915 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1915);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1915;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_474;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_141),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_78),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_25),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_121),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_51),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_24),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_143),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_83),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_28),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_90),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_144),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_62),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_50),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_61),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_126),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_80),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_124),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_50),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_24),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_73),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_21),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_9),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_21),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_64),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_116),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_74),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_109),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_47),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_6),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_47),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_26),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_32),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_1),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_2),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_101),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_55),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_93),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_104),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_96),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_167),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_118),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_75),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_18),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_164),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_2),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_95),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_51),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_140),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_34),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_130),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_85),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_23),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_9),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_94),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_86),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_55),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_41),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_7),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_105),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_60),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_91),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_44),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_15),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_180),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_35),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_39),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_99),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_179),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_66),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_166),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_12),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_112),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_171),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_3),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_67),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_89),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_15),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_63),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_64),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_67),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_136),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_153),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_170),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_165),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_84),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_113),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_31),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_154),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_23),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_150),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_128),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_56),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_127),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_4),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_119),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_107),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_12),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_30),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_17),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_45),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_17),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_148),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_1),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_147),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_40),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_108),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_181),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_133),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_20),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_33),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_71),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_97),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_32),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_172),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_123),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_102),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_82),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_61),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_139),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_146),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_62),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_5),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_56),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_27),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_92),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_22),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_182),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_79),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_117),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_114),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_35),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_178),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_34),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_25),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_168),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_65),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_26),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_87),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_156),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_68),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_19),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_98),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_110),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_132),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_7),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_0),
.Y(n_342)
);

INVx4_ASAP7_75t_R g343 ( 
.A(n_77),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_60),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_58),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_30),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_70),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_40),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_14),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_149),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_29),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_11),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_169),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_145),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_38),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_28),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_44),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_19),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_131),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_48),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_76),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_52),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_53),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_161),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_183),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_184),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_186),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_188),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_326),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_191),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_207),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_298),
.B(n_255),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_207),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_196),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_192),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_227),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_189),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_195),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_198),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_207),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_196),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_203),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_207),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_207),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_204),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_249),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_207),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_290),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_188),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_205),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_317),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_208),
.B(n_0),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_215),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_208),
.B(n_243),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_279),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_216),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_317),
.B(n_3),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_217),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_249),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_243),
.B(n_4),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_317),
.B(n_5),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_290),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_227),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_236),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_189),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_226),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_290),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_290),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_290),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_229),
.Y(n_410)
);

INVx4_ASAP7_75t_R g411 ( 
.A(n_279),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_312),
.B(n_6),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_263),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_286),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_290),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_232),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_225),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_194),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_260),
.B(n_8),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_234),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_258),
.B(n_8),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_286),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_236),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_233),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_225),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_225),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_237),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_239),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_278),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_312),
.B(n_10),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_185),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_241),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_225),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_278),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_225),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_258),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_245),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_319),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_228),
.B(n_10),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_319),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_254),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_260),
.B(n_307),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_256),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_259),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_194),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_L g446 ( 
.A(n_200),
.B(n_11),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_262),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_268),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_190),
.B(n_13),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_200),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_213),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_280),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_263),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_190),
.B(n_14),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_263),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_282),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_417),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_417),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_394),
.B(n_284),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_425),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_371),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_371),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_413),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_373),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_281),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_391),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_372),
.B(n_365),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_376),
.A2(n_211),
.B1(n_266),
.B2(n_336),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_373),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_L g475 ( 
.A(n_430),
.B(n_187),
.Y(n_475)
);

AND2x2_ASAP7_75t_SL g476 ( 
.A(n_430),
.B(n_228),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_401),
.B(n_364),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_366),
.B(n_323),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_392),
.B(n_287),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_413),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_433),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_453),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_433),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_400),
.B(n_289),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_401),
.B(n_364),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_435),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_380),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_435),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_383),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_383),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_453),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_367),
.B(n_370),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_412),
.B(n_291),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_384),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_384),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_403),
.B(n_342),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_387),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_455),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_387),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_388),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_402),
.B(n_292),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_419),
.B(n_230),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_407),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_397),
.B(n_335),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_407),
.B(n_300),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_408),
.B(n_302),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_408),
.B(n_308),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_409),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_455),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_409),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_415),
.B(n_310),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_375),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_415),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_445),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_445),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_455),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_450),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_450),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_451),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_436),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_451),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_436),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_438),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_438),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_440),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_440),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_439),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_439),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_397),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_368),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_429),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_368),
.B(n_313),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_378),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_469),
.B(n_379),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_519),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_530),
.B(n_368),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_471),
.B(n_382),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_515),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_507),
.B(n_385),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_465),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_530),
.B(n_390),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_476),
.A2(n_419),
.B1(n_454),
.B2(n_449),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_507),
.B(n_393),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_396),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_459),
.B(n_398),
.Y(n_548)
);

OAI22xp33_ASAP7_75t_L g549 ( 
.A1(n_531),
.A2(n_376),
.B1(n_404),
.B2(n_403),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_464),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_519),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_533),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_533),
.B(n_442),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_465),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_406),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_532),
.B(n_410),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_532),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_464),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_519),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_462),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_476),
.B(n_416),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_519),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_465),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_532),
.B(n_420),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_532),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_496),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_496),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_533),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_462),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_493),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_459),
.B(n_428),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_464),
.Y(n_572)
);

NAND3xp33_ASAP7_75t_L g573 ( 
.A(n_476),
.B(n_446),
.C(n_421),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_532),
.B(n_437),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_465),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_498),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_464),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_472),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_478),
.B(n_441),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_L g580 ( 
.A1(n_479),
.A2(n_404),
.B1(n_423),
.B2(n_327),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_470),
.B(n_443),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_470),
.B(n_447),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_504),
.A2(n_446),
.B1(n_421),
.B2(n_434),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_498),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_479),
.B(n_452),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_485),
.B(n_432),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_472),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_483),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_470),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_485),
.B(n_424),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_494),
.B(n_389),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_494),
.B(n_444),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_501),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_477),
.B(n_389),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_483),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_501),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_535),
.B(n_427),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_504),
.A2(n_351),
.B1(n_307),
.B2(n_288),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_506),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_506),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_477),
.B(n_389),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_535),
.B(n_448),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_R g603 ( 
.A(n_477),
.B(n_197),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_511),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_504),
.B(n_395),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_511),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_477),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_483),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_513),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_465),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_534),
.B(n_423),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_504),
.A2(n_351),
.B1(n_214),
.B2(n_219),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_534),
.B(n_456),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_486),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_533),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_483),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_504),
.A2(n_288),
.B1(n_213),
.B2(n_214),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_465),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_513),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_492),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_492),
.Y(n_622)
);

AND2x6_ASAP7_75t_L g623 ( 
.A(n_486),
.B(n_230),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_516),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_517),
.B(n_395),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_497),
.B(n_533),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_492),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_492),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_486),
.B(n_395),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_486),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_533),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_516),
.Y(n_632)
);

INVx4_ASAP7_75t_SL g633 ( 
.A(n_465),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_533),
.B(n_193),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_480),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_503),
.B(n_508),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_462),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_463),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_486),
.B(n_374),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_480),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_503),
.B(n_381),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_480),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_480),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_463),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_463),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_467),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_480),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_517),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_508),
.B(n_386),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_467),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_509),
.B(n_399),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_518),
.B(n_405),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_475),
.A2(n_295),
.B1(n_294),
.B2(n_285),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_480),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_509),
.B(n_324),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_480),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_482),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_457),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_467),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_510),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_510),
.B(n_414),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_457),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_482),
.B(n_193),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_514),
.B(n_325),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_514),
.B(n_328),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_L g666 ( 
.A1(n_518),
.A2(n_253),
.B1(n_363),
.B2(n_360),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_520),
.B(n_422),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_520),
.B(n_369),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_521),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_473),
.Y(n_670)
);

BUFx4f_ASAP7_75t_L g671 ( 
.A(n_482),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_521),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_522),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_482),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_482),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_522),
.Y(n_676)
);

INVxp33_ASAP7_75t_SL g677 ( 
.A(n_524),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_524),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_525),
.B(n_199),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_527),
.B(n_331),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_525),
.B(n_377),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_473),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_482),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_482),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_526),
.B(n_405),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_458),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_526),
.B(n_418),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_499),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_636),
.A2(n_219),
.B(n_220),
.C(n_242),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_566),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_605),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_660),
.B(n_548),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_605),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_544),
.B(n_201),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_566),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_557),
.B(n_499),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_669),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_660),
.B(n_499),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_571),
.B(n_499),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_567),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_542),
.B(n_499),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_591),
.B(n_499),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_539),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_669),
.Y(n_704)
);

INVxp33_ASAP7_75t_L g705 ( 
.A(n_614),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_565),
.B(n_499),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_565),
.B(n_512),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_541),
.Y(n_708)
);

NOR2x1p5_ASAP7_75t_L g709 ( 
.A(n_547),
.B(n_206),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_555),
.B(n_512),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_557),
.B(n_512),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_557),
.B(n_512),
.Y(n_712)
);

AO22x1_ASAP7_75t_L g713 ( 
.A1(n_586),
.A2(n_299),
.B1(n_362),
.B2(n_248),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_539),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_556),
.B(n_564),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_561),
.A2(n_334),
.B1(n_361),
.B2(n_339),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_567),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_576),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_557),
.B(n_512),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_673),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_589),
.B(n_512),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_585),
.B(n_512),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_L g723 ( 
.A(n_570),
.B(n_573),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_589),
.B(n_458),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_677),
.B(n_210),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_668),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_608),
.B(n_263),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_608),
.B(n_263),
.Y(n_728)
);

NAND2x1p5_ASAP7_75t_L g729 ( 
.A(n_553),
.B(n_199),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_573),
.B(n_523),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_673),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_546),
.B(n_218),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_625),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_612),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_625),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_538),
.B(n_460),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_681),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_538),
.B(n_460),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_551),
.B(n_461),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_576),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_551),
.B(n_461),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_559),
.B(n_466),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_559),
.B(n_466),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_607),
.B(n_263),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_584),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_607),
.B(n_263),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_562),
.B(n_579),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_678),
.Y(n_748)
);

INVx8_ASAP7_75t_L g749 ( 
.A(n_623),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_681),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_545),
.A2(n_562),
.B(n_592),
.C(n_648),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_652),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_607),
.B(n_263),
.Y(n_753)
);

BUFx8_ASAP7_75t_L g754 ( 
.A(n_652),
.Y(n_754)
);

AND2x6_ASAP7_75t_L g755 ( 
.A(n_634),
.B(n_202),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_553),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_553),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_581),
.B(n_221),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_553),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_658),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_602),
.B(n_523),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_687),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_667),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_658),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_655),
.B(n_664),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_665),
.B(n_468),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_584),
.Y(n_767)
);

NOR2xp67_ASAP7_75t_L g768 ( 
.A(n_641),
.B(n_523),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_583),
.B(n_223),
.C(n_222),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_582),
.B(n_238),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_594),
.B(n_468),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_601),
.B(n_481),
.Y(n_772)
);

NAND2x1_ASAP7_75t_L g773 ( 
.A(n_623),
.B(n_343),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_676),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_629),
.B(n_481),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_672),
.B(n_484),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_685),
.B(n_528),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_593),
.B(n_484),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_662),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_662),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_578),
.B(n_240),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_593),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_686),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_596),
.B(n_487),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_607),
.B(n_263),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_596),
.B(n_487),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_686),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_615),
.B(n_350),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_599),
.B(n_600),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_599),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_676),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_600),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_676),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_604),
.B(n_489),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_604),
.B(n_489),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_649),
.B(n_246),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_603),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_606),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_676),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_SL g800 ( 
.A(n_587),
.B(n_257),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_630),
.A2(n_353),
.B1(n_354),
.B2(n_202),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_537),
.B(n_251),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_615),
.B(n_209),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_606),
.B(n_523),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_540),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_580),
.B(n_252),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_626),
.A2(n_304),
.B1(n_271),
.B2(n_359),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_685),
.B(n_529),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_651),
.B(n_264),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_590),
.A2(n_304),
.B1(n_267),
.B2(n_359),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_610),
.B(n_527),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_661),
.B(n_269),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_687),
.B(n_529),
.Y(n_813)
);

INVx8_ASAP7_75t_L g814 ( 
.A(n_623),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_610),
.B(n_527),
.Y(n_815)
);

O2A1O1Ixp5_ASAP7_75t_L g816 ( 
.A1(n_620),
.A2(n_267),
.B(n_209),
.C(n_212),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_620),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_653),
.A2(n_250),
.B1(n_247),
.B2(n_244),
.Y(n_818)
);

OAI21xp33_ASAP7_75t_L g819 ( 
.A1(n_618),
.A2(n_598),
.B(n_613),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_624),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_624),
.B(n_632),
.Y(n_821)
);

OAI22xp33_ASAP7_75t_L g822 ( 
.A1(n_679),
.A2(n_265),
.B1(n_303),
.B2(n_250),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_597),
.B(n_639),
.C(n_574),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_632),
.A2(n_311),
.B(n_224),
.C(n_231),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_536),
.B(n_527),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_549),
.B(n_666),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_679),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_634),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_637),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_543),
.B(n_527),
.Y(n_830)
);

OAI221xp5_ASAP7_75t_L g831 ( 
.A1(n_679),
.A2(n_295),
.B1(n_362),
.B2(n_355),
.C(n_345),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_634),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_615),
.B(n_212),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_679),
.B(n_270),
.C(n_358),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_SL g835 ( 
.A(n_554),
.B(n_224),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_623),
.A2(n_265),
.B1(n_340),
.B2(n_338),
.Y(n_836)
);

CKINVDCx11_ASAP7_75t_R g837 ( 
.A(n_679),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_543),
.B(n_527),
.Y(n_838)
);

AOI221xp5_ASAP7_75t_L g839 ( 
.A1(n_634),
.A2(n_273),
.B1(n_261),
.B2(n_346),
.C(n_355),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_554),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_554),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_623),
.A2(n_248),
.B1(n_345),
.B2(n_220),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_543),
.B(n_527),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_637),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_543),
.B(n_274),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_615),
.B(n_231),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_611),
.A2(n_247),
.B(n_340),
.C(n_338),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_552),
.B(n_528),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_637),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_611),
.B(n_619),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_638),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_560),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_L g853 ( 
.A(n_623),
.B(n_235),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_554),
.B(n_235),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_611),
.B(n_244),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_560),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_611),
.B(n_271),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_638),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_619),
.B(n_276),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_680),
.B(n_275),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_737),
.B(n_342),
.Y(n_861)
);

INVx6_ASAP7_75t_L g862 ( 
.A(n_754),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_747),
.B(n_623),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_715),
.A2(n_671),
.B(n_631),
.Y(n_864)
);

OAI21xp33_ASAP7_75t_L g865 ( 
.A1(n_796),
.A2(n_293),
.B(n_283),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_692),
.B(n_619),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_SL g867 ( 
.A(n_708),
.B(n_342),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_765),
.B(n_619),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_693),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_751),
.A2(n_671),
.B1(n_657),
.B2(n_643),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_768),
.B(n_640),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_690),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_825),
.A2(n_671),
.B(n_635),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_710),
.A2(n_671),
.B(n_635),
.Y(n_874)
);

NOR2x1p5_ASAP7_75t_L g875 ( 
.A(n_797),
.B(n_296),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_699),
.A2(n_635),
.B(n_575),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_723),
.B(n_554),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_701),
.A2(n_635),
.B(n_575),
.Y(n_878)
);

O2A1O1Ixp5_ASAP7_75t_L g879 ( 
.A1(n_766),
.A2(n_650),
.B(n_644),
.C(n_569),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_750),
.B(n_342),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_823),
.A2(n_643),
.B1(n_654),
.B2(n_656),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_762),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_726),
.B(n_705),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_690),
.Y(n_884)
);

NOR2xp67_ASAP7_75t_L g885 ( 
.A(n_763),
.B(n_550),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_730),
.A2(n_702),
.B(n_722),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_689),
.A2(n_276),
.B(n_321),
.C(n_303),
.Y(n_887)
);

NOR2x2_ASAP7_75t_L g888 ( 
.A(n_839),
.B(n_800),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_754),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_689),
.A2(n_321),
.B(n_277),
.C(n_316),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_694),
.B(n_640),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_693),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_694),
.B(n_640),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_696),
.A2(n_642),
.B(n_575),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_752),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_749),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_826),
.A2(n_320),
.B(n_333),
.C(n_322),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_695),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_721),
.A2(n_647),
.B(n_640),
.Y(n_899)
);

AOI21x1_ASAP7_75t_L g900 ( 
.A1(n_696),
.A2(n_558),
.B(n_550),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_774),
.A2(n_656),
.B1(n_654),
.B2(n_643),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_761),
.B(n_554),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_796),
.B(n_647),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_703),
.B(n_647),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_714),
.B(n_647),
.Y(n_905)
);

AO21x1_ASAP7_75t_L g906 ( 
.A1(n_826),
.A2(n_311),
.B(n_277),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_697),
.B(n_704),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_L g908 ( 
.A(n_725),
.B(n_550),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_748),
.B(n_684),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_720),
.B(n_684),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_848),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_711),
.A2(n_688),
.B(n_575),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_711),
.A2(n_688),
.B(n_642),
.Y(n_913)
);

OAI21xp33_ASAP7_75t_L g914 ( 
.A1(n_806),
.A2(n_329),
.B(n_356),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_731),
.B(n_760),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_749),
.Y(n_916)
);

AOI21x1_ASAP7_75t_L g917 ( 
.A1(n_712),
.A2(n_595),
.B(n_558),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_813),
.Y(n_918)
);

INVx6_ASAP7_75t_L g919 ( 
.A(n_808),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_818),
.A2(n_315),
.B(n_316),
.C(n_645),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_764),
.B(n_779),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_712),
.A2(n_688),
.B(n_642),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_719),
.A2(n_688),
.B(n_642),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_721),
.A2(n_684),
.B(n_683),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_774),
.A2(n_654),
.B1(n_657),
.B2(n_656),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_698),
.A2(n_757),
.B(n_756),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_791),
.B(n_563),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_780),
.B(n_684),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_725),
.B(n_734),
.Y(n_929)
);

NOR2xp67_ASAP7_75t_L g930 ( 
.A(n_716),
.B(n_558),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_783),
.B(n_657),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_700),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_700),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_791),
.B(n_563),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_719),
.A2(n_683),
.B(n_552),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_819),
.A2(n_301),
.B(n_299),
.C(n_294),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_787),
.B(n_563),
.Y(n_937)
);

AOI21x1_ASAP7_75t_L g938 ( 
.A1(n_744),
.A2(n_621),
.B(n_617),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_759),
.A2(n_683),
.B(n_577),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_790),
.B(n_563),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_841),
.A2(n_707),
.B(n_706),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_717),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_799),
.A2(n_552),
.B1(n_568),
.B2(n_616),
.Y(n_943)
);

CKINVDCx8_ASAP7_75t_R g944 ( 
.A(n_805),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_781),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_799),
.B(n_563),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_808),
.B(n_568),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_744),
.A2(n_621),
.B(n_617),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_840),
.A2(n_683),
.B(n_568),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_840),
.A2(n_773),
.B(n_772),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_777),
.B(n_297),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_771),
.A2(n_616),
.B(n_563),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_SL g953 ( 
.A(n_793),
.B(n_305),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_775),
.A2(n_616),
.B(n_675),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_727),
.A2(n_609),
.B(n_572),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_776),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_793),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_850),
.A2(n_674),
.B(n_675),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_749),
.A2(n_674),
.B(n_675),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_814),
.A2(n_674),
.B(n_675),
.Y(n_960)
);

NOR2x1_ASAP7_75t_L g961 ( 
.A(n_709),
.B(n_315),
.Y(n_961)
);

AOI21x1_ASAP7_75t_L g962 ( 
.A1(n_746),
.A2(n_609),
.B(n_588),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_792),
.B(n_572),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_814),
.A2(n_674),
.B(n_675),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_813),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_828),
.A2(n_577),
.B1(n_572),
.B2(n_588),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_814),
.A2(n_674),
.B(n_675),
.Y(n_967)
);

AND2x2_ASAP7_75t_SL g968 ( 
.A(n_842),
.B(n_242),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_803),
.A2(n_846),
.B(n_833),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_717),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_798),
.B(n_577),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_848),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_718),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_718),
.B(n_633),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_740),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_740),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_810),
.A2(n_569),
.B(n_670),
.C(n_659),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_745),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_755),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_727),
.A2(n_595),
.B(n_609),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_745),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_803),
.A2(n_674),
.B(n_595),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_806),
.A2(n_272),
.B(n_285),
.C(n_301),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_767),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_746),
.A2(n_785),
.B(n_753),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_767),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_782),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_817),
.B(n_588),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_820),
.B(n_617),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_755),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_691),
.B(n_732),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_833),
.A2(n_622),
.B(n_627),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_831),
.A2(n_645),
.B(n_670),
.C(n_644),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_782),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_728),
.A2(n_622),
.B(n_627),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_789),
.B(n_621),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_733),
.A2(n_646),
.B(n_650),
.C(n_659),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_732),
.B(n_622),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_821),
.B(n_627),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_829),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_829),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_832),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_735),
.B(n_306),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_844),
.Y(n_1004)
);

AOI21xp33_ASAP7_75t_L g1005 ( 
.A1(n_812),
.A2(n_314),
.B(n_309),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_849),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_849),
.Y(n_1007)
);

AOI21xp33_ASAP7_75t_L g1008 ( 
.A1(n_812),
.A2(n_341),
.B(n_318),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_724),
.B(n_628),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_809),
.B(n_758),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_728),
.A2(n_628),
.B(n_638),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_851),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_846),
.A2(n_628),
.B(n_646),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_804),
.A2(n_682),
.B(n_663),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_802),
.A2(n_272),
.B(n_320),
.C(n_322),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_758),
.B(n_330),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_753),
.A2(n_785),
.B(n_738),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_802),
.A2(n_663),
.B1(n_682),
.B2(n_633),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_770),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_736),
.A2(n_682),
.B(n_633),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_827),
.B(n_633),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_739),
.A2(n_633),
.B(n_473),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_845),
.B(n_663),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_858),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_741),
.A2(n_743),
.B(n_742),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_729),
.A2(n_332),
.B1(n_344),
.B2(n_347),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_770),
.A2(n_333),
.B(n_337),
.C(n_348),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_729),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_858),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_842),
.A2(n_349),
.B1(n_352),
.B2(n_357),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_852),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_853),
.A2(n_491),
.B(n_505),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_788),
.A2(n_491),
.B1(n_505),
.B2(n_502),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_822),
.A2(n_491),
.B(n_505),
.C(n_502),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_830),
.A2(n_490),
.B(n_502),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_845),
.B(n_663),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_755),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_838),
.A2(n_500),
.B(n_495),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_856),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_834),
.A2(n_500),
.B(n_495),
.C(n_490),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_778),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_784),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_755),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_843),
.A2(n_500),
.B(n_495),
.Y(n_1044)
);

OAI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_801),
.A2(n_490),
.B(n_488),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_811),
.A2(n_663),
.B(n_488),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_786),
.B(n_663),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_794),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_837),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_788),
.A2(n_488),
.B(n_474),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_755),
.A2(n_663),
.B1(n_474),
.B2(n_411),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1025),
.A2(n_815),
.B(n_854),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_886),
.A2(n_854),
.B(n_795),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_1016),
.A2(n_807),
.B(n_860),
.C(n_824),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1041),
.B(n_713),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_895),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1042),
.B(n_769),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_968),
.A2(n_857),
.B1(n_855),
.B2(n_859),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_1019),
.B(n_1010),
.Y(n_1059)
);

BUFx2_ASAP7_75t_SL g1060 ( 
.A(n_889),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1048),
.B(n_836),
.Y(n_1061)
);

BUFx2_ASAP7_75t_SL g1062 ( 
.A(n_944),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_956),
.B(n_816),
.Y(n_1063)
);

CKINVDCx10_ASAP7_75t_R g1064 ( 
.A(n_862),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_956),
.B(n_847),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_933),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_1016),
.A2(n_474),
.B(n_411),
.C(n_835),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_864),
.A2(n_162),
.B(n_160),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_933),
.Y(n_1069)
);

AO22x1_ASAP7_75t_L g1070 ( 
.A1(n_1010),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_987),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_945),
.B(n_16),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_862),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_883),
.B(n_951),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_SL g1075 ( 
.A(n_883),
.B(n_1027),
.C(n_983),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_987),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_1019),
.B(n_157),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_984),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_991),
.B(n_22),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_896),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_868),
.A2(n_155),
.B(n_152),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_991),
.B(n_929),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_892),
.Y(n_1083)
);

OA22x2_ASAP7_75t_L g1084 ( 
.A1(n_914),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_921),
.B(n_909),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_872),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_863),
.A2(n_151),
.B(n_138),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_895),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_896),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_1021),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1017),
.A2(n_939),
.B(n_878),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_891),
.A2(n_135),
.B(n_129),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_903),
.A2(n_125),
.B1(n_122),
.B2(n_120),
.Y(n_1093)
);

INVx3_ASAP7_75t_SL g1094 ( 
.A(n_862),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_869),
.B(n_115),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_893),
.A2(n_111),
.B(n_103),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_884),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_909),
.B(n_33),
.Y(n_1098)
);

INVx5_ASAP7_75t_L g1099 ( 
.A(n_896),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_L g1100 ( 
.A(n_1005),
.B(n_36),
.C(n_37),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_L g1101 ( 
.A1(n_927),
.A2(n_100),
.B(n_88),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_892),
.B(n_36),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1008),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_903),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_1104)
);

OAI22x1_ASAP7_75t_L g1105 ( 
.A1(n_888),
.A2(n_875),
.B1(n_961),
.B2(n_882),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_919),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_869),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_873),
.A2(n_72),
.B(n_48),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_869),
.B(n_46),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_L g1110 ( 
.A1(n_867),
.A2(n_46),
.B(n_49),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_915),
.B(n_49),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_938),
.A2(n_52),
.B(n_53),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_876),
.A2(n_54),
.B(n_57),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_984),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_R g1115 ( 
.A(n_1049),
.B(n_54),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_998),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_882),
.B(n_59),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_998),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1004),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_965),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1004),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1007),
.Y(n_1122)
);

NAND2x1_ASAP7_75t_L g1123 ( 
.A(n_896),
.B(n_68),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_965),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_969),
.A2(n_69),
.B(n_70),
.C(n_71),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_869),
.B(n_69),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_902),
.A2(n_72),
.B(n_874),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_907),
.B(n_865),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1007),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1028),
.A2(n_911),
.B1(n_972),
.B2(n_1002),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_898),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_942),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_918),
.B(n_919),
.Y(n_1133)
);

CKINVDCx16_ASAP7_75t_R g1134 ( 
.A(n_953),
.Y(n_1134)
);

OAI22x1_ASAP7_75t_L g1135 ( 
.A1(n_957),
.A2(n_861),
.B1(n_880),
.B2(n_1028),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_970),
.Y(n_1136)
);

NOR3xp33_ASAP7_75t_L g1137 ( 
.A(n_1027),
.B(n_1026),
.C(n_983),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_919),
.Y(n_1138)
);

AOI21x1_ASAP7_75t_L g1139 ( 
.A1(n_927),
.A2(n_946),
.B(n_934),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1000),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_926),
.A2(n_908),
.B(n_885),
.C(n_930),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1021),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_SL g1143 ( 
.A1(n_1023),
.A2(n_1036),
.B(n_1014),
.C(n_1020),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_957),
.Y(n_1144)
);

NOR2x1_ASAP7_75t_SL g1145 ( 
.A(n_916),
.B(n_979),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_SL g1146 ( 
.A1(n_1015),
.A2(n_877),
.B(n_974),
.C(n_897),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_897),
.A2(n_1015),
.B(n_936),
.C(n_1030),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_902),
.A2(n_871),
.B(n_950),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_916),
.B(n_911),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1003),
.B(n_947),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_936),
.A2(n_906),
.B(n_866),
.C(n_877),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_972),
.B(n_1037),
.Y(n_1152)
);

INVxp67_ASAP7_75t_L g1153 ( 
.A(n_1031),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_975),
.A2(n_986),
.B1(n_994),
.B2(n_981),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_941),
.A2(n_934),
.B(n_946),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1000),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_916),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_976),
.B(n_978),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_SL g1159 ( 
.A(n_1037),
.B(n_968),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_894),
.A2(n_922),
.B(n_913),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_932),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_973),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1039),
.B(n_1001),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1040),
.A2(n_890),
.B(n_887),
.C(n_870),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_916),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_996),
.B(n_999),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_979),
.B(n_990),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_904),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1009),
.B(n_1006),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_905),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1012),
.B(n_1024),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1047),
.A2(n_1043),
.B(n_997),
.C(n_1045),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1043),
.A2(n_992),
.B(n_1013),
.C(n_952),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1040),
.A2(n_931),
.B(n_920),
.C(n_928),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_910),
.A2(n_940),
.B(n_937),
.C(n_963),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1029),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_971),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_977),
.A2(n_1018),
.B(n_993),
.C(n_1050),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_988),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_989),
.B(n_985),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_881),
.A2(n_966),
.B(n_974),
.C(n_1034),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_979),
.B(n_990),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1051),
.A2(n_979),
.B1(n_990),
.B2(n_924),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1033),
.A2(n_879),
.B(n_1046),
.C(n_925),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_912),
.A2(n_923),
.B(n_949),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_990),
.A2(n_943),
.B1(n_901),
.B2(n_899),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_935),
.A2(n_954),
.B(n_967),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_879),
.A2(n_980),
.B(n_955),
.C(n_995),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_L g1189 ( 
.A(n_948),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1035),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1011),
.B(n_982),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1022),
.A2(n_1032),
.B(n_1038),
.C(n_1044),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_900),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_962),
.B(n_917),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_R g1195 ( 
.A(n_959),
.B(n_960),
.Y(n_1195)
);

O2A1O1Ixp5_ASAP7_75t_L g1196 ( 
.A1(n_958),
.A2(n_1016),
.B(n_903),
.C(n_715),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_964),
.A2(n_1010),
.B(n_1016),
.C(n_796),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_933),
.Y(n_1198)
);

NOR3xp33_ASAP7_75t_L g1199 ( 
.A(n_1016),
.B(n_1010),
.C(n_726),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1025),
.A2(n_557),
.B(n_715),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_896),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1025),
.A2(n_557),
.B(n_715),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1025),
.A2(n_557),
.B(n_715),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_933),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_956),
.B(n_737),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1010),
.A2(n_1016),
.B(n_796),
.C(n_991),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1016),
.A2(n_1010),
.B(n_1027),
.C(n_826),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_933),
.Y(n_1208)
);

INVx6_ASAP7_75t_L g1209 ( 
.A(n_957),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_933),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1025),
.A2(n_557),
.B(n_715),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1025),
.A2(n_557),
.B(n_715),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1041),
.B(n_692),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1094),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1062),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1200),
.A2(n_1203),
.B(n_1202),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_1206),
.A2(n_1188),
.A3(n_1091),
.B(n_1178),
.Y(n_1217)
);

AO21x2_ASAP7_75t_L g1218 ( 
.A1(n_1197),
.A2(n_1148),
.B(n_1053),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1211),
.A2(n_1212),
.B(n_1166),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1207),
.A2(n_1196),
.B(n_1151),
.Y(n_1220)
);

O2A1O1Ixp5_ASAP7_75t_SL g1221 ( 
.A1(n_1077),
.A2(n_1059),
.B(n_1104),
.C(n_1116),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1176),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1196),
.A2(n_1052),
.B(n_1155),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1213),
.B(n_1199),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1192),
.A2(n_1193),
.B(n_1139),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1186),
.A2(n_1180),
.A3(n_1173),
.B(n_1141),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1083),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1194),
.A2(n_1191),
.B(n_1183),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1143),
.A2(n_1184),
.B(n_1085),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1161),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1112),
.A2(n_1127),
.B(n_1181),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1143),
.A2(n_1180),
.B(n_1054),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1154),
.A2(n_1059),
.B(n_1098),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1074),
.B(n_1205),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1199),
.A2(n_1106),
.B(n_1110),
.Y(n_1235)
);

NAND3x1_ASAP7_75t_L g1236 ( 
.A(n_1079),
.B(n_1117),
.C(n_1082),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1150),
.B(n_1134),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1172),
.A2(n_1175),
.B(n_1159),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1164),
.A2(n_1067),
.B(n_1189),
.Y(n_1239)
);

AOI221x1_ASAP7_75t_L g1240 ( 
.A1(n_1137),
.A2(n_1108),
.B1(n_1125),
.B2(n_1113),
.C(n_1103),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1066),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1161),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1174),
.A2(n_1101),
.B(n_1068),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1167),
.A2(n_1087),
.B(n_1152),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1061),
.A2(n_1075),
.B1(n_1055),
.B2(n_1147),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1189),
.A2(n_1128),
.B(n_1169),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1144),
.B(n_1209),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_SL g1248 ( 
.A1(n_1077),
.A2(n_1167),
.B(n_1182),
.C(n_1095),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1128),
.A2(n_1058),
.B(n_1057),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1177),
.B(n_1179),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1080),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_SL g1252 ( 
.A1(n_1100),
.A2(n_1137),
.B(n_1118),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1056),
.B(n_1088),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1162),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1152),
.A2(n_1171),
.B(n_1076),
.Y(n_1255)
);

AO21x2_ASAP7_75t_L g1256 ( 
.A1(n_1146),
.A2(n_1195),
.B(n_1075),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1158),
.A2(n_1135),
.A3(n_1130),
.B(n_1092),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1158),
.A2(n_1096),
.A3(n_1093),
.B(n_1111),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1058),
.A2(n_1190),
.B(n_1179),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1064),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1094),
.Y(n_1261)
);

INVx3_ASAP7_75t_SL g1262 ( 
.A(n_1138),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1105),
.A2(n_1084),
.B1(n_1126),
.B2(n_1109),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1073),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1120),
.B(n_1124),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1065),
.A2(n_1081),
.B(n_1145),
.Y(n_1266)
);

BUFx12f_ASAP7_75t_L g1267 ( 
.A(n_1102),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1071),
.A2(n_1210),
.A3(n_1208),
.B(n_1204),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1102),
.B(n_1170),
.Y(n_1269)
);

NOR2xp67_ASAP7_75t_L g1270 ( 
.A(n_1056),
.B(n_1088),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1168),
.B(n_1162),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1117),
.A2(n_1072),
.B(n_1153),
.C(n_1168),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1107),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1063),
.A2(n_1131),
.B(n_1132),
.Y(n_1274)
);

NAND3xp33_ASAP7_75t_SL g1275 ( 
.A(n_1115),
.B(n_1123),
.C(n_1133),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1140),
.A2(n_1156),
.B(n_1069),
.Y(n_1276)
);

INVx4_ASAP7_75t_L g1277 ( 
.A(n_1099),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1209),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1107),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1153),
.A2(n_1133),
.B(n_1136),
.C(n_1097),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1163),
.B(n_1198),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1086),
.A2(n_1084),
.B1(n_1090),
.B2(n_1142),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1119),
.A2(n_1121),
.B(n_1129),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1122),
.A2(n_1114),
.A3(n_1078),
.B(n_1165),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1099),
.A2(n_1195),
.B(n_1070),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1090),
.A2(n_1142),
.B(n_1165),
.Y(n_1286)
);

AOI221x1_ASAP7_75t_L g1287 ( 
.A1(n_1080),
.A2(n_1089),
.B1(n_1201),
.B2(n_1157),
.C(n_1060),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1099),
.A2(n_1080),
.B(n_1089),
.Y(n_1288)
);

INVx8_ASAP7_75t_L g1289 ( 
.A(n_1099),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1115),
.B(n_1209),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1149),
.A2(n_1080),
.A3(n_1089),
.B(n_1157),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1149),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1201),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1089),
.A2(n_1157),
.B(n_1201),
.C(n_1206),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1157),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1201),
.A2(n_1199),
.B1(n_1016),
.B2(n_1010),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1187),
.A2(n_1185),
.B(n_1160),
.Y(n_1297)
);

AOI221xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1206),
.A2(n_1207),
.B1(n_580),
.B2(n_826),
.C(n_806),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1010),
.C(n_1016),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1199),
.B(n_748),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1072),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1206),
.A2(n_1213),
.B1(n_1207),
.B2(n_692),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1187),
.A2(n_1185),
.B(n_1160),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1200),
.A2(n_1203),
.B(n_1202),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1148),
.A2(n_1191),
.B(n_1053),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1196),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1196),
.A2(n_1188),
.B(n_1091),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1196),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1059),
.B(n_726),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_SL g1310 ( 
.A1(n_1147),
.A2(n_1145),
.B(n_1207),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1206),
.A2(n_906),
.A3(n_1188),
.B(n_1091),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1199),
.C(n_1016),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1213),
.B(n_945),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1187),
.A2(n_1185),
.B(n_1160),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1199),
.A2(n_1016),
.B1(n_1010),
.B2(n_748),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1010),
.C(n_1016),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1200),
.A2(n_715),
.B(n_1211),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1199),
.C(n_1016),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1200),
.A2(n_1203),
.B(n_1202),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1206),
.B(n_1213),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1200),
.A2(n_715),
.B(n_1211),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1080),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1206),
.A2(n_906),
.A3(n_1188),
.B(n_1091),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1010),
.C(n_1016),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1176),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1083),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1176),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1144),
.Y(n_1328)
);

NOR2xp67_ASAP7_75t_L g1329 ( 
.A(n_1105),
.B(n_708),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1200),
.A2(n_715),
.B(n_1211),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1200),
.A2(n_715),
.B(n_1211),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_SL g1332 ( 
.A1(n_1206),
.A2(n_1197),
.B(n_1207),
.C(n_1077),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1199),
.C(n_1016),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1196),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1187),
.A2(n_1185),
.B(n_1160),
.Y(n_1335)
);

AOI31xp67_ASAP7_75t_L g1336 ( 
.A1(n_1191),
.A2(n_1193),
.A3(n_1077),
.B(n_1036),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1199),
.C(n_1016),
.Y(n_1337)
);

AO22x2_ASAP7_75t_L g1338 ( 
.A1(n_1199),
.A2(n_1137),
.B1(n_1079),
.B2(n_1104),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1196),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1206),
.A2(n_906),
.A3(n_1188),
.B(n_1091),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1200),
.A2(n_1203),
.B(n_1202),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1176),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1066),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1059),
.B(n_726),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1199),
.C(n_1016),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1206),
.A2(n_1213),
.B1(n_1207),
.B2(n_692),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1200),
.A2(n_1203),
.B(n_1202),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1206),
.B(n_1213),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1094),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1200),
.A2(n_1203),
.B(n_1202),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1206),
.B(n_1213),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1200),
.A2(n_1203),
.B(n_1202),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1200),
.A2(n_1203),
.B(n_1202),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1176),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1206),
.B(n_1213),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1187),
.A2(n_1185),
.B(n_1160),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1206),
.A2(n_906),
.A3(n_1188),
.B(n_1091),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1094),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1176),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1200),
.A2(n_715),
.B(n_1211),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1134),
.A2(n_726),
.B1(n_800),
.B2(n_867),
.Y(n_1361)
);

AOI211xp5_ASAP7_75t_L g1362 ( 
.A1(n_1199),
.A2(n_1010),
.B(n_1016),
.C(n_580),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1059),
.B(n_726),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1206),
.B(n_1213),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1080),
.Y(n_1365)
);

AOI31xp67_ASAP7_75t_L g1366 ( 
.A1(n_1191),
.A2(n_1193),
.A3(n_1077),
.B(n_1036),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1148),
.A2(n_1191),
.B(n_1053),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1206),
.B(n_1213),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1083),
.Y(n_1369)
);

OR2x6_ASAP7_75t_L g1370 ( 
.A(n_1062),
.B(n_1144),
.Y(n_1370)
);

NOR2xp67_ASAP7_75t_L g1371 ( 
.A(n_1105),
.B(n_708),
.Y(n_1371)
);

AO31x2_ASAP7_75t_L g1372 ( 
.A1(n_1206),
.A2(n_906),
.A3(n_1188),
.B(n_1091),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1222),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1313),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1260),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1289),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1241),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1325),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1327),
.Y(n_1379)
);

INVx6_ASAP7_75t_L g1380 ( 
.A(n_1289),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1315),
.A2(n_1338),
.B1(n_1300),
.B2(n_1296),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1338),
.A2(n_1224),
.B1(n_1344),
.B2(n_1363),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1362),
.A2(n_1361),
.B1(n_1235),
.B2(n_1309),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1265),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1215),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_SL g1386 ( 
.A1(n_1338),
.A2(n_1256),
.B1(n_1346),
.B2(n_1302),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1256),
.A2(n_1346),
.B1(n_1302),
.B2(n_1339),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1234),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1227),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1306),
.A2(n_1308),
.B1(n_1334),
.B2(n_1339),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1299),
.A2(n_1316),
.B1(n_1324),
.B2(n_1320),
.Y(n_1391)
);

INVx6_ASAP7_75t_L g1392 ( 
.A(n_1247),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1214),
.Y(n_1393)
);

CKINVDCx6p67_ASAP7_75t_R g1394 ( 
.A(n_1262),
.Y(n_1394)
);

INVx4_ASAP7_75t_L g1395 ( 
.A(n_1277),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1306),
.A2(n_1308),
.B1(n_1334),
.B2(n_1220),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1220),
.A2(n_1224),
.B1(n_1310),
.B2(n_1245),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1342),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1261),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1269),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1343),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1320),
.A2(n_1368),
.B1(n_1364),
.B2(n_1355),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1245),
.A2(n_1282),
.B1(n_1368),
.B2(n_1364),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1348),
.A2(n_1355),
.B1(n_1351),
.B2(n_1259),
.Y(n_1404)
);

BUFx12f_ASAP7_75t_L g1405 ( 
.A(n_1328),
.Y(n_1405)
);

BUFx4f_ASAP7_75t_L g1406 ( 
.A(n_1328),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1267),
.Y(n_1407)
);

INVx4_ASAP7_75t_SL g1408 ( 
.A(n_1291),
.Y(n_1408)
);

BUFx2_ASAP7_75t_SL g1409 ( 
.A(n_1349),
.Y(n_1409)
);

CKINVDCx11_ASAP7_75t_R g1410 ( 
.A(n_1328),
.Y(n_1410)
);

BUFx10_ASAP7_75t_L g1411 ( 
.A(n_1265),
.Y(n_1411)
);

OAI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1252),
.A2(n_1329),
.B1(n_1371),
.B2(n_1348),
.Y(n_1412)
);

BUFx4f_ASAP7_75t_SL g1413 ( 
.A(n_1358),
.Y(n_1413)
);

BUFx8_ASAP7_75t_L g1414 ( 
.A(n_1292),
.Y(n_1414)
);

OAI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1351),
.A2(n_1250),
.B1(n_1301),
.B2(n_1370),
.Y(n_1415)
);

BUFx2_ASAP7_75t_SL g1416 ( 
.A(n_1264),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1354),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1369),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1359),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_SL g1420 ( 
.A(n_1370),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1250),
.B(n_1249),
.Y(n_1421)
);

CKINVDCx6p67_ASAP7_75t_R g1422 ( 
.A(n_1370),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1268),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1263),
.A2(n_1312),
.B1(n_1318),
.B2(n_1333),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1237),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1247),
.Y(n_1426)
);

CKINVDCx16_ASAP7_75t_R g1427 ( 
.A(n_1290),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1275),
.A2(n_1298),
.B1(n_1236),
.B2(n_1332),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1249),
.A2(n_1238),
.B1(n_1282),
.B2(n_1239),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1247),
.Y(n_1430)
);

BUFx8_ASAP7_75t_L g1431 ( 
.A(n_1279),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1271),
.Y(n_1432)
);

INVx5_ASAP7_75t_L g1433 ( 
.A(n_1251),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1268),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1326),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1268),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1238),
.A2(n_1239),
.B1(n_1246),
.B2(n_1218),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1230),
.Y(n_1438)
);

INVx6_ASAP7_75t_L g1439 ( 
.A(n_1278),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1337),
.A2(n_1345),
.B1(n_1280),
.B2(n_1272),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1240),
.A2(n_1270),
.B1(n_1287),
.B2(n_1254),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1285),
.A2(n_1242),
.B1(n_1307),
.B2(n_1218),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1281),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1246),
.A2(n_1253),
.B1(n_1285),
.B2(n_1266),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_1273),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1221),
.A2(n_1229),
.B(n_1232),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1248),
.A2(n_1286),
.B1(n_1273),
.B2(n_1266),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1251),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1229),
.B(n_1232),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1293),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1295),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1286),
.A2(n_1281),
.B1(n_1307),
.B2(n_1228),
.Y(n_1452)
);

OAI22x1_ASAP7_75t_L g1453 ( 
.A1(n_1233),
.A2(n_1274),
.B1(n_1367),
.B2(n_1305),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1276),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1231),
.A2(n_1223),
.B1(n_1243),
.B2(n_1217),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1284),
.Y(n_1456)
);

CKINVDCx11_ASAP7_75t_R g1457 ( 
.A(n_1294),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1255),
.A2(n_1219),
.B1(n_1365),
.B2(n_1322),
.Y(n_1458)
);

BUFx10_ASAP7_75t_L g1459 ( 
.A(n_1365),
.Y(n_1459)
);

CKINVDCx6p67_ASAP7_75t_R g1460 ( 
.A(n_1288),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1317),
.A2(n_1321),
.B1(n_1330),
.B2(n_1331),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1244),
.A2(n_1360),
.B1(n_1283),
.B2(n_1225),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1216),
.A2(n_1341),
.B1(n_1347),
.B2(n_1350),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_SL g1464 ( 
.A(n_1257),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1216),
.A2(n_1353),
.B1(n_1319),
.B2(n_1341),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1217),
.B(n_1226),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1284),
.B(n_1323),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1304),
.A2(n_1347),
.B1(n_1319),
.B2(n_1350),
.Y(n_1468)
);

INVx4_ASAP7_75t_L g1469 ( 
.A(n_1284),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1304),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1352),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1352),
.A2(n_1353),
.B1(n_1258),
.B2(n_1226),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1258),
.A2(n_1323),
.B1(n_1357),
.B2(n_1340),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1258),
.A2(n_1323),
.B1(n_1357),
.B2(n_1340),
.Y(n_1474)
);

BUFx12f_ASAP7_75t_L g1475 ( 
.A(n_1336),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1311),
.A2(n_1372),
.B1(n_1357),
.B2(n_1340),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1372),
.A2(n_1366),
.B(n_1303),
.Y(n_1477)
);

INVx6_ASAP7_75t_L g1478 ( 
.A(n_1297),
.Y(n_1478)
);

INVx6_ASAP7_75t_L g1479 ( 
.A(n_1314),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1335),
.A2(n_1199),
.B1(n_1016),
.B2(n_1010),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1356),
.A2(n_1206),
.B1(n_1316),
.B2(n_1299),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1289),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1315),
.A2(n_1199),
.B1(n_1016),
.B2(n_1010),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1278),
.B(n_1247),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1220),
.A2(n_1232),
.B(n_1306),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1338),
.A2(n_867),
.B1(n_1010),
.B2(n_1134),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1338),
.A2(n_867),
.B1(n_1010),
.B2(n_1134),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1234),
.B(n_1074),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1315),
.A2(n_1199),
.B1(n_1016),
.B2(n_1010),
.Y(n_1489)
);

BUFx8_ASAP7_75t_L g1490 ( 
.A(n_1328),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1315),
.A2(n_1199),
.B1(n_1016),
.B2(n_1010),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1265),
.Y(n_1492)
);

CKINVDCx11_ASAP7_75t_R g1493 ( 
.A(n_1262),
.Y(n_1493)
);

CKINVDCx11_ASAP7_75t_R g1494 ( 
.A(n_1262),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1222),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1320),
.B(n_1348),
.Y(n_1496)
);

AOI21xp33_ASAP7_75t_L g1497 ( 
.A1(n_1312),
.A2(n_1333),
.B(n_1318),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1222),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1338),
.A2(n_867),
.B1(n_1010),
.B2(n_1134),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1222),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1214),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1222),
.Y(n_1502)
);

OAI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1315),
.A2(n_1016),
.B(n_1010),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1289),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1222),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1289),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1315),
.A2(n_1199),
.B1(n_1016),
.B2(n_1010),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1315),
.A2(n_1199),
.B1(n_1016),
.B2(n_1010),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1423),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1470),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1434),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1445),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1445),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1436),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1456),
.Y(n_1515)
);

INVxp33_ASAP7_75t_SL g1516 ( 
.A(n_1385),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1389),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1466),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1392),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1396),
.B(n_1390),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1396),
.B(n_1390),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1466),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1465),
.A2(n_1472),
.B(n_1468),
.Y(n_1523)
);

OAI21xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1429),
.A2(n_1402),
.B(n_1404),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1386),
.B(n_1397),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1503),
.A2(n_1508),
.B1(n_1507),
.B2(n_1491),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1386),
.B(n_1397),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1467),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1454),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1485),
.B(n_1382),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1421),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1465),
.A2(n_1472),
.B(n_1462),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1449),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1449),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_SL g1535 ( 
.A(n_1430),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1485),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1389),
.Y(n_1537)
);

AO31x2_ASAP7_75t_L g1538 ( 
.A1(n_1473),
.A2(n_1453),
.A3(n_1481),
.B(n_1391),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1478),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1483),
.A2(n_1489),
.B1(n_1424),
.B2(n_1487),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1446),
.A2(n_1461),
.B(n_1463),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1497),
.A2(n_1440),
.B(n_1424),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1481),
.B(n_1478),
.Y(n_1543)
);

NAND2x1_ASAP7_75t_L g1544 ( 
.A(n_1447),
.B(n_1469),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1473),
.A2(n_1446),
.B(n_1437),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_1471),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1464),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1408),
.B(n_1452),
.Y(n_1548)
);

AO21x2_ASAP7_75t_L g1549 ( 
.A1(n_1474),
.A2(n_1477),
.B(n_1476),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1475),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1408),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1496),
.B(n_1391),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1497),
.A2(n_1440),
.B(n_1383),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1373),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1378),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1379),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1479),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1458),
.A2(n_1444),
.B(n_1480),
.Y(n_1558)
);

INVx4_ASAP7_75t_L g1559 ( 
.A(n_1460),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1486),
.A2(n_1499),
.B1(n_1487),
.B2(n_1403),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1398),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1417),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1419),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1418),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1486),
.A2(n_1499),
.B1(n_1457),
.B2(n_1381),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1433),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1495),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1428),
.A2(n_1505),
.B(n_1502),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1498),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1500),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1442),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1412),
.A2(n_1415),
.B1(n_1387),
.B2(n_1488),
.Y(n_1572)
);

BUFx2_ASAP7_75t_SL g1573 ( 
.A(n_1420),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1377),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1442),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1438),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1432),
.B(n_1403),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1443),
.A2(n_1455),
.B(n_1387),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1455),
.Y(n_1579)
);

NAND2x1p5_ASAP7_75t_L g1580 ( 
.A(n_1376),
.B(n_1482),
.Y(n_1580)
);

AOI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1401),
.A2(n_1484),
.B(n_1492),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1435),
.Y(n_1582)
);

AOI21xp33_ASAP7_75t_L g1583 ( 
.A1(n_1441),
.A2(n_1374),
.B(n_1388),
.Y(n_1583)
);

AOI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1484),
.A2(n_1384),
.B(n_1393),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1400),
.B(n_1427),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1459),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1425),
.A2(n_1420),
.B1(n_1426),
.B2(n_1422),
.Y(n_1587)
);

OA21x2_ASAP7_75t_L g1588 ( 
.A1(n_1450),
.A2(n_1451),
.B(n_1395),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1448),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1380),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1411),
.B(n_1504),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1431),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1411),
.B(n_1506),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1546),
.B(n_1409),
.Y(n_1594)
);

AO21x2_ASAP7_75t_L g1595 ( 
.A1(n_1542),
.A2(n_1431),
.B(n_1414),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1546),
.B(n_1399),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1542),
.A2(n_1506),
.B(n_1406),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1516),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1555),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1553),
.A2(n_1406),
.B1(n_1501),
.B2(n_1416),
.C(n_1439),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_SL g1601 ( 
.A1(n_1560),
.A2(n_1493),
.B(n_1494),
.C(n_1490),
.Y(n_1601)
);

OAI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1553),
.A2(n_1506),
.B(n_1414),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1531),
.B(n_1439),
.Y(n_1603)
);

AO32x2_ASAP7_75t_L g1604 ( 
.A1(n_1560),
.A2(n_1490),
.A3(n_1413),
.B1(n_1410),
.B2(n_1394),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1510),
.B(n_1439),
.Y(n_1605)
);

AO32x2_ASAP7_75t_L g1606 ( 
.A1(n_1539),
.A2(n_1375),
.A3(n_1405),
.B1(n_1407),
.B2(n_1557),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1554),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1537),
.Y(n_1608)
);

OR2x6_ASAP7_75t_L g1609 ( 
.A(n_1543),
.B(n_1544),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1540),
.A2(n_1526),
.B1(n_1565),
.B2(n_1520),
.Y(n_1610)
);

O2A1O1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1524),
.A2(n_1583),
.B(n_1521),
.C(n_1577),
.Y(n_1611)
);

OR2x6_ASAP7_75t_L g1612 ( 
.A(n_1543),
.B(n_1544),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1533),
.B(n_1534),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1524),
.A2(n_1521),
.B1(n_1525),
.B2(n_1527),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1512),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1558),
.A2(n_1572),
.B(n_1583),
.Y(n_1616)
);

AO21x1_ASAP7_75t_L g1617 ( 
.A1(n_1525),
.A2(n_1527),
.B(n_1577),
.Y(n_1617)
);

A2O1A1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1558),
.A2(n_1523),
.B(n_1552),
.C(n_1545),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1552),
.A2(n_1585),
.B1(n_1517),
.B2(n_1513),
.Y(n_1619)
);

NAND3xp33_ASAP7_75t_L g1620 ( 
.A(n_1582),
.B(n_1530),
.C(n_1559),
.Y(n_1620)
);

AO32x2_ASAP7_75t_L g1621 ( 
.A1(n_1539),
.A2(n_1557),
.A3(n_1519),
.B1(n_1566),
.B2(n_1559),
.Y(n_1621)
);

A2O1A1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1558),
.A2(n_1523),
.B(n_1545),
.C(n_1530),
.Y(n_1622)
);

OAI211xp5_ASAP7_75t_L g1623 ( 
.A1(n_1571),
.A2(n_1575),
.B(n_1576),
.C(n_1587),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1588),
.B(n_1564),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1588),
.B(n_1564),
.Y(n_1625)
);

A2O1A1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1523),
.A2(n_1532),
.B(n_1571),
.C(n_1575),
.Y(n_1626)
);

CKINVDCx6p67_ASAP7_75t_R g1627 ( 
.A(n_1573),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1588),
.B(n_1547),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1528),
.B(n_1563),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1584),
.Y(n_1630)
);

OA21x2_ASAP7_75t_L g1631 ( 
.A1(n_1532),
.A2(n_1536),
.B(n_1579),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1541),
.A2(n_1528),
.B1(n_1562),
.B2(n_1567),
.C(n_1570),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1541),
.A2(n_1562),
.B1(n_1567),
.B2(n_1561),
.C(n_1570),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_L g1634 ( 
.A(n_1559),
.B(n_1588),
.C(n_1589),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1592),
.B(n_1593),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1543),
.B(n_1548),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1556),
.B(n_1561),
.Y(n_1637)
);

OR2x6_ASAP7_75t_L g1638 ( 
.A(n_1543),
.B(n_1548),
.Y(n_1638)
);

AO32x2_ASAP7_75t_L g1639 ( 
.A1(n_1539),
.A2(n_1557),
.A3(n_1519),
.B1(n_1566),
.B2(n_1590),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1556),
.B(n_1569),
.Y(n_1640)
);

AO32x1_ASAP7_75t_L g1641 ( 
.A1(n_1511),
.A2(n_1515),
.A3(n_1509),
.B1(n_1514),
.B2(n_1566),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1518),
.B(n_1522),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1541),
.A2(n_1569),
.B1(n_1522),
.B2(n_1518),
.C(n_1573),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1581),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1568),
.B(n_1574),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1644),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1636),
.B(n_1638),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1622),
.B(n_1549),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1610),
.A2(n_1578),
.B1(n_1543),
.B2(n_1535),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1618),
.B(n_1549),
.Y(n_1650)
);

INVx4_ASAP7_75t_R g1651 ( 
.A(n_1624),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1631),
.B(n_1645),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1610),
.A2(n_1578),
.B1(n_1535),
.B2(n_1549),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1607),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1645),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1626),
.B(n_1578),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1621),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1629),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1613),
.B(n_1538),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1641),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1613),
.B(n_1538),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1617),
.A2(n_1535),
.B1(n_1548),
.B2(n_1519),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1614),
.A2(n_1535),
.B1(n_1550),
.B2(n_1591),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1639),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1637),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1639),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1639),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1600),
.A2(n_1590),
.B(n_1580),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1640),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1634),
.B(n_1538),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1628),
.B(n_1529),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1616),
.B(n_1550),
.C(n_1586),
.Y(n_1672)
);

OR2x6_ASAP7_75t_SL g1673 ( 
.A(n_1634),
.B(n_1551),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1655),
.B(n_1633),
.Y(n_1674)
);

AND2x2_ASAP7_75t_SL g1675 ( 
.A(n_1656),
.B(n_1643),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1646),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1654),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1655),
.B(n_1608),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1646),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1659),
.B(n_1632),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1652),
.Y(n_1681)
);

OAI33xp33_ASAP7_75t_L g1682 ( 
.A1(n_1660),
.A2(n_1619),
.A3(n_1611),
.B1(n_1599),
.B2(n_1603),
.B3(n_1642),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1673),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1657),
.B(n_1625),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1659),
.B(n_1615),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1654),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1647),
.B(n_1620),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1652),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1653),
.A2(n_1614),
.B1(n_1612),
.B2(n_1609),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1657),
.B(n_1621),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1668),
.B(n_1627),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1652),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1664),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1653),
.B(n_1623),
.C(n_1601),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1671),
.B(n_1620),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1647),
.B(n_1630),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1661),
.B(n_1658),
.Y(n_1697)
);

INVx5_ASAP7_75t_L g1698 ( 
.A(n_1657),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1681),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1674),
.B(n_1664),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1690),
.B(n_1657),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1680),
.B(n_1658),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1690),
.B(n_1657),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1674),
.B(n_1666),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1683),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1677),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1690),
.B(n_1657),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1680),
.B(n_1665),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1676),
.B(n_1665),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1683),
.B(n_1672),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1676),
.B(n_1665),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1677),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1694),
.A2(n_1649),
.B1(n_1602),
.B2(n_1662),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1691),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1698),
.B(n_1684),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1686),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1679),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1698),
.B(n_1657),
.Y(n_1718)
);

NAND2x1p5_ASAP7_75t_L g1719 ( 
.A(n_1698),
.B(n_1670),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1698),
.B(n_1657),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1693),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1698),
.B(n_1657),
.Y(n_1722)
);

INVx4_ASAP7_75t_L g1723 ( 
.A(n_1698),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1698),
.B(n_1666),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1681),
.B(n_1666),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1687),
.B(n_1696),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1697),
.B(n_1666),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1687),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1686),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1679),
.B(n_1669),
.Y(n_1730)
);

INVxp67_ASAP7_75t_L g1731 ( 
.A(n_1682),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1687),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1697),
.B(n_1667),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1685),
.B(n_1669),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1693),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1731),
.B(n_1675),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1715),
.B(n_1675),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1706),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1731),
.B(n_1675),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1706),
.Y(n_1740)
);

INVxp67_ASAP7_75t_SL g1741 ( 
.A(n_1710),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1705),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1702),
.B(n_1708),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1710),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1725),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1723),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1712),
.Y(n_1747)
);

NAND2x1_ASAP7_75t_L g1748 ( 
.A(n_1723),
.B(n_1651),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1702),
.B(n_1685),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1712),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1700),
.B(n_1678),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1716),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1716),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1700),
.B(n_1678),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1729),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1725),
.Y(n_1756)
);

NAND2x1_ASAP7_75t_L g1757 ( 
.A(n_1723),
.B(n_1651),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1714),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1708),
.B(n_1695),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1715),
.B(n_1696),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1715),
.B(n_1696),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1728),
.B(n_1696),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1704),
.B(n_1681),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1704),
.B(n_1688),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1729),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1723),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1705),
.B(n_1688),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1734),
.B(n_1688),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1734),
.B(n_1692),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1713),
.B(n_1695),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1717),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1717),
.B(n_1692),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1709),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1709),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1728),
.B(n_1687),
.Y(n_1775)
);

NOR2x1_ASAP7_75t_SL g1776 ( 
.A(n_1718),
.B(n_1689),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1711),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1725),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1736),
.B(n_1714),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1739),
.B(n_1714),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1742),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1752),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1758),
.B(n_1713),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1752),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1737),
.B(n_1718),
.Y(n_1785)
);

INVx3_ASAP7_75t_L g1786 ( 
.A(n_1748),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1770),
.B(n_1711),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1771),
.B(n_1730),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1737),
.B(n_1718),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1743),
.B(n_1730),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1742),
.B(n_1724),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1749),
.B(n_1724),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1753),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1753),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1759),
.B(n_1724),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1751),
.B(n_1727),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1751),
.B(n_1727),
.Y(n_1797)
);

AND2x2_ASAP7_75t_SL g1798 ( 
.A(n_1741),
.B(n_1656),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1754),
.B(n_1733),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1767),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1776),
.B(n_1720),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1776),
.B(n_1720),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1760),
.B(n_1720),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1744),
.B(n_1773),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1738),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1774),
.B(n_1701),
.Y(n_1806)
);

NAND2x1p5_ASAP7_75t_L g1807 ( 
.A(n_1748),
.B(n_1722),
.Y(n_1807)
);

AOI32xp33_ASAP7_75t_L g1808 ( 
.A1(n_1775),
.A2(n_1656),
.A3(n_1701),
.B1(n_1703),
.B2(n_1707),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1740),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1754),
.B(n_1767),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1747),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1777),
.B(n_1775),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1745),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1750),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1781),
.B(n_1766),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1782),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1785),
.B(n_1789),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1785),
.B(n_1760),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1798),
.A2(n_1694),
.B1(n_1673),
.B2(n_1757),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1798),
.B(n_1766),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1801),
.Y(n_1821)
);

OAI222xp33_ASAP7_75t_L g1822 ( 
.A1(n_1808),
.A2(n_1719),
.B1(n_1757),
.B2(n_1689),
.C1(n_1701),
.C2(n_1707),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1783),
.A2(n_1808),
.B1(n_1779),
.B2(n_1780),
.C(n_1787),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1789),
.B(n_1761),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1807),
.A2(n_1673),
.B1(n_1670),
.B2(n_1732),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1798),
.A2(n_1673),
.B1(n_1649),
.B2(n_1662),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1781),
.B(n_1762),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1800),
.B(n_1762),
.Y(n_1828)
);

AO22x2_ASAP7_75t_L g1829 ( 
.A1(n_1801),
.A2(n_1746),
.B1(n_1722),
.B2(n_1703),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1810),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1782),
.Y(n_1831)
);

OAI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1807),
.A2(n_1719),
.B1(n_1746),
.B2(n_1732),
.C(n_1722),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1802),
.B(n_1761),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1784),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1784),
.Y(n_1835)
);

AOI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1804),
.A2(n_1682),
.B1(n_1703),
.B2(n_1707),
.C(n_1648),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1793),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1793),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1810),
.Y(n_1839)
);

A2O1A1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1802),
.A2(n_1672),
.B(n_1602),
.C(n_1656),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1819),
.A2(n_1648),
.B1(n_1812),
.B2(n_1650),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1826),
.A2(n_1836),
.B1(n_1823),
.B2(n_1817),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1830),
.B(n_1800),
.Y(n_1843)
);

OAI21xp33_ASAP7_75t_L g1844 ( 
.A1(n_1827),
.A2(n_1806),
.B(n_1791),
.Y(n_1844)
);

OAI21xp33_ASAP7_75t_L g1845 ( 
.A1(n_1817),
.A2(n_1795),
.B(n_1803),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1818),
.B(n_1803),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1818),
.B(n_1807),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1839),
.A2(n_1821),
.B1(n_1815),
.B2(n_1786),
.Y(n_1848)
);

OAI322xp33_ASAP7_75t_L g1849 ( 
.A1(n_1820),
.A2(n_1788),
.A3(n_1814),
.B1(n_1805),
.B2(n_1811),
.C1(n_1809),
.C2(n_1797),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1838),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1824),
.B(n_1786),
.Y(n_1851)
);

OAI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1820),
.A2(n_1786),
.B(n_1719),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1828),
.B(n_1598),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1824),
.B(n_1746),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1838),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1815),
.B(n_1796),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1816),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1831),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1825),
.B(n_1813),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1815),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1833),
.B(n_1813),
.Y(n_1861)
);

NAND2x1p5_ASAP7_75t_L g1862 ( 
.A(n_1848),
.B(n_1833),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1856),
.Y(n_1863)
);

A2O1A1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1842),
.A2(n_1840),
.B(n_1832),
.C(n_1835),
.Y(n_1864)
);

NOR3xp33_ASAP7_75t_L g1865 ( 
.A(n_1843),
.B(n_1860),
.C(n_1849),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1856),
.Y(n_1866)
);

AND2x2_ASAP7_75t_SL g1867 ( 
.A(n_1853),
.B(n_1834),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1861),
.B(n_1829),
.Y(n_1868)
);

AOI321xp33_ASAP7_75t_L g1869 ( 
.A1(n_1859),
.A2(n_1858),
.A3(n_1857),
.B1(n_1844),
.B2(n_1841),
.C(n_1855),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1859),
.A2(n_1840),
.B1(n_1847),
.B2(n_1846),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1861),
.B(n_1829),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1851),
.Y(n_1872)
);

NOR2x1_ASAP7_75t_SL g1873 ( 
.A(n_1847),
.B(n_1837),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1863),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1872),
.B(n_1846),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1866),
.B(n_1851),
.Y(n_1876)
);

OAI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1862),
.A2(n_1852),
.B1(n_1719),
.B2(n_1732),
.Y(n_1877)
);

NAND4xp25_ASAP7_75t_L g1878 ( 
.A(n_1869),
.B(n_1845),
.C(n_1854),
.D(n_1850),
.Y(n_1878)
);

NAND4xp25_ASAP7_75t_SL g1879 ( 
.A(n_1864),
.B(n_1854),
.C(n_1822),
.D(n_1850),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1873),
.Y(n_1880)
);

NAND4xp25_ASAP7_75t_L g1881 ( 
.A(n_1869),
.B(n_1805),
.C(n_1814),
.D(n_1811),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1867),
.B(n_1829),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1865),
.B(n_1829),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1879),
.A2(n_1870),
.B1(n_1871),
.B2(n_1868),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1882),
.B(n_1809),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1883),
.A2(n_1794),
.B1(n_1790),
.B2(n_1792),
.C(n_1796),
.Y(n_1886)
);

OAI321xp33_ASAP7_75t_L g1887 ( 
.A1(n_1878),
.A2(n_1794),
.A3(n_1799),
.B1(n_1797),
.B2(n_1672),
.C(n_1663),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1875),
.B(n_1799),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1885),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1884),
.A2(n_1877),
.B1(n_1876),
.B2(n_1880),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1888),
.A2(n_1881),
.B1(n_1874),
.B2(n_1648),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1886),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1887),
.Y(n_1893)
);

OAI31xp33_ASAP7_75t_L g1894 ( 
.A1(n_1884),
.A2(n_1732),
.A3(n_1772),
.B(n_1763),
.Y(n_1894)
);

NOR2x1_ASAP7_75t_L g1895 ( 
.A(n_1889),
.B(n_1772),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1890),
.B(n_1755),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1893),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1893),
.Y(n_1898)
);

OAI211xp5_ASAP7_75t_L g1899 ( 
.A1(n_1892),
.A2(n_1778),
.B(n_1745),
.C(n_1756),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1895),
.Y(n_1900)
);

O2A1O1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1897),
.A2(n_1894),
.B(n_1891),
.C(n_1778),
.Y(n_1901)
);

NOR3xp33_ASAP7_75t_L g1902 ( 
.A(n_1898),
.B(n_1635),
.C(n_1596),
.Y(n_1902)
);

AOI22x1_ASAP7_75t_L g1903 ( 
.A1(n_1900),
.A2(n_1896),
.B1(n_1899),
.B2(n_1756),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1903),
.A2(n_1902),
.B1(n_1901),
.B2(n_1595),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1904),
.A2(n_1764),
.B1(n_1763),
.B2(n_1765),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1904),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1906),
.B(n_1764),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_SL g1908 ( 
.A1(n_1905),
.A2(n_1735),
.B1(n_1721),
.B2(n_1726),
.Y(n_1908)
);

OAI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1907),
.A2(n_1769),
.B(n_1768),
.Y(n_1909)
);

OAI21x1_ASAP7_75t_L g1910 ( 
.A1(n_1908),
.A2(n_1769),
.B(n_1768),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_SL g1911 ( 
.A1(n_1909),
.A2(n_1735),
.B1(n_1721),
.B2(n_1726),
.Y(n_1911)
);

AOI21xp33_ASAP7_75t_L g1912 ( 
.A1(n_1911),
.A2(n_1910),
.B(n_1595),
.Y(n_1912)
);

OAI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1912),
.A2(n_1699),
.B1(n_1733),
.B2(n_1692),
.Y(n_1913)
);

OAI221xp5_ASAP7_75t_R g1914 ( 
.A1(n_1913),
.A2(n_1663),
.B1(n_1604),
.B2(n_1606),
.C(n_1726),
.Y(n_1914)
);

AOI211xp5_ASAP7_75t_L g1915 ( 
.A1(n_1914),
.A2(n_1597),
.B(n_1594),
.C(n_1605),
.Y(n_1915)
);


endmodule