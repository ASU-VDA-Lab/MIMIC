module fake_ibex_1321_n_1482 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_300, n_103, n_95, n_205, n_204, n_285, n_139, n_247, n_274, n_288, n_55, n_130, n_275, n_291, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_267, n_268, n_8, n_118, n_224, n_273, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_287, n_110, n_193, n_293, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_299, n_27, n_165, n_242, n_278, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_301, n_59, n_28, n_125, n_304, n_39, n_296, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_303, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_282, n_14, n_0, n_239, n_289, n_94, n_134, n_12, n_266, n_42, n_77, n_112, n_257, n_294, n_150, n_286, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_284, n_80, n_172, n_215, n_250, n_279, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_281, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_280, n_269, n_302, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_283, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_297, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_270, n_295, n_230, n_96, n_185, n_271, n_241, n_68, n_117, n_292, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_298, n_158, n_211, n_290, n_218, n_259, n_132, n_174, n_276, n_277, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_272, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1482);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_300;
input n_103;
input n_95;
input n_205;
input n_204;
input n_285;
input n_139;
input n_247;
input n_274;
input n_288;
input n_55;
input n_130;
input n_275;
input n_291;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_267;
input n_268;
input n_8;
input n_118;
input n_224;
input n_273;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_287;
input n_110;
input n_193;
input n_293;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_299;
input n_27;
input n_165;
input n_242;
input n_278;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_301;
input n_59;
input n_28;
input n_125;
input n_304;
input n_39;
input n_296;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_303;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_282;
input n_14;
input n_0;
input n_239;
input n_289;
input n_94;
input n_134;
input n_12;
input n_266;
input n_42;
input n_77;
input n_112;
input n_257;
input n_294;
input n_150;
input n_286;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_284;
input n_80;
input n_172;
input n_215;
input n_250;
input n_279;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_281;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_280;
input n_269;
input n_302;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_283;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_297;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_270;
input n_295;
input n_230;
input n_96;
input n_185;
input n_271;
input n_241;
input n_68;
input n_117;
input n_292;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_158;
input n_211;
input n_290;
input n_218;
input n_259;
input n_132;
input n_174;
input n_276;
input n_277;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_272;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1482;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_1340;
wire n_339;
wire n_348;
wire n_674;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_716;
wire n_923;
wire n_642;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_354;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_1047;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1433;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1369;
wire n_1297;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_141),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_36),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_4),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_11),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_159),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_100),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_238),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_49),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_208),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_132),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_214),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_153),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_269),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_301),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_23),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_86),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_199),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_71),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_144),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_242),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_149),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_233),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_118),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_38),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_75),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_223),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_155),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_160),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_251),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_75),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_295),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_78),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_98),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_175),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_112),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_171),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_192),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_86),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_24),
.Y(n_344)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_243),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_207),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_191),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_68),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_49),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_174),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_188),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_9),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_274),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_2),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_273),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_225),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_247),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_200),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_125),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_280),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_236),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_235),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_156),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_152),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_227),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_281),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_136),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_101),
.B(n_255),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_163),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_190),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_265),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_148),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_219),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_26),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_186),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_183),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_139),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_48),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_147),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_258),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_26),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_76),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_173),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_293),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_143),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_260),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_100),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_42),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_212),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_162),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_30),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_180),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_176),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_285),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_220),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_246),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_83),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_193),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_119),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_150),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_38),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_88),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_73),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_275),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_6),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_287),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_195),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_73),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_57),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_303),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_264),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_237),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_62),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_71),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_267),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_138),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_84),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_202),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_291),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_11),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_64),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_137),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_106),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_259),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_47),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_110),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_304),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_296),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_102),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_222),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_217),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_161),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_69),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_256),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_234),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_97),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_289),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_266),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_230),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_221),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_213),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_282),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_5),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_30),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_206),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_58),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_245),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_254),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_224),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_299),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_182),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_239),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_24),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_297),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_302),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_218),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_74),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_142),
.Y(n_458)
);

BUFx5_ASAP7_75t_L g459 ( 
.A(n_131),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_104),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_300),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_40),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_0),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_244),
.B(n_270),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_15),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_232),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_37),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_39),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_185),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_85),
.B(n_19),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_252),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_128),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_27),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_127),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_34),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_145),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_198),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_203),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_44),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_181),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_93),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_39),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_47),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_22),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_68),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_55),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_16),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_29),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_189),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_271),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_248),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_172),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_240),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_250),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_32),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_211),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_116),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_54),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_178),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_120),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_97),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_262),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_37),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_168),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_92),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_96),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_272),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_32),
.Y(n_508)
);

BUFx5_ASAP7_75t_L g509 ( 
.A(n_107),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_0),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_129),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_325),
.B(n_356),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_446),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_349),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_345),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_1),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_501),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_349),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_402),
.B(n_1),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_312),
.B(n_105),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_402),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_467),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_361),
.B(n_3),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_467),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_481),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_345),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_334),
.Y(n_527)
);

BUFx8_ASAP7_75t_L g528 ( 
.A(n_362),
.Y(n_528)
);

BUFx12f_ASAP7_75t_L g529 ( 
.A(n_478),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_481),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_425),
.B(n_6),
.Y(n_531)
);

INVxp33_ASAP7_75t_SL g532 ( 
.A(n_308),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_305),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_485),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_498),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_352),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_325),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_345),
.Y(n_538)
);

BUFx8_ASAP7_75t_L g539 ( 
.A(n_345),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_356),
.B(n_108),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_498),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_485),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_305),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_333),
.B(n_7),
.Y(n_544)
);

BUFx8_ASAP7_75t_SL g545 ( 
.A(n_313),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_345),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_330),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_462),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_305),
.Y(n_549)
);

AOI22x1_ASAP7_75t_R g550 ( 
.A1(n_313),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_316),
.A2(n_111),
.B(n_109),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_347),
.B(n_10),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_316),
.A2(n_114),
.B(n_113),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_400),
.B(n_115),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_336),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_331),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_330),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_331),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_347),
.B(n_12),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_331),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_331),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_489),
.Y(n_562)
);

CKINVDCx11_ASAP7_75t_R g563 ( 
.A(n_382),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_426),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_365),
.B(n_13),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_307),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_315),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_345),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_489),
.B(n_13),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_420),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_345),
.Y(n_571)
);

BUFx8_ASAP7_75t_SL g572 ( 
.A(n_382),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_459),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_364),
.A2(n_324),
.B(n_318),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_426),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_426),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_326),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_309),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_327),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_431),
.B(n_14),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_426),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_454),
.B(n_14),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_311),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_493),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_337),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_344),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_493),
.B(n_15),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_502),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_502),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_306),
.B(n_16),
.Y(n_590)
);

OA21x2_ASAP7_75t_L g591 ( 
.A1(n_364),
.A2(n_121),
.B(n_117),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_354),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_459),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_320),
.B(n_17),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_459),
.Y(n_595)
);

BUFx12f_ASAP7_75t_L g596 ( 
.A(n_352),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_459),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_459),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_342),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_443),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_372),
.Y(n_601)
);

NAND2x1p5_ASAP7_75t_L g602 ( 
.A(n_350),
.B(n_122),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_330),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_330),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_321),
.B(n_17),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_374),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_403),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_459),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_534),
.B(n_378),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_536),
.B(n_539),
.Y(n_610)
);

INVx8_ASAP7_75t_L g611 ( 
.A(n_512),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_536),
.B(n_380),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_546),
.Y(n_613)
);

BUFx6f_ASAP7_75t_SL g614 ( 
.A(n_569),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_583),
.B(n_352),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_542),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_546),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_571),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_571),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_539),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_583),
.B(n_381),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_SL g622 ( 
.A(n_552),
.B(n_372),
.Y(n_622)
);

INVx8_ASAP7_75t_L g623 ( 
.A(n_512),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_573),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_515),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_585),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_593),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_585),
.B(n_387),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_593),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_539),
.B(n_310),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_539),
.B(n_314),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_593),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_540),
.B(n_459),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_586),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_586),
.B(n_397),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_592),
.B(n_401),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_598),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_598),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_515),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_592),
.B(n_323),
.Y(n_640)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_552),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_598),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_584),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_532),
.B(n_513),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_584),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_578),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_596),
.B(n_528),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_569),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_596),
.B(n_317),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_569),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_566),
.B(n_405),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_569),
.Y(n_652)
);

CKINVDCx16_ASAP7_75t_R g653 ( 
.A(n_529),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_567),
.B(n_408),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_584),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_587),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_519),
.A2(n_335),
.B1(n_338),
.B2(n_329),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_R g658 ( 
.A(n_555),
.B(n_409),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_587),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_577),
.B(n_414),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_584),
.Y(n_661)
);

BUFx6f_ASAP7_75t_SL g662 ( 
.A(n_587),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_SL g663 ( 
.A(n_528),
.B(n_394),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_528),
.B(n_319),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_528),
.B(n_322),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_587),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_608),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_527),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_584),
.Y(n_669)
);

BUFx6f_ASAP7_75t_SL g670 ( 
.A(n_540),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_589),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_606),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_608),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_589),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_517),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_559),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_600),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_529),
.B(n_346),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_559),
.Y(n_679)
);

INVxp33_ASAP7_75t_L g680 ( 
.A(n_570),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_525),
.Y(n_681)
);

BUFx10_ASAP7_75t_L g682 ( 
.A(n_512),
.Y(n_682)
);

BUFx6f_ASAP7_75t_SL g683 ( 
.A(n_540),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_577),
.B(n_328),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_L g685 ( 
.A(n_540),
.B(n_509),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_589),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_526),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_526),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_538),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_525),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_579),
.B(n_417),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_549),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_538),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_512),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_568),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_549),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_579),
.B(n_332),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_519),
.B(n_343),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_568),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_597),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_565),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_565),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_597),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_599),
.B(n_339),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_595),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_574),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_580),
.B(n_348),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_595),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_549),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_530),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_595),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_574),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_574),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_512),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_549),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_599),
.B(n_340),
.Y(n_716)
);

XNOR2x2_ASAP7_75t_L g717 ( 
.A(n_521),
.B(n_487),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_520),
.B(n_341),
.Y(n_718)
);

INVx8_ASAP7_75t_L g719 ( 
.A(n_512),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_544),
.B(n_351),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_531),
.B(n_436),
.C(n_429),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_512),
.Y(n_722)
);

AND3x2_ASAP7_75t_L g723 ( 
.A(n_531),
.B(n_470),
.C(n_389),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_514),
.B(n_518),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_540),
.B(n_509),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_523),
.B(n_353),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_537),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_547),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_563),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_540),
.B(n_509),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_580),
.B(n_388),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_582),
.B(n_391),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_514),
.Y(n_733)
);

NOR2x1p5_ASAP7_75t_L g734 ( 
.A(n_601),
.B(n_413),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_556),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_556),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_582),
.B(n_355),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_556),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_602),
.B(n_358),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_522),
.B(n_524),
.Y(n_740)
);

AND3x2_ASAP7_75t_L g741 ( 
.A(n_550),
.B(n_433),
.C(n_421),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_602),
.B(n_359),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_545),
.Y(n_743)
);

BUFx6f_ASAP7_75t_SL g744 ( 
.A(n_540),
.Y(n_744)
);

BUFx6f_ASAP7_75t_SL g745 ( 
.A(n_554),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_562),
.B(n_588),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_516),
.B(n_473),
.C(n_468),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_562),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_588),
.B(n_360),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_535),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_541),
.B(n_366),
.Y(n_751)
);

CKINVDCx6p67_ASAP7_75t_R g752 ( 
.A(n_554),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_590),
.B(n_367),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_594),
.B(n_373),
.Y(n_754)
);

OAI22xp33_ASAP7_75t_L g755 ( 
.A1(n_521),
.A2(n_444),
.B1(n_503),
.B2(n_443),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_652),
.A2(n_554),
.B1(n_605),
.B2(n_453),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_620),
.B(n_375),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_641),
.B(n_676),
.Y(n_758)
);

OAI221xp5_ASAP7_75t_L g759 ( 
.A1(n_657),
.A2(n_702),
.B1(n_701),
.B2(n_679),
.C(n_721),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_620),
.B(n_376),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_666),
.B(n_379),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_675),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_666),
.B(n_390),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_681),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_672),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_753),
.B(n_357),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_651),
.B(n_554),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_611),
.B(n_554),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_701),
.A2(n_416),
.B1(n_423),
.B2(n_394),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_754),
.B(n_363),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_654),
.B(n_554),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_660),
.B(n_554),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_702),
.A2(n_416),
.B1(n_447),
.B2(n_423),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_612),
.B(n_369),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_656),
.A2(n_457),
.B1(n_463),
.B2(n_460),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_644),
.A2(n_548),
.B1(n_447),
.B2(n_466),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_659),
.A2(n_466),
.B1(n_469),
.B2(n_455),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_726),
.B(n_370),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_691),
.B(n_396),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_679),
.B(n_398),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_720),
.B(n_371),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_680),
.B(n_548),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_626),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_666),
.B(n_406),
.Y(n_784)
);

NOR3xp33_ASAP7_75t_L g785 ( 
.A(n_755),
.B(n_483),
.C(n_482),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_690),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_653),
.B(n_484),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_668),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_614),
.A2(n_465),
.B1(n_479),
.B2(n_475),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_684),
.B(n_377),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_634),
.B(n_486),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_748),
.B(n_415),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_690),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_694),
.B(n_418),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_615),
.A2(n_455),
.B1(n_474),
.B2(n_469),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_697),
.B(n_383),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_704),
.B(n_384),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_733),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_694),
.B(n_419),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_714),
.B(n_427),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_748),
.B(n_439),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_710),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_716),
.B(n_385),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_615),
.B(n_444),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_609),
.B(n_441),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_714),
.B(n_445),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_747),
.B(n_448),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_739),
.B(n_742),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_698),
.B(n_458),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_614),
.A2(n_508),
.B1(n_510),
.B2(n_506),
.Y(n_810)
);

BUFx8_ASAP7_75t_L g811 ( 
.A(n_614),
.Y(n_811)
);

AO22x2_ASAP7_75t_L g812 ( 
.A1(n_717),
.A2(n_392),
.B1(n_395),
.B2(n_393),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_662),
.A2(n_591),
.B1(n_403),
.B2(n_488),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_646),
.B(n_503),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_648),
.A2(n_553),
.B(n_551),
.C(n_404),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_707),
.B(n_505),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_707),
.B(n_505),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_610),
.B(n_472),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_621),
.B(n_476),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_628),
.B(n_491),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_662),
.A2(n_591),
.B1(n_403),
.B2(n_488),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_668),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_731),
.B(n_474),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_640),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_662),
.A2(n_591),
.B1(n_403),
.B2(n_488),
.Y(n_825)
);

OR2x6_ASAP7_75t_L g826 ( 
.A(n_647),
.B(n_551),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_750),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_677),
.Y(n_828)
);

OAI22xp33_ASAP7_75t_L g829 ( 
.A1(n_663),
.A2(n_496),
.B1(n_499),
.B2(n_488),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_L g830 ( 
.A(n_611),
.B(n_509),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_635),
.B(n_492),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_636),
.B(n_500),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_731),
.B(n_504),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_616),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_724),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_740),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_732),
.B(n_507),
.Y(n_837)
);

NOR3xp33_ASAP7_75t_L g838 ( 
.A(n_622),
.B(n_368),
.C(n_399),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_648),
.A2(n_553),
.B(n_407),
.C(n_411),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_727),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_751),
.B(n_410),
.Y(n_841)
);

BUFx12f_ASAP7_75t_L g842 ( 
.A(n_734),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_737),
.B(n_412),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_650),
.A2(n_499),
.B1(n_496),
.B2(n_424),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_650),
.B(n_422),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_727),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_723),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_749),
.B(n_428),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_678),
.B(n_511),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_611),
.B(n_509),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_706),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_729),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_706),
.B(n_386),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_664),
.A2(n_430),
.B(n_434),
.C(n_432),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_682),
.B(n_480),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_712),
.A2(n_435),
.B1(n_438),
.B2(n_437),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_712),
.B(n_497),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_SL g858 ( 
.A1(n_677),
.A2(n_572),
.B1(n_440),
.B2(n_442),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_713),
.B(n_449),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_713),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_625),
.B(n_450),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_625),
.B(n_451),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_746),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_643),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_630),
.B(n_452),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_631),
.B(n_456),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_752),
.A2(n_471),
.B1(n_461),
.B2(n_494),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_639),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_699),
.B(n_477),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_665),
.B(n_509),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_699),
.B(n_490),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_687),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_649),
.B(n_509),
.Y(n_873)
);

AND2x6_ASAP7_75t_SL g874 ( 
.A(n_729),
.B(n_743),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_667),
.B(n_557),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_645),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_611),
.B(n_464),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_741),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_673),
.B(n_603),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_717),
.B(n_18),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_658),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_655),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_718),
.B(n_603),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_613),
.B(n_603),
.Y(n_884)
);

BUFx5_ASAP7_75t_L g885 ( 
.A(n_722),
.Y(n_885)
);

OR2x6_ASAP7_75t_L g886 ( 
.A(n_623),
.B(n_604),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_617),
.B(n_618),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_623),
.B(n_533),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_687),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_622),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_619),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_633),
.A2(n_607),
.B1(n_604),
.B2(n_581),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_L g893 ( 
.A(n_633),
.B(n_18),
.C(n_19),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_661),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_623),
.B(n_533),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_705),
.B(n_533),
.Y(n_896)
);

INVxp33_ASAP7_75t_L g897 ( 
.A(n_661),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_719),
.B(n_688),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_719),
.Y(n_899)
);

NOR2xp67_ASAP7_75t_L g900 ( 
.A(n_728),
.B(n_20),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_685),
.B(n_20),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_705),
.B(n_543),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_725),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_903)
);

NAND3xp33_ASAP7_75t_L g904 ( 
.A(n_730),
.B(n_576),
.C(n_558),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_669),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_730),
.B(n_21),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_670),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_689),
.B(n_576),
.Y(n_908)
);

BUFx5_ASAP7_75t_L g909 ( 
.A(n_670),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_767),
.A2(n_711),
.B(n_708),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_758),
.B(n_624),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_771),
.A2(n_711),
.B(n_627),
.Y(n_912)
);

O2A1O1Ixp5_ASAP7_75t_L g913 ( 
.A1(n_808),
.A2(n_695),
.B(n_700),
.C(n_693),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_765),
.B(n_632),
.C(n_629),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_772),
.A2(n_637),
.B(n_632),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_768),
.A2(n_638),
.B(n_637),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_762),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_860),
.A2(n_642),
.B(n_638),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_851),
.A2(n_762),
.B1(n_856),
.B2(n_782),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_783),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_L g921 ( 
.A(n_878),
.B(n_25),
.Y(n_921)
);

CKINVDCx8_ASAP7_75t_R g922 ( 
.A(n_874),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_826),
.A2(n_703),
.B(n_671),
.Y(n_923)
);

NOR2xp67_ASAP7_75t_L g924 ( 
.A(n_842),
.B(n_25),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_815),
.A2(n_703),
.B(n_671),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_851),
.A2(n_859),
.B(n_857),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_783),
.A2(n_744),
.B1(n_683),
.B2(n_745),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_853),
.A2(n_845),
.B(n_839),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_789),
.B(n_683),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_886),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_824),
.A2(n_759),
.B(n_880),
.C(n_890),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_887),
.A2(n_686),
.B(n_674),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_834),
.A2(n_607),
.B(n_604),
.C(n_564),
.Y(n_933)
);

NOR2xp67_ASAP7_75t_L g934 ( 
.A(n_769),
.B(n_28),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_810),
.B(n_576),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_835),
.B(n_28),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_798),
.Y(n_937)
);

BUFx5_ASAP7_75t_L g938 ( 
.A(n_868),
.Y(n_938)
);

AO22x1_ASAP7_75t_L g939 ( 
.A1(n_811),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_810),
.B(n_576),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_811),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_L g942 ( 
.A(n_773),
.B(n_31),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_777),
.A2(n_604),
.B1(n_607),
.B2(n_564),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_836),
.B(n_35),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_809),
.B(n_36),
.Y(n_945)
);

AOI21xp33_ASAP7_75t_L g946 ( 
.A1(n_890),
.A2(n_40),
.B(n_41),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_813),
.A2(n_825),
.B(n_821),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_821),
.A2(n_825),
.B(n_756),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_775),
.B(n_41),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_775),
.B(n_42),
.Y(n_950)
);

NOR2x1_ASAP7_75t_L g951 ( 
.A(n_787),
.B(n_607),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_833),
.B(n_837),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_823),
.Y(n_953)
);

OAI321xp33_ASAP7_75t_L g954 ( 
.A1(n_829),
.A2(n_560),
.A3(n_561),
.B1(n_564),
.B2(n_575),
.C(n_581),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_791),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_814),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_816),
.B(n_43),
.Y(n_957)
);

INVxp67_ASAP7_75t_SL g958 ( 
.A(n_844),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_838),
.B(n_43),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_827),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_847),
.B(n_44),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_843),
.B(n_45),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_830),
.A2(n_736),
.B(n_735),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_843),
.B(n_46),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_850),
.A2(n_738),
.B(n_696),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_829),
.A2(n_48),
.B(n_50),
.C(n_51),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_779),
.A2(n_696),
.B(n_692),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_891),
.B(n_52),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_886),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_865),
.A2(n_581),
.B(n_564),
.C(n_575),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_903),
.A2(n_893),
.B(n_867),
.C(n_861),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_778),
.B(n_53),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_817),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_804),
.A2(n_581),
.B1(n_575),
.B2(n_561),
.Y(n_974)
);

NAND2x1p5_ASAP7_75t_L g975 ( 
.A(n_899),
.B(n_561),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_849),
.B(n_55),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_788),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_862),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_869),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_795),
.A2(n_575),
.B1(n_581),
.B2(n_58),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_776),
.A2(n_812),
.B1(n_889),
.B2(n_872),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_886),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_822),
.B(n_56),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_871),
.A2(n_56),
.B(n_59),
.C(n_60),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_790),
.B(n_59),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_866),
.A2(n_715),
.B(n_709),
.C(n_62),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_866),
.A2(n_715),
.B(n_63),
.C(n_64),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_881),
.B(n_819),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_764),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_904),
.A2(n_170),
.B(n_294),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_786),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_879),
.A2(n_169),
.B(n_292),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_790),
.B(n_61),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_796),
.B(n_61),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_877),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_774),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_797),
.B(n_65),
.Y(n_997)
);

AND2x6_ASAP7_75t_L g998 ( 
.A(n_907),
.B(n_123),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_828),
.B(n_852),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_793),
.Y(n_1000)
);

AO32x1_ASAP7_75t_L g1001 ( 
.A1(n_901),
.A2(n_66),
.A3(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_792),
.Y(n_1002)
);

AO21x1_ASAP7_75t_L g1003 ( 
.A1(n_906),
.A2(n_70),
.B(n_72),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_812),
.B(n_74),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_812),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_870),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_780),
.A2(n_77),
.B(n_79),
.Y(n_1007)
);

BUFx2_ASAP7_75t_SL g1008 ( 
.A(n_900),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_797),
.B(n_80),
.Y(n_1009)
);

AO21x1_ASAP7_75t_L g1010 ( 
.A1(n_873),
.A2(n_80),
.B(n_81),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_909),
.B(n_854),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_803),
.B(n_766),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_802),
.A2(n_184),
.B(n_290),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_818),
.A2(n_179),
.B(n_288),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_875),
.A2(n_187),
.B(n_286),
.Y(n_1015)
);

BUFx4f_ASAP7_75t_L g1016 ( 
.A(n_877),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_855),
.A2(n_898),
.B(n_760),
.Y(n_1017)
);

NAND2x1_ASAP7_75t_L g1018 ( 
.A(n_840),
.B(n_124),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_766),
.A2(n_177),
.B(n_284),
.Y(n_1019)
);

AOI33xp33_ASAP7_75t_L g1020 ( 
.A1(n_863),
.A2(n_82),
.A3(n_84),
.B1(n_85),
.B2(n_87),
.B3(n_88),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_801),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_820),
.B(n_82),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_757),
.A2(n_194),
.B(n_283),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_846),
.A2(n_196),
.B(n_279),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_831),
.A2(n_89),
.B(n_90),
.C(n_91),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_774),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_SL g1027 ( 
.A(n_909),
.B(n_126),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_907),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_805),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_832),
.A2(n_92),
.B(n_93),
.C(n_94),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_770),
.A2(n_94),
.B(n_95),
.C(n_96),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_770),
.A2(n_205),
.B(n_278),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_781),
.B(n_95),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_803),
.B(n_98),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_781),
.B(n_99),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_877),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_807),
.B(n_103),
.Y(n_1037)
);

AOI33xp33_ASAP7_75t_L g1038 ( 
.A1(n_892),
.A2(n_104),
.A3(n_130),
.B1(n_133),
.B2(n_134),
.B3(n_135),
.Y(n_1038)
);

CKINVDCx10_ASAP7_75t_R g1039 ( 
.A(n_858),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_884),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_761),
.A2(n_140),
.B(n_146),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_841),
.B(n_151),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_848),
.A2(n_154),
.B(n_157),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_763),
.B(n_158),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_841),
.B(n_164),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_909),
.B(n_165),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_784),
.A2(n_166),
.B(n_167),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_848),
.A2(n_197),
.B(n_201),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_794),
.A2(n_799),
.B(n_806),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_885),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_883),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_800),
.A2(n_204),
.B(n_209),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_897),
.A2(n_210),
.B1(n_215),
.B2(n_216),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_908),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_892),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_896),
.B(n_231),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_902),
.B(n_241),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_888),
.A2(n_249),
.B(n_253),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_895),
.B(n_298),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_919),
.A2(n_864),
.B1(n_905),
.B2(n_894),
.Y(n_1060)
);

BUFx12f_ASAP7_75t_L g1061 ( 
.A(n_999),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_928),
.A2(n_882),
.B(n_876),
.Y(n_1062)
);

NAND2x1_ASAP7_75t_L g1063 ( 
.A(n_998),
.B(n_969),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_979),
.B(n_958),
.Y(n_1064)
);

NOR2x1_ASAP7_75t_SL g1065 ( 
.A(n_969),
.B(n_885),
.Y(n_1065)
);

CKINVDCx11_ASAP7_75t_R g1066 ( 
.A(n_922),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_966),
.A2(n_885),
.B(n_257),
.C(n_261),
.Y(n_1067)
);

AOI21xp33_ASAP7_75t_SL g1068 ( 
.A1(n_941),
.A2(n_917),
.B(n_939),
.Y(n_1068)
);

AOI221x1_ASAP7_75t_L g1069 ( 
.A1(n_1007),
.A2(n_1005),
.B1(n_948),
.B2(n_1015),
.C(n_986),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_960),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_925),
.A2(n_885),
.B(n_268),
.Y(n_1071)
);

INVx6_ASAP7_75t_L g1072 ( 
.A(n_982),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_977),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_956),
.B(n_276),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_L g1075 ( 
.A(n_941),
.B(n_277),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_910),
.A2(n_912),
.B(n_967),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_1018),
.A2(n_916),
.B(n_915),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_965),
.A2(n_913),
.B(n_963),
.Y(n_1078)
);

INVxp67_ASAP7_75t_SL g1079 ( 
.A(n_938),
.Y(n_1079)
);

OAI22x1_ASAP7_75t_L g1080 ( 
.A1(n_959),
.A2(n_1004),
.B1(n_956),
.B2(n_955),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_982),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1012),
.A2(n_952),
.B(n_932),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1029),
.B(n_931),
.Y(n_1083)
);

NOR2x1_ASAP7_75t_SL g1084 ( 
.A(n_982),
.B(n_1008),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_973),
.B(n_953),
.Y(n_1085)
);

AO21x1_ASAP7_75t_L g1086 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1002),
.B(n_1021),
.Y(n_1087)
);

AO21x1_ASAP7_75t_L g1088 ( 
.A1(n_1043),
.A2(n_1048),
.B(n_1027),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_1028),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_1025),
.A2(n_1030),
.B(n_1020),
.C(n_984),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_957),
.B(n_959),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_988),
.B(n_911),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_938),
.B(n_1027),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1035),
.B(n_936),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_938),
.Y(n_1095)
);

AOI21x1_ASAP7_75t_SL g1096 ( 
.A1(n_1056),
.A2(n_1042),
.B(n_1045),
.Y(n_1096)
);

O2A1O1Ixp5_ASAP7_75t_L g1097 ( 
.A1(n_1010),
.A2(n_1003),
.B(n_1011),
.C(n_1032),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1050),
.A2(n_992),
.B(n_1013),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_1016),
.Y(n_1099)
);

OA21x2_ASAP7_75t_L g1100 ( 
.A1(n_1019),
.A2(n_954),
.B(n_970),
.Y(n_1100)
);

AOI211x1_ASAP7_75t_L g1101 ( 
.A1(n_949),
.A2(n_950),
.B(n_944),
.C(n_946),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_1028),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_SL g1103 ( 
.A1(n_990),
.A2(n_995),
.B(n_945),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_SL g1104 ( 
.A(n_1016),
.B(n_995),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1040),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_972),
.A2(n_964),
.B(n_962),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1033),
.A2(n_934),
.B(n_942),
.C(n_1031),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_983),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_989),
.A2(n_1000),
.B(n_991),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_SL g1110 ( 
.A(n_996),
.B(n_1026),
.C(n_943),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_985),
.A2(n_994),
.B(n_1034),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_968),
.Y(n_1112)
);

CKINVDCx6p67_ASAP7_75t_R g1113 ( 
.A(n_1039),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_998),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1022),
.B(n_914),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1053),
.A2(n_1057),
.B(n_929),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_993),
.A2(n_997),
.B(n_1009),
.Y(n_1117)
);

OA21x2_ASAP7_75t_L g1118 ( 
.A1(n_954),
.A2(n_990),
.B(n_933),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1006),
.B(n_976),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1024),
.A2(n_1059),
.B(n_1052),
.Y(n_1120)
);

NAND2xp33_ASAP7_75t_L g1121 ( 
.A(n_927),
.B(n_975),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1038),
.A2(n_987),
.B(n_1037),
.C(n_1044),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1041),
.A2(n_1047),
.B(n_1014),
.C(n_1017),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1058),
.A2(n_1023),
.B(n_1049),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_935),
.B(n_940),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_961),
.B(n_951),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_924),
.B(n_921),
.Y(n_1127)
);

AOI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_1036),
.A2(n_1051),
.B1(n_1054),
.B2(n_974),
.C(n_1055),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1001),
.Y(n_1129)
);

BUFx2_ASAP7_75t_SL g1130 ( 
.A(n_941),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_982),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_947),
.A2(n_839),
.A3(n_815),
.B(n_1010),
.Y(n_1132)
);

OAI22x1_ASAP7_75t_L g1133 ( 
.A1(n_959),
.A2(n_795),
.B1(n_776),
.B2(n_765),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_919),
.B(n_920),
.Y(n_1134)
);

NAND2x1p5_ASAP7_75t_L g1135 ( 
.A(n_930),
.B(n_969),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_919),
.B(n_920),
.Y(n_1136)
);

AO32x2_ASAP7_75t_L g1137 ( 
.A1(n_1005),
.A2(n_981),
.A3(n_919),
.B1(n_980),
.B2(n_1053),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_919),
.B(n_920),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_919),
.A2(n_979),
.B1(n_978),
.B2(n_641),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_947),
.A2(n_926),
.B(n_928),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_919),
.B(n_920),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_920),
.Y(n_1142)
);

BUFx4_ASAP7_75t_SL g1143 ( 
.A(n_920),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_920),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_917),
.A2(n_765),
.B1(n_777),
.B2(n_773),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_919),
.B(n_920),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_947),
.A2(n_926),
.B(n_928),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_920),
.B(n_765),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_920),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_919),
.B(n_890),
.Y(n_1150)
);

AOI31xp67_ASAP7_75t_L g1151 ( 
.A1(n_1046),
.A2(n_645),
.A3(n_655),
.B(n_643),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_937),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_919),
.B(n_920),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_920),
.Y(n_1154)
);

AOI21xp33_ASAP7_75t_L g1155 ( 
.A1(n_919),
.A2(n_765),
.B(n_658),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_920),
.Y(n_1156)
);

AOI211x1_ASAP7_75t_L g1157 ( 
.A1(n_1003),
.A2(n_919),
.B(n_981),
.C(n_759),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_918),
.Y(n_1158)
);

AO21x2_ASAP7_75t_L g1159 ( 
.A1(n_947),
.A2(n_815),
.B(n_923),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_920),
.B(n_765),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_982),
.Y(n_1161)
);

OAI22x1_ASAP7_75t_L g1162 ( 
.A1(n_959),
.A2(n_795),
.B1(n_776),
.B2(n_765),
.Y(n_1162)
);

AOI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_919),
.A2(n_765),
.B(n_658),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_920),
.B(n_765),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_919),
.B(n_920),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_947),
.A2(n_926),
.B(n_928),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_918),
.Y(n_1167)
);

AOI21xp33_ASAP7_75t_L g1168 ( 
.A1(n_919),
.A2(n_765),
.B(n_658),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_920),
.B(n_765),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_920),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_919),
.B(n_920),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_920),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_947),
.A2(n_926),
.B(n_928),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_919),
.B(n_920),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_919),
.B(n_890),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_947),
.A2(n_926),
.B(n_928),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_920),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_920),
.B(n_765),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_920),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_920),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_920),
.Y(n_1181)
);

INVx6_ASAP7_75t_SL g1182 ( 
.A(n_959),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_925),
.A2(n_815),
.B(n_839),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_919),
.B(n_920),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_947),
.A2(n_926),
.B(n_928),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_919),
.B(n_920),
.Y(n_1186)
);

AOI221xp5_ASAP7_75t_SL g1187 ( 
.A1(n_980),
.A2(n_759),
.B1(n_931),
.B2(n_973),
.C(n_971),
.Y(n_1187)
);

CKINVDCx11_ASAP7_75t_R g1188 ( 
.A(n_922),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_999),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_919),
.B(n_920),
.Y(n_1190)
);

BUFx10_ASAP7_75t_L g1191 ( 
.A(n_955),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_920),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_919),
.B(n_920),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_947),
.A2(n_926),
.B(n_928),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_920),
.B(n_765),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_919),
.B(n_920),
.Y(n_1196)
);

OAI21xp33_ASAP7_75t_L g1197 ( 
.A1(n_952),
.A2(n_765),
.B(n_680),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_SL g1198 ( 
.A1(n_948),
.A2(n_1015),
.B(n_1043),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_920),
.B(n_765),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_920),
.B(n_765),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_919),
.B(n_920),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_919),
.B(n_920),
.Y(n_1202)
);

NOR2x1_ASAP7_75t_SL g1203 ( 
.A(n_930),
.B(n_886),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_919),
.B(n_920),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_919),
.B(n_920),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1079),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1070),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1133),
.A2(n_1162),
.B1(n_1182),
.B2(n_1175),
.Y(n_1208)
);

INVx6_ASAP7_75t_L g1209 ( 
.A(n_1191),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1107),
.A2(n_1175),
.B(n_1150),
.C(n_1082),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1197),
.B(n_1145),
.Y(n_1211)
);

OAI22x1_ASAP7_75t_L g1212 ( 
.A1(n_1160),
.A2(n_1169),
.B1(n_1156),
.B2(n_1149),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1114),
.B(n_1160),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1182),
.B(n_1108),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1087),
.A2(n_1169),
.B1(n_1178),
.B2(n_1164),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1150),
.A2(n_1080),
.B1(n_1163),
.B2(n_1155),
.Y(n_1216)
);

INVx8_ASAP7_75t_L g1217 ( 
.A(n_1131),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1064),
.B(n_1157),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1143),
.Y(n_1219)
);

AO21x2_ASAP7_75t_L g1220 ( 
.A1(n_1198),
.A2(n_1147),
.B(n_1140),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_1063),
.B(n_1130),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1152),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1144),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1143),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1107),
.A2(n_1082),
.B(n_1111),
.C(n_1106),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1065),
.A2(n_1084),
.B(n_1088),
.Y(n_1226)
);

BUFx8_ASAP7_75t_L g1227 ( 
.A(n_1170),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1179),
.B(n_1148),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_SL g1229 ( 
.A1(n_1203),
.A2(n_1103),
.B(n_1086),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1205),
.A2(n_1204),
.B1(n_1202),
.B2(n_1201),
.Y(n_1230)
);

BUFx2_ASAP7_75t_R g1231 ( 
.A(n_1134),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1168),
.A2(n_1171),
.B1(n_1136),
.B2(n_1138),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1106),
.A2(n_1117),
.B(n_1111),
.C(n_1097),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1166),
.A2(n_1185),
.A3(n_1173),
.B(n_1194),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1195),
.B(n_1199),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1141),
.A2(n_1193),
.B1(n_1184),
.B2(n_1146),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1076),
.A2(n_1078),
.B(n_1077),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1153),
.A2(n_1165),
.B1(n_1190),
.B2(n_1196),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_1144),
.Y(n_1239)
);

BUFx4f_ASAP7_75t_SL g1240 ( 
.A(n_1113),
.Y(n_1240)
);

NOR2xp67_ASAP7_75t_L g1241 ( 
.A(n_1142),
.B(n_1177),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1200),
.B(n_1154),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1191),
.B(n_1068),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1176),
.A2(n_1194),
.A3(n_1129),
.B(n_1069),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1174),
.B(n_1186),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1154),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_SL g1247 ( 
.A1(n_1067),
.A2(n_1122),
.B(n_1090),
.C(n_1094),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1091),
.A2(n_1083),
.B1(n_1189),
.B2(n_1061),
.Y(n_1248)
);

BUFx10_ASAP7_75t_L g1249 ( 
.A(n_1181),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1096),
.A2(n_1098),
.B(n_1071),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1172),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1066),
.Y(n_1252)
);

OAI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1104),
.A2(n_1115),
.B1(n_1074),
.B2(n_1180),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1180),
.A2(n_1192),
.B1(n_1073),
.B2(n_1099),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1062),
.A2(n_1120),
.B(n_1124),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1085),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1109),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1101),
.A2(n_1112),
.B1(n_1060),
.B2(n_1116),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1110),
.A2(n_1119),
.B1(n_1128),
.B2(n_1121),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_1066),
.Y(n_1260)
);

AOI221xp5_ASAP7_75t_L g1261 ( 
.A1(n_1110),
.A2(n_1128),
.B1(n_1127),
.B2(n_1126),
.C(n_1125),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1099),
.B(n_1135),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1123),
.A2(n_1125),
.A3(n_1132),
.B(n_1159),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1183),
.A2(n_1100),
.B(n_1118),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1161),
.A2(n_1075),
.B1(n_1072),
.B2(n_1081),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1188),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1137),
.B(n_1102),
.Y(n_1267)
);

CKINVDCx9p33_ASAP7_75t_R g1268 ( 
.A(n_1188),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1132),
.A2(n_1151),
.A3(n_1137),
.B(n_1100),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1089),
.Y(n_1270)
);

AOI31xp67_ASAP7_75t_L g1271 ( 
.A1(n_1137),
.A2(n_1093),
.A3(n_1167),
.B(n_1158),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1092),
.B(n_919),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1092),
.B(n_919),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1079),
.B(n_1095),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1133),
.A2(n_785),
.B1(n_1162),
.B2(n_959),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_SL g1276 ( 
.A1(n_1065),
.A2(n_1084),
.B(n_1088),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1179),
.B(n_765),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1086),
.A2(n_1088),
.A3(n_1147),
.B(n_1140),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1134),
.A2(n_1138),
.B1(n_1141),
.B2(n_1136),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_1066),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1092),
.B(n_919),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1079),
.Y(n_1282)
);

AO21x2_ASAP7_75t_L g1283 ( 
.A1(n_1198),
.A2(n_1147),
.B(n_1140),
.Y(n_1283)
);

NOR3xp33_ASAP7_75t_L g1284 ( 
.A(n_1155),
.B(n_1168),
.C(n_1163),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1079),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1197),
.A2(n_765),
.B1(n_773),
.B2(n_769),
.Y(n_1286)
);

AOI21xp33_ASAP7_75t_L g1287 ( 
.A1(n_1080),
.A2(n_1187),
.B(n_1139),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1107),
.A2(n_971),
.B(n_1175),
.C(n_1150),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1087),
.B(n_920),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1087),
.B(n_920),
.Y(n_1290)
);

AOI21xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1133),
.A2(n_773),
.B(n_769),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1105),
.Y(n_1292)
);

OAI21xp33_ASAP7_75t_L g1293 ( 
.A1(n_1211),
.A2(n_1275),
.B(n_1216),
.Y(n_1293)
);

AO21x1_ASAP7_75t_SL g1294 ( 
.A1(n_1206),
.A2(n_1285),
.B(n_1282),
.Y(n_1294)
);

AOI221xp5_ASAP7_75t_L g1295 ( 
.A1(n_1291),
.A2(n_1279),
.B1(n_1287),
.B2(n_1261),
.C(n_1288),
.Y(n_1295)
);

INVxp33_ASAP7_75t_L g1296 ( 
.A(n_1277),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1270),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1207),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1222),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1257),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1233),
.A2(n_1225),
.B(n_1247),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1261),
.A2(n_1259),
.B1(n_1273),
.B2(n_1272),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1223),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1250),
.A2(n_1237),
.B(n_1255),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1282),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1289),
.B(n_1290),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_1251),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1219),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1272),
.A2(n_1273),
.B1(n_1281),
.B2(n_1230),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1228),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1209),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1242),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1209),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1209),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1256),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1217),
.Y(n_1316)
);

NAND2x1_ASAP7_75t_L g1317 ( 
.A(n_1226),
.B(n_1276),
.Y(n_1317)
);

OAI211xp5_ASAP7_75t_L g1318 ( 
.A1(n_1208),
.A2(n_1248),
.B(n_1286),
.C(n_1254),
.Y(n_1318)
);

OR2x6_ASAP7_75t_L g1319 ( 
.A(n_1221),
.B(n_1274),
.Y(n_1319)
);

INVx5_ASAP7_75t_L g1320 ( 
.A(n_1221),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1267),
.Y(n_1321)
);

CKINVDCx6p67_ASAP7_75t_R g1322 ( 
.A(n_1268),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1230),
.A2(n_1236),
.B1(n_1279),
.B2(n_1245),
.Y(n_1323)
);

BUFx4f_ASAP7_75t_SL g1324 ( 
.A(n_1280),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1234),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1218),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1234),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1245),
.B(n_1238),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1249),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1292),
.B(n_1236),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1271),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1218),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1249),
.Y(n_1333)
);

NOR2x1p5_ASAP7_75t_L g1334 ( 
.A(n_1224),
.B(n_1252),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1253),
.A2(n_1235),
.B1(n_1284),
.B2(n_1232),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1239),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1220),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1246),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1253),
.A2(n_1254),
.B1(n_1227),
.B2(n_1213),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1300),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1321),
.B(n_1263),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1321),
.B(n_1263),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1309),
.B(n_1210),
.Y(n_1343)
);

BUFx4f_ASAP7_75t_SL g1344 ( 
.A(n_1322),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1320),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1325),
.B(n_1283),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1337),
.B(n_1283),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1327),
.B(n_1220),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_1294),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1318),
.A2(n_1258),
.B1(n_1213),
.B2(n_1229),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1330),
.B(n_1278),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1328),
.B(n_1305),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1330),
.B(n_1278),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1331),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1303),
.Y(n_1355)
);

NOR2x1_ASAP7_75t_L g1356 ( 
.A(n_1319),
.B(n_1317),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1328),
.B(n_1244),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1326),
.B(n_1332),
.Y(n_1358)
);

INVxp33_ASAP7_75t_L g1359 ( 
.A(n_1355),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1340),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1340),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1351),
.B(n_1244),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1355),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1349),
.B(n_1319),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1349),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1353),
.B(n_1264),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1352),
.B(n_1312),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1352),
.B(n_1323),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1341),
.B(n_1269),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1341),
.B(n_1269),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1358),
.B(n_1341),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1354),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1345),
.B(n_1320),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1347),
.B(n_1304),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1342),
.B(n_1294),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1362),
.B(n_1342),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1363),
.B(n_1358),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1360),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1362),
.B(n_1346),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1359),
.B(n_1344),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1374),
.B(n_1346),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1372),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1371),
.B(n_1357),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1365),
.B(n_1320),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1371),
.B(n_1357),
.Y(n_1385)
);

NAND4xp25_ASAP7_75t_L g1386 ( 
.A(n_1368),
.B(n_1339),
.C(n_1335),
.D(n_1295),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1361),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1366),
.B(n_1348),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1366),
.B(n_1348),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1365),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1366),
.B(n_1348),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1375),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1388),
.B(n_1389),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1388),
.B(n_1369),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1389),
.B(n_1369),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1378),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1391),
.B(n_1369),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1387),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1387),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1390),
.Y(n_1400)
);

OAI21xp33_ASAP7_75t_L g1401 ( 
.A1(n_1392),
.A2(n_1375),
.B(n_1293),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1376),
.B(n_1367),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1376),
.B(n_1392),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1379),
.B(n_1370),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1382),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1405),
.Y(n_1406)
);

OAI21xp33_ASAP7_75t_L g1407 ( 
.A1(n_1401),
.A2(n_1386),
.B(n_1390),
.Y(n_1407)
);

OAI21xp33_ASAP7_75t_L g1408 ( 
.A1(n_1403),
.A2(n_1386),
.B(n_1390),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1396),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1403),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1400),
.Y(n_1411)
);

OAI222xp33_ASAP7_75t_L g1412 ( 
.A1(n_1402),
.A2(n_1364),
.B1(n_1384),
.B2(n_1375),
.C1(n_1383),
.C2(n_1368),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1396),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1398),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1402),
.B(n_1383),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1405),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1393),
.B(n_1344),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1398),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1404),
.B(n_1381),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1404),
.B(n_1379),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1400),
.B(n_1380),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1399),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1399),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1400),
.A2(n_1381),
.B1(n_1364),
.B2(n_1343),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1421),
.B(n_1381),
.Y(n_1425)
);

NAND2x1_ASAP7_75t_L g1426 ( 
.A(n_1411),
.B(n_1364),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_R g1427 ( 
.A(n_1417),
.B(n_1240),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1415),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1412),
.A2(n_1297),
.B(n_1356),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1419),
.B(n_1393),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1410),
.B(n_1394),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1407),
.A2(n_1381),
.B1(n_1377),
.B2(n_1385),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1408),
.A2(n_1364),
.B(n_1373),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1411),
.A2(n_1356),
.B(n_1350),
.Y(n_1434)
);

AOI211xp5_ASAP7_75t_L g1435 ( 
.A1(n_1433),
.A2(n_1297),
.B(n_1343),
.C(n_1415),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_SL g1436 ( 
.A1(n_1429),
.A2(n_1420),
.B(n_1345),
.C(n_1333),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1425),
.B(n_1419),
.Y(n_1437)
);

AOI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1428),
.A2(n_1424),
.B1(n_1423),
.B2(n_1422),
.C(n_1413),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1431),
.B(n_1322),
.Y(n_1439)
);

AOI221xp5_ASAP7_75t_L g1440 ( 
.A1(n_1434),
.A2(n_1423),
.B1(n_1422),
.B2(n_1418),
.C(n_1409),
.Y(n_1440)
);

OAI321xp33_ASAP7_75t_L g1441 ( 
.A1(n_1432),
.A2(n_1364),
.A3(n_1385),
.B1(n_1297),
.B2(n_1413),
.C(n_1409),
.Y(n_1441)
);

NOR3xp33_ASAP7_75t_L g1442 ( 
.A(n_1426),
.B(n_1266),
.C(n_1260),
.Y(n_1442)
);

OAI211xp5_ASAP7_75t_L g1443 ( 
.A1(n_1427),
.A2(n_1350),
.B(n_1297),
.C(n_1302),
.Y(n_1443)
);

NAND3xp33_ASAP7_75t_L g1444 ( 
.A(n_1425),
.B(n_1227),
.C(n_1414),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1430),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1428),
.B(n_1414),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1439),
.B(n_1324),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1442),
.B(n_1308),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1436),
.A2(n_1329),
.B(n_1243),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1437),
.B(n_1394),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1445),
.B(n_1395),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1443),
.B(n_1307),
.C(n_1297),
.Y(n_1452)
);

NOR4xp25_ASAP7_75t_L g1453 ( 
.A(n_1441),
.B(n_1315),
.C(n_1298),
.D(n_1299),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1438),
.B(n_1418),
.Y(n_1454)
);

AOI211xp5_ASAP7_75t_L g1455 ( 
.A1(n_1453),
.A2(n_1435),
.B(n_1444),
.C(n_1440),
.Y(n_1455)
);

NAND3xp33_ASAP7_75t_L g1456 ( 
.A(n_1452),
.B(n_1446),
.C(n_1308),
.Y(n_1456)
);

AOI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1454),
.A2(n_1334),
.B1(n_1364),
.B2(n_1416),
.Y(n_1457)
);

NOR2x1_ASAP7_75t_L g1458 ( 
.A(n_1448),
.B(n_1221),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1451),
.B(n_1395),
.Y(n_1459)
);

NOR3xp33_ASAP7_75t_L g1460 ( 
.A(n_1449),
.B(n_1313),
.C(n_1311),
.Y(n_1460)
);

AND4x2_ASAP7_75t_L g1461 ( 
.A(n_1447),
.B(n_1356),
.C(n_1231),
.D(n_1301),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_SL g1462 ( 
.A(n_1450),
.B(n_1320),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_L g1463 ( 
.A(n_1456),
.B(n_1241),
.Y(n_1463)
);

NOR2x1_ASAP7_75t_L g1464 ( 
.A(n_1458),
.B(n_1214),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_L g1465 ( 
.A(n_1461),
.B(n_1262),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1457),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1462),
.B(n_1296),
.Y(n_1467)
);

NOR2x1_ASAP7_75t_L g1468 ( 
.A(n_1459),
.B(n_1265),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1455),
.B(n_1406),
.Y(n_1469)
);

NOR3xp33_ASAP7_75t_L g1470 ( 
.A(n_1465),
.B(n_1460),
.C(n_1313),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1469),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1466),
.B(n_1397),
.Y(n_1472)
);

AOI21xp33_ASAP7_75t_L g1473 ( 
.A1(n_1463),
.A2(n_1296),
.B(n_1311),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1471),
.B(n_1464),
.C(n_1467),
.Y(n_1474)
);

OAI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1470),
.A2(n_1473),
.B1(n_1472),
.B2(n_1468),
.C(n_1314),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1474),
.B(n_1406),
.Y(n_1476)
);

OAI21xp33_ASAP7_75t_L g1477 ( 
.A1(n_1476),
.A2(n_1475),
.B(n_1314),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1477),
.A2(n_1215),
.B(n_1310),
.Y(n_1478)
);

XNOR2x1_ASAP7_75t_L g1479 ( 
.A(n_1478),
.B(n_1212),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1479),
.A2(n_1306),
.B(n_1338),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1480),
.B(n_1316),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1481),
.A2(n_1480),
.B1(n_1416),
.B2(n_1336),
.Y(n_1482)
);


endmodule