module fake_jpeg_24962_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_5),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_34),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_2),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_17),
.A2(n_4),
.B1(n_7),
.B2(n_9),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_23),
.Y(n_39)
);

HAxp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_9),
.CON(n_33),
.SN(n_33)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_10),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_48),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_27),
.B1(n_31),
.B2(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_19),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_12),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_40),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_54),
.B1(n_57),
.B2(n_55),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_34),
.C(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_60),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_34),
.B1(n_16),
.B2(n_23),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_64),
.B1(n_56),
.B2(n_58),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_59),
.B(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_34),
.B1(n_18),
.B2(n_20),
.Y(n_57)
);

AO21x1_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_12),
.B(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_41),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_40),
.B1(n_37),
.B2(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_67),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_47),
.B(n_51),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_76),
.B(n_71),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_61),
.B1(n_59),
.B2(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_76),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_81),
.A2(n_84),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_67),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_89),
.C(n_90),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_74),
.C(n_77),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_97),
.Y(n_99)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_90),
.B(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

OAI321xp33_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_69),
.A3(n_73),
.B1(n_80),
.B2(n_82),
.C(n_94),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_98),
.B(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_99),
.Y(n_102)
);


endmodule