module fake_netlist_1_3646_n_443 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_12, n_9, n_17, n_14, n_10, n_15, n_42, n_24, n_19, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_443);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_443;
wire n_117;
wire n_361;
wire n_185;
wire n_57;
wire n_407;
wire n_284;
wire n_278;
wire n_60;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_73;
wire n_97;
wire n_167;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_59;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_61;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_69;
wire n_204;
wire n_430;
wire n_88;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_56;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_58;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_55;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g55 ( .A(n_36), .Y(n_55) );
INVx1_ASAP7_75t_L g56 ( .A(n_26), .Y(n_56) );
INVx1_ASAP7_75t_L g57 ( .A(n_25), .Y(n_57) );
CKINVDCx16_ASAP7_75t_R g58 ( .A(n_44), .Y(n_58) );
BUFx6f_ASAP7_75t_L g59 ( .A(n_53), .Y(n_59) );
INVx1_ASAP7_75t_L g60 ( .A(n_49), .Y(n_60) );
INVx1_ASAP7_75t_L g61 ( .A(n_43), .Y(n_61) );
INVx1_ASAP7_75t_L g62 ( .A(n_24), .Y(n_62) );
CKINVDCx5p33_ASAP7_75t_R g63 ( .A(n_27), .Y(n_63) );
INVxp33_ASAP7_75t_SL g64 ( .A(n_0), .Y(n_64) );
INVxp67_ASAP7_75t_L g65 ( .A(n_47), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_14), .Y(n_66) );
INVx1_ASAP7_75t_L g67 ( .A(n_13), .Y(n_67) );
INVxp67_ASAP7_75t_SL g68 ( .A(n_52), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_38), .Y(n_69) );
INVxp33_ASAP7_75t_SL g70 ( .A(n_50), .Y(n_70) );
CKINVDCx5p33_ASAP7_75t_R g71 ( .A(n_51), .Y(n_71) );
INVxp67_ASAP7_75t_SL g72 ( .A(n_39), .Y(n_72) );
INVxp67_ASAP7_75t_L g73 ( .A(n_35), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_17), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_46), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_48), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_2), .Y(n_77) );
INVx1_ASAP7_75t_SL g78 ( .A(n_37), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_5), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_17), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_45), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_2), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_21), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_11), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_13), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_4), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_32), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_33), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_40), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_6), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_41), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_29), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_18), .Y(n_93) );
INVx3_ASAP7_75t_L g94 ( .A(n_61), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_61), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_90), .Y(n_96) );
INVx3_ASAP7_75t_L g97 ( .A(n_62), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_90), .Y(n_98) );
NAND2xp5_ASAP7_75t_L g99 ( .A(n_66), .B(n_0), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_62), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_92), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_92), .Y(n_102) );
BUFx2_ASAP7_75t_L g103 ( .A(n_58), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_59), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g105 ( .A1(n_79), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_59), .Y(n_106) );
INVx4_ASAP7_75t_L g107 ( .A(n_59), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_66), .B(n_1), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_59), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_67), .B(n_3), .Y(n_110) );
INVx3_ASAP7_75t_L g111 ( .A(n_59), .Y(n_111) );
AND2x4_ASAP7_75t_L g112 ( .A(n_55), .B(n_5), .Y(n_112) );
NAND2xp33_ASAP7_75t_L g113 ( .A(n_63), .B(n_34), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_56), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_57), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_112), .B(n_74), .Y(n_116) );
AND2x4_ASAP7_75t_L g117 ( .A(n_112), .B(n_80), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_96), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_96), .B(n_63), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_98), .B(n_71), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_94), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_94), .Y(n_122) );
BUFx4f_ASAP7_75t_L g123 ( .A(n_112), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_111), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_112), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_94), .Y(n_126) );
BUFx10_ASAP7_75t_L g127 ( .A(n_112), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_103), .B(n_71), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_98), .B(n_65), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_107), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_94), .Y(n_131) );
INVx2_ASAP7_75t_SL g132 ( .A(n_95), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_94), .Y(n_133) );
NAND3x1_ASAP7_75t_L g134 ( .A(n_99), .B(n_60), .C(n_91), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_104), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_97), .B(n_95), .Y(n_136) );
INVx1_ASAP7_75t_SL g137 ( .A(n_103), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_111), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_97), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_137), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_118), .B(n_114), .Y(n_141) );
BUFx4f_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_121), .Y(n_143) );
BUFx4f_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_136), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_136), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_121), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_127), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_122), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_119), .B(n_100), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_136), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_132), .B(n_97), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_122), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
NOR2x2_ASAP7_75t_L g155 ( .A(n_137), .B(n_77), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_128), .B(n_114), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_123), .Y(n_157) );
INVxp67_ASAP7_75t_SL g158 ( .A(n_125), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_119), .B(n_100), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_131), .Y(n_161) );
AOI22xp5_ASAP7_75t_SL g162 ( .A1(n_119), .A2(n_77), .B1(n_93), .B2(n_105), .Y(n_162) );
NOR2x1_ASAP7_75t_L g163 ( .A(n_116), .B(n_113), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_133), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_120), .B(n_101), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_127), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_145), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_141), .A2(n_123), .B1(n_125), .B2(n_120), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_154), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_159), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
INVx1_ASAP7_75t_SL g178 ( .A(n_159), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_160), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_157), .B(n_116), .Y(n_180) );
AOI22xp33_ASAP7_75t_SL g181 ( .A1(n_162), .A2(n_105), .B1(n_64), .B2(n_93), .Y(n_181) );
NOR2xp33_ASAP7_75t_SL g182 ( .A(n_157), .B(n_127), .Y(n_182) );
BUFx2_ASAP7_75t_SL g183 ( .A(n_157), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_161), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_161), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_141), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_162), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_143), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_141), .B(n_123), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_143), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_164), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_141), .B(n_132), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_150), .A2(n_125), .B1(n_117), .B2(n_116), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_167), .B(n_127), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
NAND2xp33_ASAP7_75t_L g196 ( .A(n_169), .B(n_132), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
INVxp67_ASAP7_75t_SL g198 ( .A(n_142), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_170), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_181), .A2(n_146), .B1(n_145), .B2(n_144), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_173), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_176), .B(n_156), .Y(n_203) );
OAI22xp33_ASAP7_75t_L g204 ( .A1(n_187), .A2(n_155), .B1(n_142), .B2(n_144), .Y(n_204) );
OR2x6_ASAP7_75t_L g205 ( .A(n_183), .B(n_157), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_186), .A2(n_142), .B1(n_144), .B2(n_166), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_173), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_198), .B(n_166), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_170), .Y(n_209) );
AOI22x1_ASAP7_75t_L g210 ( .A1(n_173), .A2(n_104), .B1(n_109), .B2(n_106), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_186), .A2(n_166), .B1(n_144), .B2(n_163), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_174), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_174), .Y(n_213) );
OAI221xp5_ASAP7_75t_L g214 ( .A1(n_181), .A2(n_129), .B1(n_151), .B2(n_166), .C(n_110), .Y(n_214) );
OAI221xp5_ASAP7_75t_L g215 ( .A1(n_178), .A2(n_129), .B1(n_151), .B2(n_110), .C(n_158), .Y(n_215) );
O2A1O1Ixp5_ASAP7_75t_SL g216 ( .A1(n_175), .A2(n_89), .B(n_75), .C(n_76), .Y(n_216) );
OAI22xp33_ASAP7_75t_L g217 ( .A1(n_178), .A2(n_64), .B1(n_145), .B2(n_146), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_175), .Y(n_218) );
OAI22xp33_ASAP7_75t_L g219 ( .A1(n_193), .A2(n_146), .B1(n_145), .B2(n_108), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_188), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_188), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_188), .Y(n_222) );
NOR2xp67_ASAP7_75t_SL g223 ( .A(n_183), .B(n_148), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_189), .A2(n_180), .B1(n_194), .B2(n_145), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_202), .B(n_189), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_214), .A2(n_193), .B1(n_192), .B2(n_172), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_205), .B(n_198), .Y(n_227) );
OAI211xp5_ASAP7_75t_L g228 ( .A1(n_201), .A2(n_99), .B(n_108), .C(n_86), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_202), .Y(n_229) );
AOI32xp33_ASAP7_75t_L g230 ( .A1(n_204), .A2(n_194), .A3(n_84), .B1(n_85), .B2(n_82), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_207), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_212), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_219), .A2(n_192), .B1(n_177), .B2(n_184), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_207), .A2(n_196), .B(n_190), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_220), .B(n_190), .Y(n_235) );
AOI221xp5_ASAP7_75t_L g236 ( .A1(n_215), .A2(n_101), .B1(n_102), .B2(n_117), .C(n_116), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g237 ( .A1(n_200), .A2(n_182), .B1(n_185), .B2(n_184), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_220), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_221), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_212), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_217), .A2(n_134), .B1(n_199), .B2(n_185), .Y(n_241) );
AOI21x1_ASAP7_75t_L g242 ( .A1(n_223), .A2(n_199), .B(n_177), .Y(n_242) );
AOI22x1_ASAP7_75t_SL g243 ( .A1(n_209), .A2(n_88), .B1(n_68), .B2(n_72), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_226), .A2(n_213), .B1(n_218), .B2(n_221), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_239), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_239), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_227), .B(n_222), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_239), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_232), .B(n_213), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_236), .A2(n_208), .B1(n_224), .B2(n_203), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_227), .Y(n_251) );
OAI31xp33_ASAP7_75t_L g252 ( .A1(n_228), .A2(n_206), .A3(n_208), .B(n_218), .Y(n_252) );
AO22x1_ASAP7_75t_L g253 ( .A1(n_227), .A2(n_208), .B1(n_222), .B2(n_70), .Y(n_253) );
OAI221xp5_ASAP7_75t_L g254 ( .A1(n_230), .A2(n_211), .B1(n_205), .B2(n_102), .C(n_182), .Y(n_254) );
AOI33xp33_ASAP7_75t_L g255 ( .A1(n_232), .A2(n_69), .A3(n_87), .B1(n_81), .B2(n_83), .B3(n_117), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_233), .A2(n_216), .B(n_134), .Y(n_256) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_242), .A2(n_210), .B(n_191), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_239), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_240), .Y(n_259) );
OA222x2_ASAP7_75t_L g260 ( .A1(n_240), .A2(n_205), .B1(n_191), .B2(n_179), .C1(n_195), .C2(n_190), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_229), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_235), .B(n_195), .Y(n_263) );
AOI22xp33_ASAP7_75t_SL g264 ( .A1(n_243), .A2(n_205), .B1(n_179), .B2(n_180), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_259), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_259), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_249), .B(n_262), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_249), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_263), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_249), .Y(n_270) );
INVx8_ASAP7_75t_L g271 ( .A(n_247), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_263), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_263), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g274 ( .A(n_264), .B(n_216), .C(n_243), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_251), .B(n_239), .Y(n_275) );
AOI211xp5_ASAP7_75t_L g276 ( .A1(n_253), .A2(n_237), .B(n_113), .C(n_241), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_247), .B(n_225), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_262), .Y(n_278) );
OAI31xp33_ASAP7_75t_L g279 ( .A1(n_254), .A2(n_225), .A3(n_180), .B(n_235), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_261), .Y(n_280) );
OAI211xp5_ASAP7_75t_SL g281 ( .A1(n_255), .A2(n_252), .B(n_250), .C(n_73), .Y(n_281) );
OAI211xp5_ASAP7_75t_L g282 ( .A1(n_252), .A2(n_88), .B(n_97), .C(n_115), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_254), .A2(n_238), .B1(n_231), .B2(n_134), .Y(n_283) );
OAI211xp5_ASAP7_75t_SL g284 ( .A1(n_244), .A2(n_115), .B(n_97), .C(n_78), .Y(n_284) );
NAND4xp25_ASAP7_75t_L g285 ( .A(n_244), .B(n_115), .C(n_117), .D(n_107), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_251), .B(n_231), .Y(n_286) );
OAI33xp33_ASAP7_75t_L g287 ( .A1(n_260), .A2(n_106), .A3(n_109), .B1(n_8), .B2(n_9), .B3(n_10), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_251), .B(n_238), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_261), .B(n_195), .Y(n_289) );
NOR3xp33_ASAP7_75t_SL g290 ( .A(n_256), .B(n_234), .C(n_152), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_271), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_265), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_266), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_267), .B(n_261), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_269), .B(n_247), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_268), .B(n_247), .Y(n_296) );
OAI21xp5_ASAP7_75t_SL g297 ( .A1(n_279), .A2(n_256), .B(n_247), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_278), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_271), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_272), .B(n_245), .Y(n_300) );
AOI332xp33_ASAP7_75t_L g301 ( .A1(n_270), .A2(n_115), .A3(n_111), .B1(n_11), .B2(n_12), .B3(n_14), .C1(n_15), .C2(n_16), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_273), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_288), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_277), .B(n_253), .Y(n_304) );
INVxp33_ASAP7_75t_L g305 ( .A(n_286), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_280), .B(n_245), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_289), .B(n_271), .Y(n_307) );
NAND2x1_ASAP7_75t_SL g308 ( .A(n_286), .B(n_246), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_275), .B(n_246), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_275), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_290), .B(n_246), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_283), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_279), .B(n_246), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_276), .B(n_248), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_274), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_285), .B(n_248), .Y(n_316) );
OAI211xp5_ASAP7_75t_SL g317 ( .A1(n_276), .A2(n_139), .B(n_124), .C(n_138), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_274), .B(n_258), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_282), .B(n_258), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_287), .B(n_258), .Y(n_320) );
NAND3xp33_ASAP7_75t_L g321 ( .A(n_281), .B(n_104), .C(n_107), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_284), .B(n_258), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_265), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_281), .B(n_6), .Y(n_324) );
OR2x6_ASAP7_75t_L g325 ( .A(n_271), .B(n_258), .Y(n_325) );
NAND4xp75_ASAP7_75t_L g326 ( .A(n_279), .B(n_257), .C(n_12), .D(n_7), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_265), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_267), .B(n_258), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_298), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_291), .B(n_19), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_292), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_295), .B(n_257), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_293), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_303), .B(n_257), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_294), .B(n_104), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_315), .B(n_242), .Y(n_336) );
NOR2xp33_ASAP7_75t_R g337 ( .A(n_299), .B(n_20), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_323), .Y(n_338) );
NAND2xp33_ASAP7_75t_SL g339 ( .A(n_305), .B(n_223), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_314), .B(n_104), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_327), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_308), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_302), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_300), .B(n_197), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_294), .B(n_22), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_296), .Y(n_346) );
NOR2xp33_ASAP7_75t_SL g347 ( .A(n_326), .B(n_171), .Y(n_347) );
NAND2xp33_ASAP7_75t_SL g348 ( .A(n_305), .B(n_171), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_304), .B(n_23), .Y(n_349) );
INVxp67_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_310), .B(n_28), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_325), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_307), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_328), .B(n_30), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_311), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_328), .B(n_309), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_306), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_306), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_311), .Y(n_360) );
NAND2xp33_ASAP7_75t_SL g361 ( .A(n_313), .B(n_171), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_325), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_312), .B(n_31), .Y(n_363) );
OAI31xp33_ASAP7_75t_L g364 ( .A1(n_324), .A2(n_153), .A3(n_168), .B(n_165), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_335), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_355), .A2(n_324), .B1(n_297), .B2(n_313), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_358), .Y(n_367) );
OAI211xp5_ASAP7_75t_SL g368 ( .A1(n_364), .A2(n_316), .B(n_301), .C(n_321), .Y(n_368) );
XNOR2xp5_ASAP7_75t_L g369 ( .A(n_360), .B(n_309), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_346), .B(n_312), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_331), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_335), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_359), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_357), .B(n_318), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_350), .B(n_322), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_339), .B(n_319), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_338), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_341), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_329), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_329), .Y(n_381) );
INVxp67_ASAP7_75t_L g382 ( .A(n_340), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_343), .Y(n_383) );
OAI21xp33_ASAP7_75t_L g384 ( .A1(n_356), .A2(n_317), .B(n_210), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_337), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_339), .A2(n_171), .B1(n_135), .B2(n_146), .C(n_153), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_334), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_362), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_362), .Y(n_389) );
XOR2x2_ASAP7_75t_L g390 ( .A(n_330), .B(n_42), .Y(n_390) );
AOI32xp33_ASAP7_75t_L g391 ( .A1(n_361), .A2(n_148), .A3(n_147), .B1(n_149), .B2(n_153), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_345), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_349), .B(n_352), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_345), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_348), .B(n_135), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_332), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_332), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_352), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_342), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_344), .Y(n_400) );
XNOR2xp5_ASAP7_75t_L g401 ( .A(n_354), .B(n_54), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_351), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_348), .Y(n_403) );
XNOR2xp5_ASAP7_75t_L g404 ( .A(n_363), .B(n_148), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_336), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_347), .Y(n_406) );
AOI211xp5_ASAP7_75t_L g407 ( .A1(n_337), .A2(n_169), .B(n_148), .C(n_130), .Y(n_407) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_335), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_353), .Y(n_409) );
OAI21xp5_ASAP7_75t_SL g410 ( .A1(n_362), .A2(n_264), .B(n_291), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_337), .A2(n_362), .B1(n_291), .B2(n_299), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_411), .A2(n_385), .B1(n_410), .B2(n_366), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_367), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_377), .A2(n_408), .B1(n_409), .B2(n_396), .Y(n_414) );
NOR2x1p5_ASAP7_75t_L g415 ( .A(n_408), .B(n_399), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_L g416 ( .A1(n_407), .A2(n_377), .B(n_396), .C(n_391), .Y(n_416) );
XNOR2xp5_ASAP7_75t_L g417 ( .A(n_390), .B(n_369), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_373), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_375), .A2(n_382), .B1(n_393), .B2(n_400), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_368), .A2(n_389), .B1(n_388), .B2(n_373), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_376), .A2(n_379), .B1(n_371), .B2(n_378), .C(n_387), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_399), .A2(n_394), .B1(n_392), .B2(n_370), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g425 ( .A1(n_374), .A2(n_398), .B(n_403), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_412), .A2(n_405), .B1(n_384), .B2(n_383), .C(n_380), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_414), .B(n_412), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g428 ( .A1(n_417), .A2(n_401), .B1(n_406), .B2(n_386), .Y(n_428) );
AO22x2_ASAP7_75t_L g429 ( .A1(n_419), .A2(n_398), .B1(n_395), .B2(n_381), .Y(n_429) );
AOI211xp5_ASAP7_75t_L g430 ( .A1(n_416), .A2(n_421), .B(n_425), .C(n_422), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_413), .B(n_365), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_431), .Y(n_432) );
OAI221xp5_ASAP7_75t_R g433 ( .A1(n_427), .A2(n_420), .B1(n_424), .B2(n_415), .C(n_404), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_429), .Y(n_434) );
NAND3xp33_ASAP7_75t_SL g435 ( .A(n_426), .B(n_418), .C(n_395), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_428), .A2(n_423), .B1(n_372), .B2(n_402), .Y(n_436) );
INVx3_ASAP7_75t_SL g437 ( .A(n_433), .Y(n_437) );
INVx4_ASAP7_75t_L g438 ( .A(n_434), .Y(n_438) );
INVx4_ASAP7_75t_L g439 ( .A(n_438), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_439), .A2(n_437), .B1(n_436), .B2(n_430), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_440), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_441), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_442), .A2(n_439), .B1(n_435), .B2(n_432), .Y(n_443) );
endmodule