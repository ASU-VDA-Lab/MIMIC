module fake_jpeg_21052_n_165 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_3),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx6p67_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_16),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_19),
.B1(n_11),
.B2(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_23),
.A2(n_20),
.B1(n_11),
.B2(n_19),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_40),
.B(n_43),
.C(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_13),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_24),
.A2(n_11),
.B1(n_12),
.B2(n_20),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_22),
.B1(n_17),
.B2(n_18),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_54),
.B1(n_56),
.B2(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_18),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_32),
.B(n_9),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_28),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_37),
.C(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_56),
.B1(n_47),
.B2(n_41),
.Y(n_80)
);

NOR2xp67_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_9),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_72),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_30),
.C(n_26),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_82),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_45),
.B(n_51),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_64),
.B(n_72),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_84),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_53),
.B1(n_55),
.B2(n_66),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_91),
.B(n_15),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_15),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_76),
.B(n_89),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_67),
.B1(n_61),
.B2(n_41),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_87),
.Y(n_115)
);

AOI322xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_67),
.A3(n_63),
.B1(n_15),
.B2(n_28),
.C1(n_25),
.C2(n_26),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_82),
.C(n_81),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_66),
.C(n_50),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_102),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_88),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_25),
.B1(n_29),
.B2(n_73),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_30),
.C(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_83),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_13),
.B(n_21),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_105),
.A2(n_81),
.B1(n_88),
.B2(n_83),
.Y(n_112)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_74),
.B(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_109),
.B(n_113),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_117),
.B1(n_106),
.B2(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_103),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_94),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_100),
.B1(n_101),
.B2(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_127),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_98),
.C(n_102),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_108),
.C(n_114),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_117),
.A2(n_94),
.B1(n_106),
.B2(n_21),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_115),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_136),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_135),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_137),
.C(n_124),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_21),
.C(n_16),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_126),
.B(n_8),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_21),
.C(n_16),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_120),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_142),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_123),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_144),
.A2(n_130),
.B1(n_138),
.B2(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_145),
.A2(n_127),
.B1(n_129),
.B2(n_3),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_150),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_1),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_2),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_8),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_140),
.B1(n_3),
.B2(n_4),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

AOI21x1_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_2),
.B(n_4),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_148),
.B(n_7),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_156),
.B(n_5),
.Y(n_159)
);

OAI21x1_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_159),
.B(n_153),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_157),
.B(n_155),
.C(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_7),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_7),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_164),
.Y(n_165)
);


endmodule