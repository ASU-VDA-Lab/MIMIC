module fake_netlist_1_8788_n_1187 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1187);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1187;
wire n_1173;
wire n_663;
wire n_791;
wire n_707;
wire n_513;
wire n_361;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_1122;
wire n_779;
wire n_993;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_1177;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_1185;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_1179;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1174;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1125;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_1183;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1025;
wire n_1011;
wire n_1132;
wire n_880;
wire n_1101;
wire n_1159;
wire n_630;
wire n_1155;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_1160;
wire n_1184;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_1046;
wire n_460;
wire n_950;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_1186;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_1157;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1017;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_1178;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_1181;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_1066;
wire n_1055;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1146;
wire n_287;
wire n_1108;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
INVx1_ASAP7_75t_L g252 ( .A(n_96), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_43), .Y(n_253) );
INVx1_ASAP7_75t_SL g254 ( .A(n_220), .Y(n_254) );
INVxp33_ASAP7_75t_L g255 ( .A(n_92), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_229), .Y(n_256) );
CKINVDCx14_ASAP7_75t_R g257 ( .A(n_130), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_59), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_157), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_156), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_240), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_138), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_166), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g265 ( .A(n_49), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_116), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_49), .Y(n_267) );
CKINVDCx16_ASAP7_75t_R g268 ( .A(n_34), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_63), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_210), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_31), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_172), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_86), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_62), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_63), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_246), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_50), .Y(n_277) );
INVxp33_ASAP7_75t_SL g278 ( .A(n_30), .Y(n_278) );
CKINVDCx16_ASAP7_75t_R g279 ( .A(n_44), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_5), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_12), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_109), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_26), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_38), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_215), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_40), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_191), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_53), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_189), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_33), .Y(n_290) );
INVxp33_ASAP7_75t_L g291 ( .A(n_120), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_52), .Y(n_292) );
INVxp67_ASAP7_75t_SL g293 ( .A(n_134), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_173), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_201), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_131), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_107), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_115), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_221), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_21), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_159), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_177), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_205), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_11), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_82), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_234), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_198), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_233), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_117), .Y(n_309) );
INVxp67_ASAP7_75t_SL g310 ( .A(n_181), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_0), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_30), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_202), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_182), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_66), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_200), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_110), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_75), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_6), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_5), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_238), .Y(n_321) );
INVxp67_ASAP7_75t_L g322 ( .A(n_10), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_87), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_148), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_28), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_37), .Y(n_326) );
CKINVDCx14_ASAP7_75t_R g327 ( .A(n_62), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_46), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_196), .Y(n_329) );
CKINVDCx16_ASAP7_75t_R g330 ( .A(n_136), .Y(n_330) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_174), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_250), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_126), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_61), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_139), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_175), .Y(n_336) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_84), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_245), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_18), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_183), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_26), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_52), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_55), .Y(n_343) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_216), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_46), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_152), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_118), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_147), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_127), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_197), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_145), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_14), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_211), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_164), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_53), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_119), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_25), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_129), .Y(n_358) );
INVxp33_ASAP7_75t_SL g359 ( .A(n_135), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_40), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_178), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_128), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_16), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g364 ( .A(n_237), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_207), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_11), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_165), .Y(n_367) );
INVxp33_ASAP7_75t_SL g368 ( .A(n_243), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_101), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_158), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_142), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_228), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_21), .Y(n_373) );
INVx2_ASAP7_75t_SL g374 ( .A(n_102), .Y(n_374) );
INVxp33_ASAP7_75t_SL g375 ( .A(n_59), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_32), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_149), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_83), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_125), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_122), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_111), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_95), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_140), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_137), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_179), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_327), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_304), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_329), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_329), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_329), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_329), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_271), .B(n_0), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_255), .B(n_1), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_275), .B(n_253), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_304), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_271), .B(n_1), .Y(n_397) );
NAND2xp33_ASAP7_75t_L g398 ( .A(n_255), .B(n_74), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_374), .B(n_2), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_347), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_374), .B(n_2), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_360), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_360), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_347), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_327), .Y(n_405) );
AND2x6_ASAP7_75t_L g406 ( .A(n_296), .B(n_76), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_347), .Y(n_407) );
OAI22xp5_ASAP7_75t_SL g408 ( .A1(n_277), .A2(n_3), .B1(n_4), .B2(n_6), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_265), .A2(n_3), .B1(n_4), .B2(n_7), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_366), .Y(n_410) );
BUFx2_ASAP7_75t_SL g411 ( .A(n_273), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_296), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_366), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_339), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_270), .B(n_7), .Y(n_415) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_298), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_263), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_330), .Y(n_418) );
AND2x6_ASAP7_75t_L g419 ( .A(n_397), .B(n_298), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_397), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_397), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_397), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_386), .B(n_291), .Y(n_423) );
AND2x6_ASAP7_75t_L g424 ( .A(n_394), .B(n_393), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_395), .B(n_268), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_417), .B(n_263), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_412), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_386), .B(n_291), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_417), .Y(n_430) );
AND2x6_ASAP7_75t_L g431 ( .A(n_393), .B(n_318), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_388), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_387), .B(n_337), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_417), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_387), .B(n_294), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_396), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_388), .Y(n_437) );
NAND2xp33_ASAP7_75t_SL g438 ( .A(n_405), .B(n_273), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_396), .B(n_344), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_411), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_411), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_402), .Y(n_442) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_388), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_402), .B(n_317), .Y(n_444) );
AND2x6_ASAP7_75t_L g445 ( .A(n_399), .B(n_318), .Y(n_445) );
INVx4_ASAP7_75t_L g446 ( .A(n_406), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_403), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_410), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_412), .B(n_252), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_410), .B(n_323), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_413), .Y(n_452) );
INVxp33_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_413), .B(n_364), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_418), .B(n_324), .Y(n_455) );
NAND2xp33_ASAP7_75t_R g456 ( .A(n_414), .B(n_278), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_398), .B(n_322), .C(n_274), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_401), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_412), .B(n_256), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_412), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_414), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_414), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_408), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_412), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_452), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_420), .A2(n_406), .B1(n_375), .B2(n_278), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_453), .B(n_359), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_441), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_453), .B(n_359), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_425), .B(n_279), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_452), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g473 ( .A(n_440), .B(n_258), .Y(n_473) );
INVx5_ASAP7_75t_L g474 ( .A(n_419), .Y(n_474) );
BUFx4f_ASAP7_75t_L g475 ( .A(n_424), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_427), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_429), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_446), .B(n_259), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_446), .B(n_260), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_442), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_447), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_448), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_435), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_433), .B(n_264), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_421), .B(n_262), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_424), .A2(n_406), .B1(n_375), .B2(n_269), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_458), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_439), .B(n_295), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_424), .A2(n_406), .B1(n_281), .B2(n_283), .Y(n_490) );
INVx2_ASAP7_75t_SL g491 ( .A(n_435), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_454), .Y(n_492) );
AND2x6_ASAP7_75t_L g493 ( .A(n_422), .B(n_272), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_428), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_449), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_459), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_419), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_424), .B(n_295), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_458), .Y(n_499) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_455), .B(n_409), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_424), .B(n_336), .Y(n_501) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_427), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_422), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_430), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_434), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_457), .B(n_276), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_444), .B(n_336), .Y(n_507) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_419), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_419), .Y(n_509) );
OR2x6_ASAP7_75t_L g510 ( .A(n_444), .B(n_408), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_451), .B(n_282), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_426), .A2(n_308), .B1(n_309), .B2(n_289), .Y(n_512) );
INVx4_ASAP7_75t_L g513 ( .A(n_419), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_445), .B(n_368), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_438), .Y(n_515) );
NAND3xp33_ASAP7_75t_SL g516 ( .A(n_464), .B(n_325), .C(n_274), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_431), .Y(n_517) );
AO22x1_ASAP7_75t_L g518 ( .A1(n_431), .A2(n_368), .B1(n_326), .B2(n_334), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_450), .B(n_285), .Y(n_519) );
BUFx3_ASAP7_75t_L g520 ( .A(n_445), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_431), .B(n_308), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_431), .B(n_362), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_465), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_461), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_445), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_450), .B(n_369), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_460), .B(n_257), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_460), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_456), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_461), .B(n_257), .Y(n_530) );
AND3x2_ASAP7_75t_SL g531 ( .A(n_456), .B(n_280), .C(n_277), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_462), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_465), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_463), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_443), .A2(n_321), .B1(n_340), .B2(n_309), .Y(n_535) );
BUFx4f_ASAP7_75t_L g536 ( .A(n_443), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_432), .B(n_261), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_432), .A2(n_406), .B1(n_284), .B2(n_286), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_432), .B(n_314), .Y(n_539) );
NOR2x1p5_ASAP7_75t_L g540 ( .A(n_432), .B(n_325), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_437), .B(n_351), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_437), .Y(n_542) );
AND2x6_ASAP7_75t_L g543 ( .A(n_437), .B(n_287), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_443), .B(n_365), .Y(n_544) );
BUFx4f_ASAP7_75t_L g545 ( .A(n_424), .Y(n_545) );
INVx5_ASAP7_75t_L g546 ( .A(n_419), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_423), .B(n_335), .Y(n_547) );
NOR2xp33_ASAP7_75t_SL g548 ( .A(n_513), .B(n_321), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_494), .Y(n_549) );
INVxp67_ASAP7_75t_SL g550 ( .A(n_535), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_478), .B(n_512), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_503), .Y(n_552) );
INVx3_ASAP7_75t_L g553 ( .A(n_513), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_491), .Y(n_554) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_508), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_473), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_503), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_486), .A2(n_310), .B(n_293), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_487), .A2(n_371), .B1(n_340), .B2(n_280), .Y(n_559) );
BUFx2_ASAP7_75t_L g560 ( .A(n_484), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_486), .A2(n_331), .B(n_299), .Y(n_561) );
AOI21xp33_ASAP7_75t_L g562 ( .A1(n_514), .A2(n_301), .B(n_297), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_477), .A2(n_288), .B(n_290), .C(n_267), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_492), .B(n_326), .Y(n_564) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_508), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_481), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_482), .A2(n_311), .B(n_312), .C(n_292), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_469), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_483), .A2(n_319), .B(n_320), .C(n_315), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_495), .B(n_334), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_468), .B(n_342), .Y(n_571) );
O2A1O1Ixp5_ASAP7_75t_L g572 ( .A1(n_511), .A2(n_303), .B(n_305), .C(n_302), .Y(n_572) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_514), .A2(n_341), .B(n_343), .C(n_328), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_468), .B(n_342), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_471), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_472), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_466), .Y(n_577) );
BUFx3_ASAP7_75t_L g578 ( .A(n_521), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_487), .A2(n_300), .B1(n_363), .B2(n_357), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_479), .A2(n_307), .B(n_306), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_504), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_496), .B(n_376), .Y(n_582) );
NAND2x1p5_ASAP7_75t_L g583 ( .A(n_474), .B(n_339), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_510), .B(n_345), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g585 ( .A1(n_511), .A2(n_372), .B(n_384), .C(n_300), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_521), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_505), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_532), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_534), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_479), .A2(n_316), .B(n_313), .Y(n_590) );
INVx2_ASAP7_75t_SL g591 ( .A(n_540), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_518), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_529), .A2(n_406), .B1(n_352), .B2(n_373), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_515), .Y(n_594) );
INVx4_ASAP7_75t_L g595 ( .A(n_508), .Y(n_595) );
INVx2_ASAP7_75t_SL g596 ( .A(n_475), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_528), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_485), .Y(n_598) );
INVx5_ASAP7_75t_L g599 ( .A(n_508), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_475), .A2(n_355), .B1(n_373), .B2(n_352), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_545), .A2(n_333), .B1(n_338), .B2(n_332), .Y(n_601) );
INVx5_ASAP7_75t_L g602 ( .A(n_474), .Y(n_602) );
BUFx2_ASAP7_75t_L g603 ( .A(n_493), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_489), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_470), .B(n_339), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_474), .B(n_346), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_470), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_510), .A2(n_406), .B1(n_339), .B2(n_416), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_502), .Y(n_609) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_509), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_493), .B(n_348), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_493), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_547), .B(n_254), .Y(n_613) );
OAI22xp5_ASAP7_75t_SL g614 ( .A1(n_510), .A2(n_353), .B1(n_354), .B2(n_350), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_474), .B(n_356), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_493), .B(n_358), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_500), .A2(n_367), .B1(n_370), .B2(n_361), .Y(n_617) );
BUFx12f_ASAP7_75t_L g618 ( .A(n_493), .Y(n_618) );
BUFx12f_ASAP7_75t_L g619 ( .A(n_543), .Y(n_619) );
INVx4_ASAP7_75t_L g620 ( .A(n_546), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_502), .Y(n_621) );
INVx4_ASAP7_75t_L g622 ( .A(n_546), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_502), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_507), .B(n_377), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_516), .Y(n_625) );
INVx3_ASAP7_75t_SL g626 ( .A(n_506), .Y(n_626) );
BUFx2_ASAP7_75t_L g627 ( .A(n_509), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_498), .Y(n_628) );
BUFx12f_ASAP7_75t_L g629 ( .A(n_543), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_545), .B(n_8), .Y(n_630) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_546), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_501), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_480), .A2(n_379), .B(n_378), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_497), .Y(n_634) );
INVx4_ASAP7_75t_L g635 ( .A(n_546), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_520), .Y(n_636) );
INVx2_ASAP7_75t_SL g637 ( .A(n_517), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_526), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_516), .A2(n_416), .B1(n_381), .B2(n_382), .Y(n_639) );
AOI21x1_ASAP7_75t_L g640 ( .A1(n_480), .A2(n_383), .B(n_380), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_502), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_522), .Y(n_642) );
OR2x6_ASAP7_75t_L g643 ( .A(n_531), .B(n_385), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_467), .A2(n_266), .B1(n_349), .B2(n_414), .C(n_416), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_543), .Y(n_645) );
BUFx12f_ASAP7_75t_L g646 ( .A(n_543), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_467), .B(n_416), .Y(n_647) );
BUFx12f_ASAP7_75t_L g648 ( .A(n_543), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_519), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_531), .B(n_8), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_490), .B(n_416), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_490), .B(n_9), .Y(n_652) );
AOI21xp33_ASAP7_75t_L g653 ( .A1(n_525), .A2(n_416), .B(n_392), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_519), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_520), .Y(n_655) );
INVx4_ASAP7_75t_L g656 ( .A(n_536), .Y(n_656) );
INVx4_ASAP7_75t_L g657 ( .A(n_536), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_527), .Y(n_658) );
NAND2x1p5_ASAP7_75t_L g659 ( .A(n_476), .B(n_390), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_530), .Y(n_660) );
CKINVDCx16_ASAP7_75t_R g661 ( .A(n_537), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_539), .Y(n_662) );
INVx3_ASAP7_75t_L g663 ( .A(n_533), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_541), .B(n_388), .Y(n_664) );
BUFx2_ASAP7_75t_L g665 ( .A(n_544), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_488), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_524), .A2(n_392), .B(n_390), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_538), .A2(n_407), .B1(n_404), .B2(n_400), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_533), .B(n_9), .Y(n_669) );
BUFx2_ASAP7_75t_L g670 ( .A(n_488), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_499), .B(n_400), .Y(n_671) );
INVx3_ASAP7_75t_L g672 ( .A(n_499), .Y(n_672) );
AO21x2_ASAP7_75t_L g673 ( .A1(n_651), .A2(n_407), .B(n_404), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_566), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_551), .B(n_10), .Y(n_675) );
AOI22x1_ASAP7_75t_L g676 ( .A1(n_658), .A2(n_523), .B1(n_542), .B2(n_391), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_587), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_581), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_588), .Y(n_679) );
OR2x2_ASAP7_75t_L g680 ( .A(n_564), .B(n_12), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_589), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_605), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_564), .B(n_13), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_647), .A2(n_389), .B(n_388), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_559), .B(n_15), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_568), .Y(n_686) );
NAND2x1p5_ASAP7_75t_L g687 ( .A(n_656), .B(n_389), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_666), .Y(n_688) );
OAI21x1_ASAP7_75t_L g689 ( .A1(n_583), .A2(n_391), .B(n_389), .Y(n_689) );
OR2x6_ASAP7_75t_L g690 ( .A(n_618), .B(n_16), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_559), .B(n_17), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_670), .Y(n_692) );
INVx4_ASAP7_75t_SL g693 ( .A(n_619), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_L g694 ( .A1(n_573), .A2(n_17), .B(n_18), .C(n_19), .Y(n_694) );
BUFx2_ASAP7_75t_L g695 ( .A(n_556), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_597), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_548), .B(n_389), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_577), .Y(n_698) );
OAI22xp5_ASAP7_75t_SL g699 ( .A1(n_643), .A2(n_19), .B1(n_20), .B2(n_22), .Y(n_699) );
OAI21x1_ASAP7_75t_L g700 ( .A1(n_583), .A2(n_391), .B(n_78), .Y(n_700) );
INVx3_ASAP7_75t_L g701 ( .A(n_656), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_560), .Y(n_702) );
OAI21x1_ASAP7_75t_L g703 ( .A1(n_640), .A2(n_391), .B(n_79), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_672), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_548), .B(n_20), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_598), .B(n_23), .Y(n_706) );
NAND2x1p5_ASAP7_75t_L g707 ( .A(n_657), .B(n_24), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_604), .B(n_27), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_579), .A2(n_28), .B1(n_29), .B2(n_31), .Y(n_709) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_554), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_575), .B(n_29), .Y(n_711) );
OAI21x1_ASAP7_75t_L g712 ( .A1(n_659), .A2(n_80), .B(n_77), .Y(n_712) );
INVx5_ASAP7_75t_L g713 ( .A(n_629), .Y(n_713) );
OAI21x1_ASAP7_75t_L g714 ( .A1(n_659), .A2(n_85), .B(n_81), .Y(n_714) );
NAND2x1_ASAP7_75t_L g715 ( .A(n_657), .B(n_88), .Y(n_715) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_655), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_579), .A2(n_32), .B1(n_33), .B2(n_34), .Y(n_717) );
AND2x4_ASAP7_75t_L g718 ( .A(n_549), .B(n_35), .Y(n_718) );
BUFx2_ASAP7_75t_L g719 ( .A(n_643), .Y(n_719) );
OAI21x1_ASAP7_75t_L g720 ( .A1(n_664), .A2(n_90), .B(n_89), .Y(n_720) );
OA21x2_ASAP7_75t_L g721 ( .A1(n_653), .A2(n_93), .B(n_91), .Y(n_721) );
AOI21x1_ASAP7_75t_L g722 ( .A1(n_611), .A2(n_97), .B(n_94), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_582), .Y(n_723) );
OA21x2_ASAP7_75t_L g724 ( .A1(n_667), .A2(n_99), .B(n_98), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_582), .Y(n_725) );
BUFx2_ASAP7_75t_L g726 ( .A(n_578), .Y(n_726) );
OA21x2_ASAP7_75t_L g727 ( .A1(n_667), .A2(n_103), .B(n_100), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_570), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_650), .A2(n_35), .B1(n_36), .B2(n_37), .Y(n_729) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_625), .A2(n_36), .B1(n_38), .B2(n_39), .Y(n_730) );
NAND2x1_ASAP7_75t_L g731 ( .A(n_620), .B(n_104), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_624), .A2(n_590), .B(n_580), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_638), .B(n_39), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_570), .Y(n_734) );
INVxp67_ASAP7_75t_L g735 ( .A(n_600), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_576), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_607), .B(n_41), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_550), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_628), .B(n_42), .Y(n_739) );
OAI21x1_ASAP7_75t_L g740 ( .A1(n_609), .A2(n_162), .B(n_249), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_562), .A2(n_44), .B(n_45), .Y(n_741) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_555), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_586), .B(n_45), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_624), .A2(n_163), .B(n_248), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_649), .Y(n_745) );
AND2x4_ASAP7_75t_L g746 ( .A(n_603), .B(n_47), .Y(n_746) );
OAI21x1_ASAP7_75t_L g747 ( .A1(n_621), .A2(n_161), .B(n_247), .Y(n_747) );
AO31x2_ASAP7_75t_L g748 ( .A1(n_601), .A2(n_47), .A3(n_48), .B(n_50), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_623), .A2(n_167), .B(n_244), .Y(n_749) );
OAI21x1_ASAP7_75t_L g750 ( .A1(n_641), .A2(n_160), .B(n_241), .Y(n_750) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_555), .Y(n_751) );
BUFx3_ASAP7_75t_L g752 ( .A(n_646), .Y(n_752) );
AOI22xp33_ASAP7_75t_SL g753 ( .A1(n_614), .A2(n_48), .B1(n_51), .B2(n_54), .Y(n_753) );
OAI21x1_ASAP7_75t_L g754 ( .A1(n_671), .A2(n_155), .B(n_239), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_669), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_584), .B(n_51), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_632), .B(n_54), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_654), .Y(n_758) );
AND2x4_ASAP7_75t_L g759 ( .A(n_612), .B(n_56), .Y(n_759) );
OAI21x1_ASAP7_75t_L g760 ( .A1(n_671), .A2(n_169), .B(n_236), .Y(n_760) );
OAI21xp5_ASAP7_75t_L g761 ( .A1(n_562), .A2(n_57), .B(n_58), .Y(n_761) );
OAI21x1_ASAP7_75t_L g762 ( .A1(n_616), .A2(n_168), .B(n_235), .Y(n_762) );
INVx3_ASAP7_75t_L g763 ( .A(n_620), .Y(n_763) );
AO21x2_ASAP7_75t_L g764 ( .A1(n_580), .A2(n_154), .B(n_232), .Y(n_764) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_555), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_662), .Y(n_766) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_565), .Y(n_767) );
OAI21x1_ASAP7_75t_L g768 ( .A1(n_590), .A2(n_153), .B(n_231), .Y(n_768) );
OA21x2_ASAP7_75t_L g769 ( .A1(n_608), .A2(n_151), .B(n_230), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g770 ( .A1(n_563), .A2(n_569), .B1(n_567), .B2(n_585), .C(n_571), .Y(n_770) );
BUFx2_ASAP7_75t_L g771 ( .A(n_648), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_596), .B(n_60), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_633), .A2(n_170), .B(n_227), .Y(n_773) );
NAND2x1_ASAP7_75t_L g774 ( .A(n_622), .B(n_105), .Y(n_774) );
AND2x4_ASAP7_75t_L g775 ( .A(n_592), .B(n_61), .Y(n_775) );
NAND2x1p5_ASAP7_75t_L g776 ( .A(n_599), .B(n_64), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_552), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_642), .B(n_65), .Y(n_778) );
OAI21x1_ASAP7_75t_L g779 ( .A1(n_553), .A2(n_171), .B(n_226), .Y(n_779) );
INVx3_ASAP7_75t_L g780 ( .A(n_622), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_571), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_781) );
NAND2x1p5_ASAP7_75t_L g782 ( .A(n_599), .B(n_67), .Y(n_782) );
INVx3_ASAP7_75t_SL g783 ( .A(n_594), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_574), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_561), .A2(n_176), .B(n_225), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_557), .Y(n_786) );
OAI21xp5_ASAP7_75t_L g787 ( .A1(n_561), .A2(n_68), .B(n_69), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_574), .A2(n_180), .B(n_224), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_613), .B(n_70), .Y(n_789) );
AOI221xp5_ASAP7_75t_L g790 ( .A1(n_601), .A2(n_70), .B1(n_71), .B2(n_72), .C(n_73), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_652), .A2(n_71), .B1(n_72), .B2(n_73), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_665), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_617), .B(n_106), .Y(n_793) );
AOI221xp5_ASAP7_75t_SL g794 ( .A1(n_644), .A2(n_108), .B1(n_112), .B2(n_113), .C(n_114), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_663), .Y(n_795) );
BUFx3_ASAP7_75t_L g796 ( .A(n_591), .Y(n_796) );
INVx8_ASAP7_75t_L g797 ( .A(n_602), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_630), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_661), .B(n_121), .Y(n_799) );
NAND3xp33_ASAP7_75t_SL g800 ( .A(n_639), .B(n_123), .C(n_124), .Y(n_800) );
NAND2x1p5_ASAP7_75t_L g801 ( .A(n_599), .B(n_251), .Y(n_801) );
OA21x2_ASAP7_75t_L g802 ( .A1(n_572), .A2(n_132), .B(n_133), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_698), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_784), .B(n_626), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_692), .B(n_634), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_685), .A2(n_660), .B1(n_606), .B2(n_615), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_691), .A2(n_606), .B1(n_615), .B2(n_558), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_792), .B(n_734), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_674), .Y(n_809) );
AOI21xp33_ASAP7_75t_SL g810 ( .A1(n_783), .A2(n_668), .B(n_593), .Y(n_810) );
INVx3_ASAP7_75t_L g811 ( .A(n_797), .Y(n_811) );
OAI22xp33_ASAP7_75t_L g812 ( .A1(n_709), .A2(n_645), .B1(n_627), .B2(n_599), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_770), .B(n_558), .Y(n_813) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_797), .Y(n_814) );
AOI21x1_ASAP7_75t_L g815 ( .A1(n_684), .A2(n_668), .B(n_637), .Y(n_815) );
NAND2xp5_ASAP7_75t_SL g816 ( .A(n_794), .B(n_565), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_677), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_735), .A2(n_610), .B1(n_595), .B2(n_636), .Y(n_818) );
INVx4_ASAP7_75t_SL g819 ( .A(n_690), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_738), .A2(n_610), .B1(n_636), .B2(n_553), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_678), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_732), .A2(n_565), .B(n_636), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g823 ( .A1(n_711), .A2(n_737), .B1(n_725), .B2(n_723), .C(n_791), .Y(n_823) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_746), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_679), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g826 ( .A1(n_719), .A2(n_602), .B1(n_635), .B2(n_610), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_681), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_695), .B(n_602), .Y(n_828) );
AOI221xp5_ASAP7_75t_L g829 ( .A1(n_791), .A2(n_635), .B1(n_631), .B2(n_602), .C(n_144), .Y(n_829) );
OAI22xp33_ASAP7_75t_L g830 ( .A1(n_709), .A2(n_631), .B1(n_141), .B2(n_143), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_710), .B(n_702), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_699), .A2(n_631), .B1(n_146), .B2(n_150), .Y(n_832) );
INVx1_ASAP7_75t_SL g833 ( .A(n_686), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_699), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_834) );
OA21x2_ASAP7_75t_L g835 ( .A1(n_684), .A2(n_223), .B(n_187), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_688), .Y(n_836) );
OA21x2_ASAP7_75t_L g837 ( .A1(n_794), .A2(n_222), .B(n_188), .Y(n_837) );
INVxp67_ASAP7_75t_SL g838 ( .A(n_759), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_706), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_696), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_790), .A2(n_190), .B1(n_192), .B2(n_193), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_790), .A2(n_194), .B1(n_195), .B2(n_199), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_706), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g844 ( .A(n_752), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_690), .B(n_203), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_690), .B(n_204), .Y(n_846) );
OAI221xp5_ASAP7_75t_L g847 ( .A1(n_798), .A2(n_206), .B1(n_208), .B2(n_209), .C(n_212), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_730), .A2(n_761), .B1(n_741), .B2(n_789), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_730), .A2(n_213), .B1(n_214), .B2(n_217), .Y(n_849) );
OAI21x1_ASAP7_75t_L g850 ( .A1(n_689), .A2(n_218), .B(n_219), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_756), .B(n_708), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_736), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_741), .A2(n_761), .B1(n_675), .B2(n_717), .Y(n_853) );
AND2x4_ASAP7_75t_L g854 ( .A(n_693), .B(n_713), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_682), .A2(n_708), .B1(n_680), .B2(n_683), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_718), .A2(n_733), .B1(n_787), .B2(n_729), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_743), .B(n_733), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_755), .A2(n_778), .B1(n_739), .B2(n_757), .Y(n_858) );
BUFx2_ASAP7_75t_L g859 ( .A(n_716), .Y(n_859) );
AOI222xp33_ASAP7_75t_L g860 ( .A1(n_775), .A2(n_787), .B1(n_772), .B2(n_705), .C1(n_726), .C2(n_693), .Y(n_860) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_776), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_707), .Y(n_862) );
AOI222xp33_ASAP7_75t_L g863 ( .A1(n_775), .A2(n_693), .B1(n_781), .B2(n_778), .C1(n_757), .C2(n_739), .Y(n_863) );
AOI22xp33_ASAP7_75t_SL g864 ( .A1(n_782), .A2(n_713), .B1(n_799), .B2(n_797), .Y(n_864) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_742), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_745), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_758), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_753), .A2(n_729), .B1(n_793), .B2(n_771), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_748), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_800), .A2(n_697), .B1(n_701), .B2(n_786), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_713), .B(n_777), .Y(n_871) );
INVx2_ASAP7_75t_SL g872 ( .A(n_796), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_748), .B(n_701), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_673), .Y(n_874) );
AND2x4_ASAP7_75t_L g875 ( .A(n_763), .B(n_780), .Y(n_875) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_801), .A2(n_800), .B1(n_744), .B2(n_769), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_673), .Y(n_877) );
OA21x2_ASAP7_75t_L g878 ( .A1(n_754), .A2(n_760), .B(n_762), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_795), .B(n_704), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_748), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_687), .A2(n_676), .B1(n_769), .B2(n_744), .Y(n_881) );
OA21x2_ASAP7_75t_L g882 ( .A1(n_703), .A2(n_750), .B(n_747), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_687), .B(n_764), .Y(n_883) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_742), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_779), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_768), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_788), .B(n_785), .Y(n_887) );
OA21x2_ASAP7_75t_L g888 ( .A1(n_740), .A2(n_749), .B(n_773), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_764), .A2(n_802), .B1(n_715), .B2(n_721), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_742), .B(n_767), .Y(n_890) );
AO21x2_ASAP7_75t_L g891 ( .A1(n_722), .A2(n_700), .B(n_720), .Y(n_891) );
A2O1A1Ixp33_ASAP7_75t_L g892 ( .A1(n_731), .A2(n_774), .B(n_714), .C(n_712), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_724), .Y(n_893) );
INVxp33_ASAP7_75t_L g894 ( .A(n_751), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_727), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_767), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_751), .B(n_765), .Y(n_897) );
INVx2_ASAP7_75t_SL g898 ( .A(n_765), .Y(n_898) );
AOI211xp5_ASAP7_75t_L g899 ( .A1(n_765), .A2(n_614), .B(n_730), .C(n_699), .Y(n_899) );
A2O1A1Ixp33_ASAP7_75t_L g900 ( .A1(n_694), .A2(n_732), .B(n_709), .C(n_741), .Y(n_900) );
AND2x4_ASAP7_75t_L g901 ( .A(n_693), .B(n_728), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_766), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_766), .Y(n_903) );
OAI22xp33_ASAP7_75t_L g904 ( .A1(n_709), .A2(n_548), .B1(n_691), .B2(n_685), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_784), .B(n_728), .Y(n_905) );
AOI222xp33_ASAP7_75t_L g906 ( .A1(n_699), .A2(n_408), .B1(n_464), .B2(n_614), .C1(n_730), .C2(n_728), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_698), .Y(n_907) );
BUFx6f_ASAP7_75t_L g908 ( .A(n_797), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_735), .A2(n_535), .B1(n_559), .B2(n_551), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_766), .Y(n_910) );
AOI221xp5_ASAP7_75t_L g911 ( .A1(n_728), .A2(n_575), .B1(n_471), .B2(n_734), .C(n_607), .Y(n_911) );
BUFx3_ASAP7_75t_L g912 ( .A(n_814), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_906), .A2(n_904), .B1(n_848), .B2(n_856), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_869), .Y(n_914) );
BUFx8_ASAP7_75t_L g915 ( .A(n_814), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_880), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_838), .B(n_803), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_838), .B(n_907), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_873), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_836), .B(n_825), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_866), .Y(n_921) );
OAI221xp5_ASAP7_75t_L g922 ( .A1(n_911), .A2(n_899), .B1(n_868), .B2(n_848), .C(n_823), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_867), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_852), .B(n_839), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_843), .B(n_809), .Y(n_925) );
INVx2_ASAP7_75t_L g926 ( .A(n_874), .Y(n_926) );
INVx2_ASAP7_75t_SL g927 ( .A(n_814), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_840), .B(n_817), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_821), .B(n_827), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_905), .B(n_808), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_902), .Y(n_931) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_805), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_903), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_910), .Y(n_934) );
INVx3_ASAP7_75t_SL g935 ( .A(n_814), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_856), .B(n_824), .Y(n_936) );
AND2x4_ASAP7_75t_L g937 ( .A(n_890), .B(n_897), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_861), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_877), .Y(n_939) );
INVx2_ASAP7_75t_L g940 ( .A(n_893), .Y(n_940) );
OR2x2_ASAP7_75t_L g941 ( .A(n_824), .B(n_909), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_851), .B(n_855), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_861), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_885), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_858), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_855), .B(n_813), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_886), .Y(n_947) );
INVx3_ASAP7_75t_L g948 ( .A(n_908), .Y(n_948) );
INVx2_ASAP7_75t_L g949 ( .A(n_895), .Y(n_949) );
BUFx3_ASAP7_75t_L g950 ( .A(n_908), .Y(n_950) );
BUFx2_ASAP7_75t_L g951 ( .A(n_865), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_857), .B(n_875), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_815), .Y(n_953) );
OR2x2_ASAP7_75t_L g954 ( .A(n_904), .B(n_831), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_883), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_884), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_884), .Y(n_957) );
OR2x2_ASAP7_75t_L g958 ( .A(n_862), .B(n_859), .Y(n_958) );
OR2x2_ASAP7_75t_L g959 ( .A(n_806), .B(n_804), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_860), .A2(n_863), .B1(n_819), .B2(n_812), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_875), .B(n_806), .Y(n_961) );
INVx1_ASAP7_75t_SL g962 ( .A(n_833), .Y(n_962) );
INVx1_ASAP7_75t_SL g963 ( .A(n_844), .Y(n_963) );
INVx2_ASAP7_75t_SL g964 ( .A(n_854), .Y(n_964) );
INVx3_ASAP7_75t_L g965 ( .A(n_811), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_879), .B(n_819), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_900), .Y(n_967) );
OAI31xp33_ASAP7_75t_L g968 ( .A1(n_812), .A2(n_830), .A3(n_845), .B(n_846), .Y(n_968) );
INVx3_ASAP7_75t_L g969 ( .A(n_811), .Y(n_969) );
INVx3_ASAP7_75t_L g970 ( .A(n_896), .Y(n_970) );
BUFx2_ASAP7_75t_L g971 ( .A(n_865), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_879), .B(n_819), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_900), .B(n_849), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_849), .B(n_901), .Y(n_974) );
INVxp67_ASAP7_75t_SL g975 ( .A(n_830), .Y(n_975) );
AND2x4_ASAP7_75t_L g976 ( .A(n_898), .B(n_822), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_816), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_901), .B(n_853), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_864), .A2(n_853), .B1(n_807), .B2(n_842), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_816), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_835), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_807), .B(n_834), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_834), .B(n_828), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_878), .Y(n_984) );
INVx2_ASAP7_75t_SL g985 ( .A(n_854), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_832), .B(n_894), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_832), .B(n_841), .Y(n_987) );
INVx4_ASAP7_75t_L g988 ( .A(n_871), .Y(n_988) );
OR2x2_ASAP7_75t_L g989 ( .A(n_872), .B(n_887), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_841), .B(n_842), .Y(n_990) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_829), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_878), .Y(n_992) );
INVx2_ASAP7_75t_SL g993 ( .A(n_850), .Y(n_993) );
NOR2xp33_ASAP7_75t_L g994 ( .A(n_810), .B(n_847), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_930), .B(n_820), .Y(n_995) );
BUFx2_ASAP7_75t_L g996 ( .A(n_951), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_942), .B(n_826), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_955), .B(n_837), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_913), .B(n_818), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_925), .B(n_870), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_919), .B(n_878), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_922), .A2(n_870), .B1(n_876), .B2(n_881), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_946), .B(n_889), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_929), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_946), .B(n_889), .Y(n_1005) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_915), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_936), .B(n_891), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_936), .B(n_891), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g1009 ( .A1(n_979), .A2(n_876), .B1(n_892), .B2(n_888), .C(n_882), .Y(n_1009) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_951), .Y(n_1010) );
NAND3xp33_ASAP7_75t_L g1011 ( .A(n_994), .B(n_888), .C(n_882), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_928), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_921), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_925), .B(n_932), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_924), .B(n_882), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_921), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_967), .B(n_917), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_923), .Y(n_1018) );
NAND2xp5_ASAP7_75t_SL g1019 ( .A(n_968), .B(n_960), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_924), .B(n_920), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_958), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_923), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_920), .B(n_952), .Y(n_1023) );
INVx2_ASAP7_75t_SL g1024 ( .A(n_915), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_940), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_917), .B(n_918), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_918), .B(n_945), .Y(n_1027) );
BUFx3_ASAP7_75t_L g1028 ( .A(n_915), .Y(n_1028) );
OR2x2_ASAP7_75t_L g1029 ( .A(n_954), .B(n_989), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_945), .B(n_978), .Y(n_1030) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_989), .B(n_941), .Y(n_1031) );
AOI221xp5_ASAP7_75t_L g1032 ( .A1(n_931), .A2(n_934), .B1(n_933), .B2(n_973), .C(n_952), .Y(n_1032) );
INVx2_ASAP7_75t_SL g1033 ( .A(n_915), .Y(n_1033) );
AND2x4_ASAP7_75t_L g1034 ( .A(n_914), .B(n_916), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_978), .B(n_914), .Y(n_1035) );
AND2x4_ASAP7_75t_L g1036 ( .A(n_916), .B(n_976), .Y(n_1036) );
BUFx3_ASAP7_75t_L g1037 ( .A(n_935), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_931), .Y(n_1038) );
AOI33xp33_ASAP7_75t_L g1039 ( .A1(n_934), .A2(n_962), .A3(n_963), .B1(n_938), .B2(n_943), .B3(n_973), .Y(n_1039) );
AND2x4_ASAP7_75t_L g1040 ( .A(n_976), .B(n_944), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_958), .Y(n_1041) );
OAI31xp33_ASAP7_75t_L g1042 ( .A1(n_959), .A2(n_982), .A3(n_974), .B(n_987), .Y(n_1042) );
AND2x4_ASAP7_75t_L g1043 ( .A(n_976), .B(n_944), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_988), .B(n_961), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_956), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_988), .B(n_961), .Y(n_1046) );
INVx2_ASAP7_75t_SL g1047 ( .A(n_912), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_956), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_937), .B(n_939), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_957), .Y(n_1050) );
OAI31xp33_ASAP7_75t_SL g1051 ( .A1(n_966), .A2(n_972), .A3(n_975), .B(n_983), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_947), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_1021), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1013), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1004), .B(n_937), .Y(n_1055) );
AND4x1_ASAP7_75t_L g1056 ( .A(n_1051), .B(n_972), .C(n_966), .D(n_987), .Y(n_1056) );
OR2x2_ASAP7_75t_L g1057 ( .A(n_1031), .B(n_926), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1030), .B(n_949), .Y(n_1058) );
NAND2xp5_ASAP7_75t_SL g1059 ( .A(n_1039), .B(n_971), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1016), .Y(n_1060) );
AND2x4_ASAP7_75t_SL g1061 ( .A(n_1024), .B(n_1033), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1025), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1003), .B(n_1005), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1052), .Y(n_1064) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_1029), .B(n_939), .Y(n_1065) );
INVx2_ASAP7_75t_L g1066 ( .A(n_1025), .Y(n_1066) );
INVxp67_ASAP7_75t_L g1067 ( .A(n_1006), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1018), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1034), .Y(n_1069) );
INVx5_ASAP7_75t_SL g1070 ( .A(n_1028), .Y(n_1070) );
HB1xp67_ASAP7_75t_L g1071 ( .A(n_996), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1022), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g1073 ( .A(n_1010), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1038), .Y(n_1074) );
OR2x2_ASAP7_75t_L g1075 ( .A(n_1029), .B(n_939), .Y(n_1075) );
INVx1_ASAP7_75t_SL g1076 ( .A(n_1037), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1003), .B(n_949), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_1035), .B(n_971), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1014), .Y(n_1079) );
OAI31xp33_ASAP7_75t_L g1080 ( .A1(n_1019), .A2(n_991), .A3(n_985), .B(n_964), .Y(n_1080) );
OR2x2_ASAP7_75t_L g1081 ( .A(n_1035), .B(n_1026), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1045), .Y(n_1082) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_1036), .B(n_976), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_1026), .B(n_992), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1048), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1005), .B(n_992), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1050), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1012), .B(n_937), .Y(n_1088) );
AND2x4_ASAP7_75t_L g1089 ( .A(n_1036), .B(n_980), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1007), .B(n_977), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1010), .B(n_984), .Y(n_1091) );
INVxp33_ASAP7_75t_SL g1092 ( .A(n_1037), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1007), .B(n_977), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1008), .B(n_984), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1020), .B(n_983), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1034), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1064), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1063), .B(n_1042), .Y(n_1098) );
INVx1_ASAP7_75t_SL g1099 ( .A(n_1061), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1086), .B(n_1001), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1094), .B(n_1001), .Y(n_1101) );
INVx2_ASAP7_75t_L g1102 ( .A(n_1062), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_1071), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1064), .Y(n_1104) );
AND2x4_ASAP7_75t_L g1105 ( .A(n_1083), .B(n_1036), .Y(n_1105) );
NOR2xp33_ASAP7_75t_L g1106 ( .A(n_1067), .B(n_1033), .Y(n_1106) );
AND2x4_ASAP7_75t_L g1107 ( .A(n_1083), .B(n_1040), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1094), .B(n_1049), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1054), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_1063), .B(n_1032), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_1081), .B(n_1015), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1060), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1081), .B(n_1027), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1068), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1072), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_1073), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1077), .B(n_1049), .Y(n_1117) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_1053), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1079), .B(n_1041), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1074), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1077), .B(n_1043), .Y(n_1121) );
INVxp67_ASAP7_75t_SL g1122 ( .A(n_1059), .Y(n_1122) );
NOR2xp67_ASAP7_75t_L g1123 ( .A(n_1084), .B(n_1011), .Y(n_1123) );
OAI31xp33_ASAP7_75t_L g1124 ( .A1(n_1080), .A2(n_1061), .A3(n_1092), .B(n_1076), .Y(n_1124) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1062), .Y(n_1125) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1066), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_1098), .B(n_1039), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1110), .B(n_1058), .Y(n_1128) );
INVx2_ASAP7_75t_L g1129 ( .A(n_1102), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1109), .Y(n_1130) );
INVx2_ASAP7_75t_SL g1131 ( .A(n_1099), .Y(n_1131) );
OAI32xp33_ASAP7_75t_L g1132 ( .A1(n_1113), .A2(n_1078), .A3(n_1084), .B1(n_1057), .B2(n_1069), .Y(n_1132) );
OAI332xp33_ASAP7_75t_L g1133 ( .A1(n_1119), .A2(n_1095), .A3(n_999), .B1(n_997), .B2(n_1023), .B3(n_1082), .C1(n_1085), .C2(n_1087), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1118), .B(n_1058), .Y(n_1134) );
INVx1_ASAP7_75t_SL g1135 ( .A(n_1113), .Y(n_1135) );
OAI32xp33_ASAP7_75t_L g1136 ( .A1(n_1111), .A2(n_1057), .A3(n_1069), .B1(n_1065), .B2(n_1075), .Y(n_1136) );
NAND2xp5_ASAP7_75t_SL g1137 ( .A(n_1124), .B(n_1056), .Y(n_1137) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1102), .Y(n_1138) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1125), .Y(n_1139) );
INVx2_ASAP7_75t_SL g1140 ( .A(n_1105), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1112), .Y(n_1141) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_1106), .A2(n_1070), .B1(n_1088), .B2(n_1055), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_1123), .A2(n_1046), .B1(n_1044), .B2(n_995), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1112), .Y(n_1144) );
OAI321xp33_ASAP7_75t_L g1145 ( .A1(n_1122), .A2(n_1002), .A3(n_1096), .B1(n_1093), .B2(n_1090), .C(n_1075), .Y(n_1145) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_1111), .B(n_1065), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1114), .Y(n_1147) );
AOI21xp5_ASAP7_75t_L g1148 ( .A1(n_1137), .A2(n_1116), .B(n_1103), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1146), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1146), .Y(n_1150) );
OAI31xp33_ASAP7_75t_L g1151 ( .A1(n_1137), .A2(n_1115), .A3(n_1120), .B(n_1107), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1130), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1141), .Y(n_1153) );
AOI322xp5_ASAP7_75t_L g1154 ( .A1(n_1135), .A2(n_1100), .A3(n_1101), .B1(n_1117), .B2(n_1108), .C1(n_1121), .C2(n_1115), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1144), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_1131), .A2(n_1070), .B1(n_1105), .B2(n_1107), .Y(n_1156) );
INVx2_ASAP7_75t_SL g1157 ( .A(n_1131), .Y(n_1157) );
NOR2xp33_ASAP7_75t_L g1158 ( .A(n_1133), .B(n_1097), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1147), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1134), .Y(n_1160) );
AOI222xp33_ASAP7_75t_L g1161 ( .A1(n_1127), .A2(n_1104), .B1(n_1097), .B2(n_1121), .C1(n_1117), .C2(n_1009), .Y(n_1161) );
AOI21xp33_ASAP7_75t_L g1162 ( .A1(n_1158), .A2(n_1145), .B(n_1143), .Y(n_1162) );
AOI22xp5_ASAP7_75t_L g1163 ( .A1(n_1161), .A2(n_1142), .B1(n_1143), .B2(n_1140), .Y(n_1163) );
O2A1O1Ixp33_ASAP7_75t_L g1164 ( .A1(n_1148), .A2(n_1132), .B(n_1136), .C(n_1128), .Y(n_1164) );
OAI221xp5_ASAP7_75t_L g1165 ( .A1(n_1151), .A2(n_1139), .B1(n_1138), .B2(n_1129), .C(n_1000), .Y(n_1165) );
NAND2xp5_ASAP7_75t_SL g1166 ( .A(n_1157), .B(n_1070), .Y(n_1166) );
NAND5xp2_ASAP7_75t_L g1167 ( .A(n_1154), .B(n_990), .C(n_986), .D(n_1017), .E(n_998), .Y(n_1167) );
AOI21xp33_ASAP7_75t_SL g1168 ( .A1(n_1156), .A2(n_1047), .B(n_927), .Y(n_1168) );
AOI21xp33_ASAP7_75t_SL g1169 ( .A1(n_1149), .A2(n_1047), .B(n_927), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_1162), .A2(n_1160), .B1(n_1150), .B2(n_1089), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1163), .Y(n_1171) );
BUFx6f_ASAP7_75t_L g1172 ( .A(n_1166), .Y(n_1172) );
AOI221xp5_ASAP7_75t_L g1173 ( .A1(n_1164), .A2(n_1159), .B1(n_1152), .B2(n_1155), .C(n_1153), .Y(n_1173) );
NOR4xp25_ASAP7_75t_L g1174 ( .A(n_1171), .B(n_1165), .C(n_1166), .D(n_969), .Y(n_1174) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_1170), .A2(n_1168), .B1(n_1169), .B2(n_1167), .Y(n_1175) );
NOR3x2_ASAP7_75t_L g1176 ( .A(n_1173), .B(n_950), .C(n_1091), .Y(n_1176) );
CKINVDCx6p67_ASAP7_75t_R g1177 ( .A(n_1172), .Y(n_1177) );
NAND4xp25_ASAP7_75t_L g1178 ( .A(n_1175), .B(n_950), .C(n_1172), .D(n_969), .Y(n_1178) );
INVx2_ASAP7_75t_L g1179 ( .A(n_1177), .Y(n_1179) );
AO22x2_ASAP7_75t_L g1180 ( .A1(n_1176), .A2(n_969), .B1(n_965), .B2(n_1125), .Y(n_1180) );
HB1xp67_ASAP7_75t_L g1181 ( .A(n_1179), .Y(n_1181) );
OR3x1_ASAP7_75t_L g1182 ( .A(n_1178), .B(n_1174), .C(n_981), .Y(n_1182) );
INVx2_ASAP7_75t_L g1183 ( .A(n_1181), .Y(n_1183) );
OAI22x1_ASAP7_75t_L g1184 ( .A1(n_1183), .A2(n_1182), .B1(n_1180), .B2(n_965), .Y(n_1184) );
OAI22xp33_ASAP7_75t_L g1185 ( .A1(n_1184), .A2(n_948), .B1(n_1091), .B2(n_1126), .Y(n_1185) );
OAI22xp33_ASAP7_75t_L g1186 ( .A1(n_1185), .A2(n_993), .B1(n_970), .B2(n_953), .Y(n_1186) );
AOI21xp5_ASAP7_75t_L g1187 ( .A1(n_1186), .A2(n_993), .B(n_953), .Y(n_1187) );
endmodule