module fake_jpeg_23759_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx4f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_3),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_14),
.B(n_16),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g15 ( 
.A1(n_9),
.A2(n_4),
.B(n_5),
.C(n_2),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_5),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_19),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_5),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_2),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_21),
.Y(n_25)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_27),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_10),
.B1(n_8),
.B2(n_13),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_28),
.B1(n_27),
.B2(n_29),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_14),
.C(n_16),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.C(n_35),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_8),
.C(n_20),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_16),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_22),
.C(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_40),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_17),
.C(n_6),
.Y(n_40)
);

OAI221xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.C(n_36),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_43),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_6),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_42),
.C(n_6),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_0),
.C(n_1),
.Y(n_46)
);


endmodule