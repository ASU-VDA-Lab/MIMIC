module fake_jpeg_21290_n_88 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_88);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_5),
.B(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_1),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_21),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_22),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_16),
.C(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_23),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_51),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_31),
.B1(n_29),
.B2(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_49),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_13),
.B1(n_19),
.B2(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_29),
.B1(n_15),
.B2(n_32),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_20),
.B1(n_32),
.B2(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_52),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_16),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_54),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

OR2x4_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_65),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_1),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_51),
.B1(n_43),
.B2(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_59),
.C(n_61),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_56),
.Y(n_71)
);

AOI221xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_64),
.B1(n_57),
.B2(n_55),
.C(n_18),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_62),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_42),
.B1(n_49),
.B2(n_48),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_73),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_9),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_79),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_72),
.B1(n_71),
.B2(n_20),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_80),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_7),
.B(n_2),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_78),
.B1(n_81),
.B2(n_8),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_84),
.Y(n_88)
);


endmodule