module fake_jpeg_16066_n_85 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_85);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_85;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx6_ASAP7_75t_SL g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_24),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_1),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_27),
.C(n_19),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_17),
.B1(n_10),
.B2(n_13),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_36),
.B1(n_14),
.B2(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_27),
.Y(n_39)
);

CKINVDCx12_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_37),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_10),
.B1(n_19),
.B2(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_27),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_10),
.B1(n_11),
.B2(n_16),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_46),
.B(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_47),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_25),
.B(n_21),
.C(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_14),
.B1(n_15),
.B2(n_20),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_18),
.Y(n_56)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_20),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_50),
.B(n_46),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_40),
.C(n_38),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_21),
.C(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_57),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_46),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_62),
.B(n_63),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_55),
.C(n_49),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_46),
.Y(n_62)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_51),
.B1(n_50),
.B2(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_SL g71 ( 
.A(n_67),
.B(n_62),
.C(n_61),
.Y(n_71)
);

FAx1_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_18),
.CI(n_28),
.CON(n_69),
.SN(n_69)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_69),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_34),
.C(n_7),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_66),
.C(n_67),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_34),
.C(n_9),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_77),
.B(n_34),
.Y(n_79)
);

AOI322xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_72),
.A3(n_71),
.B1(n_70),
.B2(n_8),
.C1(n_9),
.C2(n_6),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_79),
.C(n_80),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_76),
.B(n_5),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_4),
.C(n_5),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_82),
.B1(n_4),
.B2(n_6),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_4),
.Y(n_85)
);


endmodule