module real_jpeg_24170_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_1),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_1),
.A2(n_34),
.B1(n_51),
.B2(n_52),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_1),
.A2(n_34),
.B1(n_65),
.B2(n_66),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_46),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_2),
.A2(n_46),
.B1(n_65),
.B2(n_66),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_31),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_4),
.A2(n_37),
.B1(n_51),
.B2(n_52),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_4),
.A2(n_37),
.B1(n_65),
.B2(n_66),
.Y(n_136)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_7),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_69),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_69),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_8),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_145),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_8),
.A2(n_51),
.B1(n_52),
.B2(n_145),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_145),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_9),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_9),
.A2(n_65),
.B1(n_66),
.B2(n_147),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_147),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_147),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_10),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_10),
.B(n_101),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_10),
.B(n_61),
.C(n_65),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_10),
.B(n_57),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_10),
.A2(n_88),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_12),
.A2(n_115),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_12),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_154),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_12),
.A2(n_51),
.B1(n_52),
.B2(n_154),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_154),
.Y(n_224)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_15),
.Y(n_167)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_15),
.Y(n_217)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_15),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_121),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_102),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_19),
.B(n_102),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_72),
.C(n_84),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_20),
.A2(n_72),
.B1(n_73),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_20),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_42),
.B2(n_71),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_21),
.A2(n_22),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_22),
.B(n_43),
.C(n_70),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_35),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_23),
.A2(n_97),
.B1(n_152),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_25),
.B1(n_33),
.B2(n_38),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_24),
.A2(n_27),
.B(n_149),
.C(n_169),
.Y(n_168)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_25),
.B(n_26),
.C(n_31),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_26),
.A2(n_27),
.B1(n_50),
.B2(n_53),
.Y(n_54)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

HAxp5_ASAP7_75t_SL g242 ( 
.A(n_27),
.B(n_150),
.CON(n_242),
.SN(n_242)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_27),
.B(n_51),
.C(n_53),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_29),
.Y(n_113)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

HAxp5_ASAP7_75t_SL g149 ( 
.A(n_31),
.B(n_150),
.CON(n_149),
.SN(n_149)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_33),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_36),
.B(n_101),
.Y(n_100)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_40),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_40),
.A2(n_101),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_40),
.A2(n_101),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_40),
.A2(n_101),
.B1(n_160),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_58),
.B2(n_70),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_55),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_47),
.A2(n_109),
.B(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_47),
.A2(n_49),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_47),
.A2(n_55),
.B(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_57),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_48),
.B(n_56),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_48),
.A2(n_57),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_48),
.A2(n_57),
.B1(n_179),
.B2(n_242),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_49),
.A2(n_76),
.B(n_111),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_50),
.A2(n_52),
.B(n_242),
.C(n_243),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_52),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_52),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_57),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_70),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B(n_67),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_59),
.A2(n_67),
.B(n_94),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_59),
.A2(n_64),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_59),
.A2(n_64),
.B1(n_199),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_59),
.A2(n_79),
.B(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_59),
.A2(n_64),
.B1(n_93),
.B2(n_138),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_64),
.A2(n_81),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_64),
.B(n_150),
.Y(n_233)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_66),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_73),
.A2(n_74),
.B(n_78),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_80),
.A2(n_83),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_84),
.B(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_95),
.B(n_96),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_85),
.A2(n_86),
.B1(n_320),
.B2(n_322),
.Y(n_319)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_87),
.A2(n_92),
.B1(n_95),
.B2(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_87),
.A2(n_95),
.B1(n_96),
.B2(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_90),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_88),
.A2(n_131),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_88),
.B(n_136),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_88),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_88),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_88),
.A2(n_167),
.B1(n_215),
.B2(n_224),
.Y(n_234)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_89),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_91),
.B(n_185),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_91),
.A2(n_133),
.B(n_213),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_92),
.Y(n_302)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_96),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_100),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_97),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_99),
.B(n_101),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_118),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_110),
.Y(n_286)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_327),
.B(n_332),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_314),
.B(n_326),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_297),
.B(n_313),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_187),
.B(n_274),
.C(n_296),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_171),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_126),
.B(n_171),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_155),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_139),
.B2(n_140),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_128),
.B(n_140),
.C(n_155),
.Y(n_275)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_130),
.B(n_137),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.C(n_148),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_150),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_163),
.B2(n_170),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_158),
.B(n_161),
.C(n_170),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_168),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.C(n_176),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_172),
.B(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_175),
.B(n_176),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_183),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_177),
.B(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_259)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_186),
.B(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_273),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_268),
.B(n_272),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_254),
.B(n_267),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_238),
.B(n_253),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_210),
.B(n_237),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_200),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_200),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_194),
.A2(n_196),
.B1(n_197),
.B2(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_205),
.C(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_206),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_208),
.Y(n_218)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_221),
.B(n_236),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_219),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_218),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_232),
.B(n_235),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_233),
.B(n_234),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_252),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_252),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_247),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_248),
.C(n_251),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_244),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_250),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_256),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_263),
.C(n_265),
.Y(n_271)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_271),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_276),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_295),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_287),
.B1(n_293),
.B2(n_294),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_282),
.C(n_284),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_283),
.Y(n_307)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_293),
.C(n_295),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_292),
.Y(n_310)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_298),
.B(n_299),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_312),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_303),
.C(n_312),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_310),
.B2(n_311),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_309),
.C(n_311),
.Y(n_325)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_316),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_325),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_323),
.B2(n_324),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_323),
.C(n_325),
.Y(n_328)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_320),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);


endmodule