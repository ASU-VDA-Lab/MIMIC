module real_jpeg_28907_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_334, n_335, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_334;
input n_335;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_0),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_0),
.A2(n_26),
.B1(n_50),
.B2(n_52),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_0),
.A2(n_26),
.B1(n_55),
.B2(n_56),
.Y(n_265)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_1),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_3),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_108),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_108),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_3),
.A2(n_50),
.B1(n_52),
.B2(n_108),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_4),
.A2(n_43),
.B1(n_50),
.B2(n_52),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_258)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_6),
.A2(n_36),
.B1(n_55),
.B2(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_6),
.A2(n_36),
.B1(n_50),
.B2(n_52),
.Y(n_155)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_8),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_98),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_8),
.A2(n_50),
.B1(n_52),
.B2(n_98),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_98),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_9),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_9),
.A2(n_45),
.B1(n_55),
.B2(n_56),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_10),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_28),
.B(n_32),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_10),
.B(n_30),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_55),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_10),
.B(n_55),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_10),
.B(n_69),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_10),
.A2(n_118),
.B1(n_135),
.B2(n_201),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_10),
.A2(n_31),
.B(n_216),
.Y(n_215)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_12),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_93),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_12),
.A2(n_50),
.B1(n_52),
.B2(n_93),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_93),
.Y(n_220)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_15),
.A2(n_55),
.B1(n_56),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_15),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_15),
.A2(n_50),
.B1(n_52),
.B2(n_101),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_101),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_101),
.Y(n_283)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_16),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_91),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_17),
.A2(n_55),
.B1(n_56),
.B2(n_91),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_17),
.A2(n_50),
.B1(n_52),
.B2(n_91),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_79),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_77),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_37),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_23),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_73)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_25),
.A2(n_34),
.B(n_105),
.C(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_27),
.A2(n_30),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_27),
.A2(n_30),
.B1(n_143),
.B2(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_27),
.A2(n_30),
.B1(n_162),
.B2(n_256),
.Y(n_255)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_30),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_31),
.A2(n_62),
.B(n_64),
.C(n_67),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_65),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_31),
.A2(n_56),
.A3(n_65),
.B1(n_217),
.B2(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_32),
.B(n_105),
.Y(n_217)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_70),
.C(n_72),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_38),
.A2(n_39),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_58),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_40),
.B(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_42),
.A2(n_74),
.B1(n_76),
.B2(n_283),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_46),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_46),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_46),
.A2(n_58),
.B1(n_309),
.B2(n_316),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_57),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_47),
.A2(n_53),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_47),
.A2(n_53),
.B1(n_133),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_47),
.A2(n_53),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_47),
.A2(n_53),
.B1(n_176),
.B2(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_47),
.B(n_105),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_47),
.A2(n_53),
.B1(n_97),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_47),
.A2(n_53),
.B1(n_57),
.B2(n_265),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_48),
.A2(n_52),
.A3(n_55),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_49),
.B(n_50),
.Y(n_180)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_50),
.B(n_206),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_55),
.B(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_58),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_60),
.A2(n_69),
.B1(n_90),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_60),
.A2(n_69),
.B1(n_146),
.B2(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_60),
.A2(n_69),
.B1(n_164),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_67),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_67),
.B1(n_89),
.B2(n_92),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_61),
.A2(n_67),
.B1(n_92),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_61),
.A2(n_67),
.B1(n_124),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_61),
.A2(n_67),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_65),
.Y(n_226)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_68),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_70),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_74),
.A2(n_76),
.B1(n_107),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_74),
.A2(n_76),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_324),
.B(n_330),
.Y(n_79)
);

OAI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_300),
.A3(n_319),
.B1(n_322),
.B2(n_323),
.C(n_334),
.Y(n_80)
);

AOI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_252),
.A3(n_289),
.B1(n_294),
.B2(n_299),
.C(n_335),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_148),
.C(n_166),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_128),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_84),
.B(n_128),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_109),
.C(n_120),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_85),
.B(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_103),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_94),
.B2(n_95),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_95),
.C(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_99),
.A2(n_102),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_99),
.A2(n_102),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_105),
.B(n_118),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_109),
.A2(n_120),
.B1(n_121),
.B2(n_250),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_109),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_112),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_113),
.A2(n_114),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_135),
.B1(n_137),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_118),
.A2(n_135),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_118),
.A2(n_135),
.B1(n_195),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_118),
.A2(n_135),
.B1(n_190),
.B2(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_118),
.A2(n_135),
.B(n_155),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.C(n_127),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_122),
.B(n_237),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_125),
.B(n_127),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_126),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_138),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_138),
.C(n_139),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_134),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_147),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_144),
.C(n_147),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_149),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_150),
.B(n_151),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_165),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_153),
.B(n_158),
.C(n_165),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_154),
.B(n_156),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_157),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_246),
.B(n_251),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_232),
.B(n_245),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_210),
.B(n_231),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_191),
.B(n_209),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_181),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_181),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_186),
.C(n_188),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_187),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_189),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_198),
.B(n_208),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_193),
.B(n_197),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_203),
.B(n_207),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_200),
.B(n_202),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_211),
.B(n_212),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_223),
.B1(n_229),
.B2(n_230),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_222),
.C(n_230),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_234),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_241),
.C(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_241),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_248),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_269),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_253),
.B(n_269),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_260),
.C(n_268),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_260),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_254),
.Y(n_331)
);

FAx1_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.CI(n_259),
.CON(n_254),
.SN(n_254)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_257),
.C(n_259),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_256),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_258),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_266),
.B2(n_267),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_261),
.B(n_267),
.Y(n_285)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_267),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_266),
.A2(n_281),
.B(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_287),
.B2(n_288),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_278),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_278),
.C(n_288),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_276),
.B(n_277),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_276),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_275),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_302),
.C(n_311),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g321 ( 
.A(n_277),
.B(n_302),
.CI(n_311),
.CON(n_321),
.SN(n_321)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_278)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_295),
.B(n_298),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_291),
.B(n_292),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_312),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_312),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_310),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_304),
.B1(n_314),
.B2(n_317),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_306),
.C(n_309),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_317),
.C(n_318),
.Y(n_325)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_318),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_321),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_321),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);


endmodule