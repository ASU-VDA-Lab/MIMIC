module real_aes_1717_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_103;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_0), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_1), .B(n_188), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_2), .B(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g146 ( .A(n_3), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_4), .B(n_522), .Y(n_521) );
NAND2xp33_ASAP7_75t_SL g603 ( .A(n_5), .B(n_175), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_6), .B(n_155), .Y(n_179) );
INVx1_ASAP7_75t_L g596 ( .A(n_7), .Y(n_596) );
INVx1_ASAP7_75t_L g201 ( .A(n_8), .Y(n_201) );
CKINVDCx16_ASAP7_75t_R g827 ( .A(n_9), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_10), .Y(n_217) );
AND2x2_ASAP7_75t_L g519 ( .A(n_11), .B(n_232), .Y(n_519) );
INVx2_ASAP7_75t_L g154 ( .A(n_12), .Y(n_154) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_13), .Y(n_115) );
AND3x1_ASAP7_75t_L g824 ( .A(n_13), .B(n_36), .C(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g189 ( .A(n_14), .Y(n_189) );
AOI221x1_ASAP7_75t_L g599 ( .A1(n_15), .A2(n_206), .B1(n_524), .B2(n_600), .C(n_602), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_16), .B(n_522), .Y(n_583) );
INVx1_ASAP7_75t_L g119 ( .A(n_17), .Y(n_119) );
INVx1_ASAP7_75t_L g186 ( .A(n_18), .Y(n_186) );
INVx1_ASAP7_75t_SL g261 ( .A(n_19), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_20), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_21), .B(n_166), .Y(n_165) );
AOI33xp33_ASAP7_75t_L g238 ( .A1(n_22), .A2(n_51), .A3(n_143), .B1(n_161), .B2(n_239), .B3(n_240), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_23), .A2(n_524), .B(n_525), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_24), .B(n_188), .Y(n_526) );
AOI221xp5_ASAP7_75t_SL g570 ( .A1(n_25), .A2(n_41), .B1(n_522), .B2(n_524), .C(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g210 ( .A(n_26), .Y(n_210) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_27), .A2(n_91), .B(n_154), .Y(n_153) );
OR2x2_ASAP7_75t_L g156 ( .A(n_27), .B(n_91), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_28), .B(n_191), .Y(n_587) );
INVxp67_ASAP7_75t_L g598 ( .A(n_29), .Y(n_598) );
AND2x2_ASAP7_75t_L g545 ( .A(n_30), .B(n_231), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_31), .B(n_199), .Y(n_258) );
INVxp33_ASAP7_75t_L g829 ( .A(n_32), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_33), .A2(n_524), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_34), .B(n_191), .Y(n_572) );
AND2x2_ASAP7_75t_L g149 ( .A(n_35), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g160 ( .A(n_35), .Y(n_160) );
AND2x2_ASAP7_75t_L g175 ( .A(n_35), .B(n_146), .Y(n_175) );
OR2x6_ASAP7_75t_L g117 ( .A(n_36), .B(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_37), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_38), .B(n_199), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_39), .A2(n_140), .B1(n_152), .B2(n_155), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_40), .B(n_172), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_42), .A2(n_81), .B1(n_158), .B2(n_524), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_43), .B(n_166), .Y(n_262) );
AOI22xp5_ASAP7_75t_SL g123 ( .A1(n_44), .A2(n_71), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_44), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_45), .B(n_188), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_46), .B(n_177), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_47), .B(n_166), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_48), .Y(n_151) );
AND2x2_ASAP7_75t_L g563 ( .A(n_49), .B(n_231), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_50), .B(n_231), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_52), .B(n_166), .Y(n_229) );
INVx1_ASAP7_75t_L g144 ( .A(n_53), .Y(n_144) );
INVx1_ASAP7_75t_L g168 ( .A(n_53), .Y(n_168) );
AND2x2_ASAP7_75t_L g230 ( .A(n_54), .B(n_231), .Y(n_230) );
AOI221xp5_ASAP7_75t_L g198 ( .A1(n_55), .A2(n_74), .B1(n_158), .B2(n_199), .C(n_200), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_56), .B(n_199), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_57), .B(n_522), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_58), .B(n_152), .Y(n_219) );
AOI21xp5_ASAP7_75t_SL g249 ( .A1(n_59), .A2(n_158), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g536 ( .A(n_60), .B(n_231), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_61), .B(n_191), .Y(n_561) );
INVx1_ASAP7_75t_L g182 ( .A(n_62), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_63), .B(n_188), .Y(n_534) );
AND2x2_ASAP7_75t_SL g588 ( .A(n_64), .B(n_232), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_65), .A2(n_524), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g228 ( .A(n_66), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_67), .B(n_191), .Y(n_527) );
AND2x2_ASAP7_75t_SL g552 ( .A(n_68), .B(n_177), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_69), .A2(n_158), .B(n_227), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_70), .A2(n_89), .B1(n_506), .B2(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_70), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_71), .Y(n_124) );
INVx1_ASAP7_75t_L g150 ( .A(n_72), .Y(n_150) );
INVx1_ASAP7_75t_L g170 ( .A(n_72), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_73), .B(n_199), .Y(n_241) );
AND2x2_ASAP7_75t_L g263 ( .A(n_75), .B(n_206), .Y(n_263) );
INVx1_ASAP7_75t_L g183 ( .A(n_76), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_77), .A2(n_158), .B(n_260), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g157 ( .A1(n_78), .A2(n_158), .B(n_164), .C(n_176), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_79), .B(n_522), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_80), .A2(n_84), .B1(n_199), .B2(n_522), .Y(n_550) );
INVx1_ASAP7_75t_L g120 ( .A(n_82), .Y(n_120) );
AND2x2_ASAP7_75t_SL g247 ( .A(n_83), .B(n_206), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_85), .A2(n_158), .B1(n_236), .B2(n_237), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_86), .B(n_188), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_87), .B(n_188), .Y(n_573) );
OAI22xp5_ASAP7_75t_SL g809 ( .A1(n_88), .A2(n_810), .B1(n_811), .B2(n_813), .Y(n_809) );
INVx1_ASAP7_75t_L g813 ( .A(n_88), .Y(n_813) );
NOR3xp33_ASAP7_75t_L g132 ( .A(n_89), .B(n_133), .C(n_360), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_89), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_90), .A2(n_524), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g251 ( .A(n_92), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_93), .B(n_191), .Y(n_533) );
AND2x2_ASAP7_75t_L g242 ( .A(n_94), .B(n_206), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_95), .A2(n_208), .B(n_209), .C(n_211), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_96), .B(n_522), .Y(n_562) );
INVxp67_ASAP7_75t_L g601 ( .A(n_97), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_98), .B(n_191), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_99), .A2(n_524), .B(n_585), .Y(n_584) );
BUFx2_ASAP7_75t_L g107 ( .A(n_100), .Y(n_107) );
BUFx2_ASAP7_75t_SL g804 ( .A(n_100), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_101), .B(n_166), .Y(n_252) );
AOI21xp33_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_820), .B(n_828), .Y(n_102) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_122), .B(n_802), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_109), .A2(n_806), .B(n_817), .Y(n_805) );
NOR2xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_121), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g819 ( .A(n_114), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x6_ASAP7_75t_SL g130 ( .A(n_115), .B(n_117), .Y(n_130) );
OR2x6_ASAP7_75t_SL g511 ( .A(n_115), .B(n_116), .Y(n_511) );
OR2x2_ASAP7_75t_L g801 ( .A(n_115), .B(n_117), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g823 ( .A(n_118), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_126), .B(n_793), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_123), .A2(n_794), .B(n_797), .Y(n_793) );
INVxp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AO22x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_131), .B1(n_510), .B2(n_512), .Y(n_127) );
INVx4_ASAP7_75t_SL g795 ( .A(n_128), .Y(n_795) );
INVx3_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_131), .A2(n_512), .B1(n_795), .B2(n_796), .Y(n_794) );
AOI211x1_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_402), .B(n_503), .C(n_507), .Y(n_131) );
INVxp67_ASAP7_75t_L g505 ( .A(n_133), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_133), .B(n_447), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_307), .C(n_340), .Y(n_133) );
AOI211xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_264), .B(n_273), .C(n_297), .Y(n_134) );
OAI21xp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_193), .B(n_243), .Y(n_135) );
OR2x2_ASAP7_75t_L g317 ( .A(n_136), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g445 ( .A(n_136), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g429 ( .A(n_137), .B(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_137), .A2(n_450), .B1(n_453), .B2(n_454), .Y(n_449) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_178), .Y(n_137) );
INVx1_ASAP7_75t_L g296 ( .A(n_138), .Y(n_296) );
AND2x4_ASAP7_75t_L g313 ( .A(n_138), .B(n_294), .Y(n_313) );
INVx2_ASAP7_75t_L g335 ( .A(n_138), .Y(n_335) );
AND2x2_ASAP7_75t_L g383 ( .A(n_138), .B(n_246), .Y(n_383) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_138), .Y(n_397) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_157), .Y(n_138) );
NOR3xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_147), .C(n_151), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g199 ( .A(n_142), .B(n_148), .Y(n_199) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
OR2x6_ASAP7_75t_L g173 ( .A(n_143), .B(n_162), .Y(n_173) );
INVxp33_ASAP7_75t_L g239 ( .A(n_143), .Y(n_239) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g163 ( .A(n_144), .B(n_146), .Y(n_163) );
AND2x4_ASAP7_75t_L g191 ( .A(n_144), .B(n_169), .Y(n_191) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x6_ASAP7_75t_L g524 ( .A(n_149), .B(n_163), .Y(n_524) );
INVx2_ASAP7_75t_L g162 ( .A(n_150), .Y(n_162) );
AND2x6_ASAP7_75t_L g188 ( .A(n_150), .B(n_167), .Y(n_188) );
INVx4_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_152), .B(n_216), .Y(n_215) );
AOI21x1_ASAP7_75t_L g556 ( .A1(n_152), .A2(n_557), .B(n_563), .Y(n_556) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx4f_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
AND2x4_ASAP7_75t_L g155 ( .A(n_154), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_SL g232 ( .A(n_154), .B(n_156), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_155), .B(n_174), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_155), .A2(n_249), .B(n_253), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_155), .A2(n_521), .B(n_523), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_155), .B(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_155), .B(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_155), .B(n_601), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_155), .B(n_184), .C(n_603), .Y(n_602) );
INVxp67_ASAP7_75t_L g218 ( .A(n_158), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_158), .A2(n_199), .B1(n_595), .B2(n_597), .Y(n_594) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_163), .Y(n_158) );
NOR2x1p5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx1_ASAP7_75t_L g240 ( .A(n_161), .Y(n_240) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_171), .B(n_174), .Y(n_164) );
INVx1_ASAP7_75t_L g184 ( .A(n_166), .Y(n_184) );
AND2x4_ASAP7_75t_L g522 ( .A(n_166), .B(n_175), .Y(n_522) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_169), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g181 ( .A1(n_173), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_SL g200 ( .A1(n_173), .A2(n_174), .B(n_201), .C(n_202), .Y(n_200) );
INVxp67_ASAP7_75t_L g208 ( .A(n_173), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_173), .A2(n_174), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_173), .A2(n_174), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_SL g260 ( .A1(n_173), .A2(n_174), .B(n_261), .C(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g236 ( .A(n_174), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_174), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_174), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_174), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_174), .A2(n_560), .B(n_561), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_174), .A2(n_572), .B(n_573), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_174), .A2(n_586), .B(n_587), .Y(n_585) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_175), .Y(n_211) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_176), .A2(n_234), .B(n_242), .Y(n_233) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_176), .A2(n_234), .B(n_242), .Y(n_278) );
AOI21x1_ASAP7_75t_L g548 ( .A1(n_176), .A2(n_549), .B(n_552), .Y(n_548) );
INVx2_ASAP7_75t_SL g176 ( .A(n_177), .Y(n_176) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_177), .A2(n_198), .B(n_203), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_177), .A2(n_583), .B(n_584), .Y(n_582) );
AND2x2_ASAP7_75t_L g254 ( .A(n_178), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g283 ( .A(n_178), .Y(n_283) );
INVx3_ASAP7_75t_L g294 ( .A(n_178), .Y(n_294) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_185), .B(n_192), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_184), .B(n_210), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B1(n_189), .B2(n_190), .Y(n_185) );
INVxp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVxp67_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_193), .A2(n_378), .B1(n_380), .B2(n_382), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_193), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_221), .Y(n_194) );
INVx3_ASAP7_75t_L g267 ( .A(n_195), .Y(n_267) );
AND2x2_ASAP7_75t_L g275 ( .A(n_195), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_195), .Y(n_305) );
NAND2x1_ASAP7_75t_SL g394 ( .A(n_195), .B(n_266), .Y(n_394) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_204), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g272 ( .A(n_197), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_197), .B(n_278), .Y(n_290) );
AND2x2_ASAP7_75t_L g303 ( .A(n_197), .B(n_204), .Y(n_303) );
AND2x4_ASAP7_75t_L g310 ( .A(n_197), .B(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_197), .Y(n_359) );
INVx1_ASAP7_75t_L g369 ( .A(n_197), .Y(n_369) );
INVxp67_ASAP7_75t_L g452 ( .A(n_197), .Y(n_452) );
INVx1_ASAP7_75t_L g220 ( .A(n_199), .Y(n_220) );
INVx1_ASAP7_75t_L g270 ( .A(n_204), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_204), .B(n_280), .Y(n_289) );
INVx2_ASAP7_75t_L g357 ( .A(n_204), .Y(n_357) );
INVx1_ASAP7_75t_L g400 ( .A(n_204), .Y(n_400) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_214), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B1(n_212), .B2(n_213), .Y(n_205) );
INVx3_ASAP7_75t_L g213 ( .A(n_206), .Y(n_213) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_213), .A2(n_224), .B(n_230), .Y(n_223) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_213), .A2(n_224), .B(n_230), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_218), .B1(n_219), .B2(n_220), .Y(n_214) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g326 ( .A(n_221), .B(n_303), .Y(n_326) );
AND2x2_ASAP7_75t_L g475 ( .A(n_221), .B(n_399), .Y(n_475) );
AND2x2_ASAP7_75t_L g481 ( .A(n_221), .B(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_221), .B(n_442), .Y(n_492) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_233), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NOR2x1_ASAP7_75t_L g271 ( .A(n_223), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g418 ( .A(n_223), .B(n_357), .Y(n_418) );
AND2x2_ASAP7_75t_L g422 ( .A(n_223), .B(n_277), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_231), .Y(n_256) );
OA21x2_ASAP7_75t_L g569 ( .A1(n_231), .A2(n_570), .B(n_574), .Y(n_569) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g266 ( .A(n_233), .Y(n_266) );
INVx2_ASAP7_75t_L g311 ( .A(n_233), .Y(n_311) );
AND2x2_ASAP7_75t_L g356 ( .A(n_233), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_235), .B(n_241), .Y(n_234) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_254), .Y(n_244) );
OR2x6_ASAP7_75t_L g424 ( .A(n_245), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g428 ( .A(n_245), .B(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx4_ASAP7_75t_L g287 ( .A(n_246), .Y(n_287) );
AND2x4_ASAP7_75t_L g295 ( .A(n_246), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g330 ( .A(n_246), .B(n_255), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_246), .B(n_353), .Y(n_376) );
AND2x2_ASAP7_75t_L g392 ( .A(n_246), .B(n_283), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_246), .B(n_348), .Y(n_446) );
INVx2_ASAP7_75t_L g461 ( .A(n_246), .Y(n_461) );
OR2x6_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x2_ASAP7_75t_L g306 ( .A(n_254), .B(n_295), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_254), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_SL g410 ( .A(n_254), .B(n_333), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_254), .B(n_346), .Y(n_439) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_255), .Y(n_285) );
AND2x2_ASAP7_75t_L g293 ( .A(n_255), .B(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_255), .Y(n_316) );
INVx2_ASAP7_75t_L g319 ( .A(n_255), .Y(n_319) );
INVx1_ASAP7_75t_L g352 ( .A(n_255), .Y(n_352) );
INVx1_ASAP7_75t_L g430 ( .A(n_255), .Y(n_430) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_263), .Y(n_255) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_256), .A2(n_530), .B(n_536), .Y(n_529) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_256), .A2(n_539), .B(n_545), .Y(n_538) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_256), .A2(n_539), .B(n_545), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_266), .B(n_269), .Y(n_342) );
AND4x1_ASAP7_75t_SL g432 ( .A(n_266), .B(n_407), .C(n_433), .D(n_435), .Y(n_432) );
OR2x2_ASAP7_75t_L g486 ( .A(n_266), .B(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g378 ( .A(n_267), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AND2x2_ASAP7_75t_L g321 ( .A(n_270), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_270), .B(n_279), .Y(n_444) );
AND2x2_ASAP7_75t_L g390 ( .A(n_271), .B(n_356), .Y(n_390) );
OAI32xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_281), .A3(n_286), .B1(n_288), .B2(n_291), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g441 ( .A(n_276), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g454 ( .A(n_276), .B(n_372), .Y(n_454) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g417 ( .A(n_277), .Y(n_417) );
AND2x2_ASAP7_75t_L g451 ( .A(n_277), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_278), .B(n_280), .Y(n_379) );
INVx3_ASAP7_75t_L g302 ( .A(n_279), .Y(n_302) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_279), .B(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_280), .Y(n_339) );
AND2x2_ASAP7_75t_L g358 ( .A(n_280), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g386 ( .A(n_282), .Y(n_386) );
NAND2x1_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g332 ( .A(n_283), .Y(n_332) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_283), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_286), .B(n_473), .Y(n_472) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g324 ( .A(n_287), .B(n_292), .Y(n_324) );
AND2x4_ASAP7_75t_L g346 ( .A(n_287), .B(n_296), .Y(n_346) );
AND2x4_ASAP7_75t_SL g396 ( .A(n_287), .B(n_397), .Y(n_396) );
NOR2x1_ASAP7_75t_L g408 ( .A(n_287), .B(n_364), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_288), .A2(n_484), .B1(n_486), .B2(n_488), .Y(n_483) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx2_ASAP7_75t_SL g496 ( .A(n_289), .Y(n_496) );
INVx2_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_293), .B(n_299), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_293), .A2(n_495), .B1(n_498), .B2(n_501), .Y(n_497) );
INVx1_ASAP7_75t_L g353 ( .A(n_294), .Y(n_353) );
AND2x2_ASAP7_75t_L g426 ( .A(n_294), .B(n_335), .Y(n_426) );
INVx2_ASAP7_75t_L g299 ( .A(n_295), .Y(n_299) );
OAI21xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_300), .B(n_304), .Y(n_297) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_301), .A2(n_456), .B1(n_459), .B2(n_460), .Y(n_455) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_302), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_302), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g471 ( .A(n_302), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NOR3xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_323), .C(n_327), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_312), .B1(n_317), .B2(n_320), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g337 ( .A(n_310), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g398 ( .A(n_310), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g411 ( .A(n_310), .B(n_400), .Y(n_411) );
AND2x2_ASAP7_75t_L g459 ( .A(n_310), .B(n_418), .Y(n_459) );
AND2x2_ASAP7_75t_L g495 ( .A(n_310), .B(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx4_ASAP7_75t_L g364 ( .A(n_313), .Y(n_364) );
AND2x2_ASAP7_75t_L g460 ( .A(n_313), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_L g465 ( .A(n_316), .Y(n_465) );
AND2x2_ASAP7_75t_L g473 ( .A(n_316), .B(n_426), .Y(n_473) );
INVx1_ASAP7_75t_L g375 ( .A(n_318), .Y(n_375) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g348 ( .A(n_319), .Y(n_348) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_321), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_322), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_331), .B(n_336), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_329), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AOI21xp33_ASAP7_75t_SL g340 ( .A1(n_332), .A2(n_341), .B(n_343), .Y(n_340) );
AND2x2_ASAP7_75t_L g381 ( .A(n_332), .B(n_346), .Y(n_381) );
AND2x4_ASAP7_75t_L g350 ( .A(n_333), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_333), .B(n_430), .Y(n_438) );
INVx2_ASAP7_75t_SL g466 ( .A(n_333), .Y(n_466) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI21xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_349), .B(n_354), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_346), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_346), .B(n_351), .Y(n_494) );
AND2x2_ASAP7_75t_L g391 ( .A(n_347), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g395 ( .A(n_347), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g434 ( .A(n_347), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_347), .B(n_364), .Y(n_453) );
INVx1_ASAP7_75t_L g482 ( .A(n_347), .Y(n_482) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_SL g351 ( .A(n_352), .B(n_353), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_352), .B(n_426), .Y(n_458) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g366 ( .A(n_356), .Y(n_366) );
AND2x2_ASAP7_75t_L g372 ( .A(n_357), .B(n_369), .Y(n_372) );
INVxp67_ASAP7_75t_L g508 ( .A(n_360), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_360), .B(n_403), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_387), .Y(n_360) );
NOR3xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_377), .C(n_384), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B1(n_370), .B2(n_373), .Y(n_362) );
INVx2_ASAP7_75t_L g401 ( .A(n_364), .Y(n_401) );
NAND2xp5_ASAP7_75t_R g419 ( .A(n_364), .B(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx3_ASAP7_75t_L g415 ( .A(n_368), .Y(n_415) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g467 ( .A(n_371), .Y(n_467) );
INVx2_ASAP7_75t_L g487 ( .A(n_372), .Y(n_487) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_374), .A2(n_491), .B1(n_493), .B2(n_495), .Y(n_490) );
NOR2x1_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
NOR3xp33_ASAP7_75t_L g384 ( .A(n_378), .B(n_383), .C(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI222xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_391), .B1(n_393), .B2(n_395), .C1(n_398), .C2(n_401), .Y(n_387) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_392), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g420 ( .A(n_396), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_396), .B(n_465), .Y(n_488) );
INVx1_ASAP7_75t_L g442 ( .A(n_399), .Y(n_442) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_399), .A2(n_478), .B(n_479), .Y(n_477) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g421 ( .A(n_400), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g435 ( .A(n_400), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_447), .Y(n_402) );
INVxp67_ASAP7_75t_L g509 ( .A(n_403), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_412), .C(n_431), .Y(n_403) );
NOR2x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_419), .B1(n_421), .B2(n_423), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_L g480 ( .A(n_415), .Y(n_480) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
AND2x2_ASAP7_75t_L g450 ( .A(n_418), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_427), .Y(n_423) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_427), .A2(n_469), .B1(n_472), .B2(n_474), .Y(n_468) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g498 ( .A(n_430), .B(n_499), .Y(n_498) );
NOR3xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_436), .C(n_443), .Y(n_431) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g485 ( .A(n_434), .B(n_460), .Y(n_485) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B(n_440), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVxp67_ASAP7_75t_L g504 ( .A(n_447), .Y(n_504) );
NAND4xp75_ASAP7_75t_L g447 ( .A(n_448), .B(n_462), .C(n_476), .D(n_489), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_455), .Y(n_448) );
NAND2x1p5_ASAP7_75t_L g502 ( .A(n_451), .B(n_496), .Y(n_502) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g500 ( .A(n_461), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_467), .B(n_468), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_466), .B(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_481), .B(n_483), .Y(n_476) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_497), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B(n_506), .Y(n_503) );
AOI21xp5_ASAP7_75t_SL g507 ( .A1(n_506), .A2(n_508), .B(n_509), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_510), .Y(n_796) );
CKINVDCx11_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_723), .Y(n_513) );
NOR4xp25_ASAP7_75t_SL g514 ( .A(n_515), .B(n_616), .C(n_660), .D(n_687), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_579), .B1(n_589), .B2(n_604), .C(n_606), .Y(n_515) );
AOI32xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_546), .A3(n_553), .B1(n_564), .B2(n_575), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_517), .B(n_759), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_517), .A2(n_729), .B1(n_787), .B2(n_790), .Y(n_786) );
AND2x4_ASAP7_75t_SL g517 ( .A(n_518), .B(n_528), .Y(n_517) );
INVx5_ASAP7_75t_L g578 ( .A(n_518), .Y(n_578) );
OR2x2_ASAP7_75t_L g605 ( .A(n_518), .B(n_577), .Y(n_605) );
AND2x4_ASAP7_75t_L g607 ( .A(n_518), .B(n_538), .Y(n_607) );
INVx2_ASAP7_75t_L g622 ( .A(n_518), .Y(n_622) );
OR2x2_ASAP7_75t_L g634 ( .A(n_518), .B(n_547), .Y(n_634) );
AND2x2_ASAP7_75t_L g641 ( .A(n_518), .B(n_537), .Y(n_641) );
AND2x2_ASAP7_75t_SL g683 ( .A(n_518), .B(n_566), .Y(n_683) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_518), .Y(n_740) );
OR2x6_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx3_ASAP7_75t_SL g635 ( .A(n_528), .Y(n_635) );
AND2x2_ASAP7_75t_L g654 ( .A(n_528), .B(n_578), .Y(n_654) );
AOI32xp33_ASAP7_75t_L g769 ( .A1(n_528), .A2(n_640), .A3(n_670), .B1(n_700), .B2(n_735), .Y(n_769) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_537), .Y(n_528) );
AND2x2_ASAP7_75t_L g609 ( .A(n_529), .B(n_547), .Y(n_609) );
OR2x2_ASAP7_75t_L g625 ( .A(n_529), .B(n_538), .Y(n_625) );
INVx1_ASAP7_75t_L g648 ( .A(n_529), .Y(n_648) );
INVx2_ASAP7_75t_L g664 ( .A(n_529), .Y(n_664) );
AND2x2_ASAP7_75t_L g701 ( .A(n_529), .B(n_566), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_529), .B(n_538), .Y(n_720) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_529), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g756 ( .A(n_538), .B(n_547), .Y(n_756) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_538), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_544), .Y(n_539) );
OR2x2_ASAP7_75t_L g604 ( .A(n_546), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g610 ( .A(n_546), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g623 ( .A(n_546), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g785 ( .A(n_546), .B(n_654), .Y(n_785) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g714 ( .A(n_547), .B(n_664), .Y(n_714) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_548), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_553), .B(n_681), .Y(n_783) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_554), .B(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g568 ( .A(n_555), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g590 ( .A(n_555), .Y(n_590) );
AND2x2_ASAP7_75t_L g614 ( .A(n_555), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_555), .B(n_592), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_555), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g672 ( .A(n_555), .Y(n_672) );
OR2x2_ASAP7_75t_L g691 ( .A(n_555), .B(n_618), .Y(n_691) );
INVx1_ASAP7_75t_L g698 ( .A(n_555), .Y(n_698) );
NOR2xp33_ASAP7_75t_R g750 ( .A(n_555), .B(n_581), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_555), .B(n_593), .Y(n_754) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_562), .Y(n_557) );
AOI32xp33_ASAP7_75t_L g777 ( .A1(n_564), .A2(n_613), .A3(n_778), .B1(n_779), .B2(n_780), .Y(n_777) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx2_ASAP7_75t_L g644 ( .A(n_566), .Y(n_644) );
AND2x4_ASAP7_75t_L g663 ( .A(n_566), .B(n_664), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_566), .B(n_635), .Y(n_692) );
OR2x2_ASAP7_75t_L g746 ( .A(n_566), .B(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g704 ( .A(n_567), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g762 ( .A(n_567), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_568), .B(n_581), .Y(n_728) );
AND2x2_ASAP7_75t_L g765 ( .A(n_568), .B(n_731), .Y(n_765) );
INVx2_ASAP7_75t_L g615 ( .A(n_569), .Y(n_615) );
INVx2_ASAP7_75t_L g618 ( .A(n_569), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_569), .B(n_581), .Y(n_638) );
INVx1_ASAP7_75t_L g669 ( .A(n_569), .Y(n_669) );
OR2x2_ASAP7_75t_L g695 ( .A(n_569), .B(n_581), .Y(n_695) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_569), .Y(n_747) );
BUFx3_ASAP7_75t_L g776 ( .A(n_569), .Y(n_776) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g645 ( .A(n_576), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_576), .B(n_663), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_576), .B(n_734), .Y(n_733) );
AND2x4_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_577), .B(n_648), .Y(n_647) );
OAI21xp33_ASAP7_75t_L g677 ( .A1(n_577), .A2(n_644), .B(n_662), .Y(n_677) );
OAI32xp33_ASAP7_75t_L g699 ( .A1(n_578), .A2(n_700), .A3(n_702), .B1(n_704), .B2(n_706), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_578), .B(n_663), .Y(n_772) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g705 ( .A(n_580), .Y(n_705) );
NOR2x1p5_ASAP7_75t_L g775 ( .A(n_580), .B(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_L g591 ( .A(n_581), .B(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_SL g613 ( .A(n_581), .B(n_593), .Y(n_613) );
OR2x2_ASAP7_75t_L g617 ( .A(n_581), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g652 ( .A(n_581), .Y(n_652) );
AND2x2_ASAP7_75t_L g670 ( .A(n_581), .B(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g681 ( .A(n_581), .B(n_593), .Y(n_681) );
OR2x2_ASAP7_75t_L g743 ( .A(n_581), .B(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g760 ( .A(n_581), .B(n_691), .Y(n_760) );
INVx1_ASAP7_75t_L g792 ( .A(n_581), .Y(n_792) );
OR2x6_ASAP7_75t_L g581 ( .A(n_582), .B(n_588), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_590), .B(n_669), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_591), .B(n_703), .Y(n_702) );
AOI222xp33_ASAP7_75t_L g707 ( .A1(n_591), .A2(n_708), .B1(n_713), .B2(n_715), .C1(n_718), .C2(n_721), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_591), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g735 ( .A(n_591), .B(n_614), .Y(n_735) );
AND2x2_ASAP7_75t_L g697 ( .A(n_592), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g712 ( .A(n_592), .B(n_617), .Y(n_712) );
INVx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_593), .B(n_618), .Y(n_650) );
AND2x4_ASAP7_75t_L g671 ( .A(n_593), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g731 ( .A(n_593), .B(n_652), .Y(n_731) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_599), .Y(n_593) );
INVx1_ASAP7_75t_SL g611 ( .A(n_605), .Y(n_611) );
NAND2xp33_ASAP7_75t_SL g780 ( .A(n_605), .B(n_635), .Y(n_780) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B(n_610), .C(n_612), .Y(n_606) );
INVx2_ASAP7_75t_SL g657 ( .A(n_607), .Y(n_657) );
AND2x2_ASAP7_75t_L g661 ( .A(n_608), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_609), .B(n_657), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_609), .A2(n_647), .B(n_683), .C(n_684), .Y(n_682) );
AND2x2_ASAP7_75t_L g759 ( .A(n_609), .B(n_740), .Y(n_759) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x4_ASAP7_75t_L g658 ( .A(n_613), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g763 ( .A(n_613), .Y(n_763) );
OAI211xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B(n_626), .C(n_653), .Y(n_616) );
INVx2_ASAP7_75t_L g628 ( .A(n_617), .Y(n_628) );
OR2x2_ASAP7_75t_L g675 ( .A(n_617), .B(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_618), .Y(n_659) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_621), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g713 ( .A(n_621), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_621), .B(n_701), .Y(n_767) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI222xp33_ASAP7_75t_L g725 ( .A1(n_623), .A2(n_726), .B1(n_727), .B2(n_729), .C1(n_732), .C2(n_735), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_624), .A2(n_689), .B1(n_692), .B2(n_693), .C(n_699), .Y(n_688) );
AND2x2_ASAP7_75t_L g726 ( .A(n_624), .B(n_683), .Y(n_726) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp33_ASAP7_75t_SL g639 ( .A(n_625), .B(n_640), .Y(n_639) );
AOI221x1_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_631), .B1(n_636), .B2(n_639), .C(n_642), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
AND2x2_ASAP7_75t_L g779 ( .A(n_629), .B(n_717), .Y(n_779) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g637 ( .A(n_630), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
OAI32xp33_ASAP7_75t_L g745 ( .A1(n_635), .A2(n_676), .A3(n_746), .B1(n_748), .B2(n_752), .Y(n_745) );
OAI21xp33_ASAP7_75t_SL g764 ( .A1(n_636), .A2(n_765), .B(n_766), .Y(n_764) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B(n_649), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
OR2x2_ASAP7_75t_L g646 ( .A(n_644), .B(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g719 ( .A(n_644), .B(n_720), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_648), .A2(n_674), .B1(n_677), .B2(n_678), .C(n_682), .Y(n_673) );
INVx1_ASAP7_75t_L g749 ( .A(n_648), .Y(n_749) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_648), .Y(n_755) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
OAI21xp33_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B(n_658), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_657), .B(n_722), .Y(n_721) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_665), .B(n_673), .Y(n_660) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_664), .Y(n_734) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_667), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVxp67_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g686 ( .A(n_669), .Y(n_686) );
INVx1_ASAP7_75t_L g676 ( .A(n_671), .Y(n_676) );
AND2x2_ASAP7_75t_SL g685 ( .A(n_671), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_671), .B(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_671), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g690 ( .A(n_681), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_686), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_688), .B(n_707), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g703 ( .A(n_691), .Y(n_703) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_SL g717 ( .A(n_695), .Y(n_717) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_697), .B(n_775), .Y(n_774) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_698), .Y(n_711) );
BUFx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_709), .B(n_712), .Y(n_708) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g722 ( .A(n_714), .Y(n_722) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g741 ( .A(n_720), .Y(n_741) );
NOR4xp25_ASAP7_75t_L g723 ( .A(n_724), .B(n_757), .C(n_768), .D(n_781), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_736), .Y(n_724) );
O2A1O1Ixp33_ASAP7_75t_L g736 ( .A1(n_726), .A2(n_737), .B(n_742), .C(n_745), .Y(n_736) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_739), .B(n_741), .Y(n_738) );
OAI211xp5_ASAP7_75t_L g748 ( .A1(n_739), .A2(n_749), .B(n_750), .C(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
OAI21xp33_ASAP7_75t_SL g752 ( .A1(n_753), .A2(n_755), .B(n_756), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_SL g787 ( .A(n_756), .B(n_788), .Y(n_787) );
OAI221xp5_ASAP7_75t_SL g757 ( .A1(n_758), .A2(n_760), .B1(n_761), .B2(n_762), .C(n_764), .Y(n_757) );
INVx1_ASAP7_75t_SL g761 ( .A(n_759), .Y(n_761) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NAND3xp33_ASAP7_75t_SL g768 ( .A(n_769), .B(n_770), .C(n_777), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI21xp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_784), .B(n_786), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVxp33_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
INVx1_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .Y(n_802) );
INVx1_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
XNOR2x1_ASAP7_75t_L g807 ( .A(n_808), .B(n_814), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AND2x2_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_SL g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_822), .Y(n_831) );
AND2x2_ASAP7_75t_SL g822 ( .A(n_823), .B(n_824), .Y(n_822) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
endmodule