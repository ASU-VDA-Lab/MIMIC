module fake_jpeg_3104_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_63),
.Y(n_66)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_53),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_46),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_49),
.B1(n_53),
.B2(n_55),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_74),
.B1(n_63),
.B2(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_44),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_55),
.B(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_54),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_49),
.B1(n_55),
.B2(n_42),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_78),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_61),
.B1(n_50),
.B2(n_42),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_84),
.B1(n_3),
.B2(n_4),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_60),
.B(n_62),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_87),
.B(n_0),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_63),
.B1(n_46),
.B2(n_51),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_90),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_43),
.B1(n_45),
.B2(n_2),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_1),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_86),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_21),
.Y(n_100)
);

AO21x2_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_75),
.B(n_19),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_97),
.B(n_13),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_98),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_91),
.B1(n_8),
.B2(n_9),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_4),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_108),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_5),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_5),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_6),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_24),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_10),
.B(n_11),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_117),
.B(n_22),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_26),
.B1(n_40),
.B2(n_38),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_11),
.B(n_12),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_126),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_25),
.C(n_37),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_104),
.C(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_29),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_104),
.B1(n_110),
.B2(n_94),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_129),
.A2(n_118),
.B1(n_112),
.B2(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_128),
.Y(n_131)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

AOI221xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_139),
.B1(n_140),
.B2(n_120),
.C(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_14),
.B(n_41),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_121),
.C(n_122),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_133),
.Y(n_150)
);

OAI322xp33_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_112),
.A3(n_136),
.B1(n_140),
.B2(n_137),
.C1(n_135),
.C2(n_30),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_145),
.A2(n_129),
.B1(n_134),
.B2(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_147),
.B(n_139),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_151),
.B(n_145),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_154),
.B(n_152),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_142),
.Y(n_157)
);

AOI21x1_ASAP7_75t_SL g158 ( 
.A1(n_157),
.A2(n_150),
.B(n_144),
.Y(n_158)
);

AOI21x1_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_146),
.B(n_148),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_144),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_23),
.B1(n_27),
.B2(n_33),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_161),
.Y(n_162)
);


endmodule