module fake_ibex_1625_n_4963 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4963);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4963;

wire n_4557;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_3548;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_4204;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_962;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_3479;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_2343;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_4423;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3472;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_4801;
wire n_3639;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_4569;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_4567;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1306;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1960;
wire n_937;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_3565;
wire n_3883;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_2147;
wire n_2253;
wire n_4479;
wire n_3858;
wire n_4173;
wire n_1078;
wire n_4422;
wire n_1865;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_1653;
wire n_1375;
wire n_1118;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_3060;
wire n_4124;
wire n_971;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_3293;
wire n_2550;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_1108;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_1209;
wire n_3732;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_1121;
wire n_4823;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_4757;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_1042;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_1987;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_4374;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_1008;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_1210;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_1246;
wire n_4231;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_2361;
wire n_4128;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_3544;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_2046;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_4679;
wire n_1345;
wire n_4456;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_1471;
wire n_3441;
wire n_4559;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_2010;
wire n_2733;
wire n_3796;
wire n_1836;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_4321;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_4024;
wire n_3975;
wire n_3164;
wire n_1448;
wire n_3034;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_1967;
wire n_1095;
wire n_3834;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_4851;
wire n_1122;
wire n_3387;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_3428;
wire n_2427;
wire n_1127;
wire n_947;
wire n_1004;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_2422;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_972;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_3339;
wire n_3673;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_1340;
wire n_2562;
wire n_3269;
wire n_2223;
wire n_3876;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_4339;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3686;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_1517;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_977;
wire n_1895;
wire n_1860;
wire n_1763;
wire n_3912;
wire n_1607;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_933;
wire n_2221;
wire n_1774;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1021;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_4729;
wire n_1617;
wire n_2639;
wire n_3099;
wire n_1001;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_1017;
wire n_2049;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_4417;
wire n_1550;
wire n_1169;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1072;
wire n_2194;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_3096;
wire n_1278;
wire n_2059;
wire n_4730;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_4082;
wire n_4367;
wire n_3273;
wire n_950;
wire n_4282;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_4919;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_2871;
wire n_2764;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_985;
wire n_4611;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_1459;
wire n_4032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_995;
wire n_1303;
wire n_1994;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_946;
wire n_4895;
wire n_3354;
wire n_4069;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_2574;
wire n_1887;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_2228;
wire n_4474;
wire n_1518;
wire n_4350;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_1010;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_4911;
wire n_1329;
wire n_2409;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_3742;
wire n_3532;
wire n_4686;
wire n_4682;
wire n_2914;
wire n_1833;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_4733;
wire n_987;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_1166;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_4962;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_4644;
wire n_1012;
wire n_960;
wire n_4412;
wire n_4266;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_1230;
wire n_3622;
wire n_3857;
wire n_2357;
wire n_4354;
wire n_2937;
wire n_3728;
wire n_4401;
wire n_4727;
wire n_4296;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1033;
wire n_990;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_4539;
wire n_1205;
wire n_2969;
wire n_3550;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_1002;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_3789;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_984;
wire n_2978;
wire n_3502;
wire n_3935;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_4926;
wire n_4688;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_1930;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_969;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_3484;
wire n_2485;
wire n_4477;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_948;
wire n_3726;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_4491;
wire n_4672;
wire n_2421;
wire n_3237;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_4433;
wire n_3030;
wire n_4503;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_3221;
wire n_4511;
wire n_3210;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_1301;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_4610;
wire n_4067;
wire n_4393;
wire n_3777;
wire n_4553;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_2257;
wire n_4856;
wire n_1467;
wire n_3217;
wire n_2511;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_3633;
wire n_1731;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3788;
wire n_3448;
wire n_2076;
wire n_974;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_959;
wire n_1312;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_2829;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_965;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_936;
wire n_2176;
wire n_2805;
wire n_2319;
wire n_3757;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_3787;
wire n_3445;
wire n_2080;
wire n_2554;
wire n_1676;
wire n_1013;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_1014;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_3394;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_3488;
wire n_2832;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_2142;
wire n_3703;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_954;
wire n_4734;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_998;
wire n_1729;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_4579;
wire n_943;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1775;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_3074;
wire n_4640;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_2170;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_997;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_3350;
wire n_4873;
wire n_945;
wire n_3936;
wire n_1560;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_4636;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_4609;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_1011;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_2442;
wire n_1067;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_1331;
wire n_1223;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_1294;
wire n_1351;
wire n_1380;
wire n_3336;
wire n_1291;
wire n_3763;
wire n_4284;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_1662;
wire n_3443;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_1660;
wire n_4000;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_1962;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_2309;
wire n_2274;
wire n_3712;
wire n_2143;
wire n_4637;
wire n_4021;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_4643;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_1241;
wire n_2589;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_1238;
wire n_3959;
wire n_976;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_1644;
wire n_4586;
wire n_3860;
wire n_1871;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_1149;
wire n_4905;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_1261;
wire n_3327;
wire n_1114;
wire n_3647;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1018;
wire n_1669;
wire n_1885;
wire n_1989;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_1175;
wire n_4408;
wire n_1221;
wire n_3875;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_4565;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_1507;
wire n_1206;
wire n_3576;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_956;
wire n_4597;
wire n_1812;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_1798;
wire n_4562;
wire n_1584;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_941;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_3050;
wire n_2666;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_4516;
wire n_2913;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_4196;
wire n_2371;
wire n_3898;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_2671;
wire n_3296;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_3207;
wire n_953;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_3036;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_3332;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_3861;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_955;
wire n_2619;
wire n_2917;
wire n_2726;
wire n_3738;
wire n_1640;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_1355;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_4590;
wire n_4602;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_1780;
wire n_1091;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_1743;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_4883;
wire n_1079;
wire n_3559;
wire n_4943;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_3750;
wire n_3838;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_4159;
wire n_4372;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_3819;
wire n_3334;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_1233;
wire n_3653;
wire n_4360;
wire n_4897;
wire n_963;
wire n_2139;
wire n_3693;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_1829;
wire n_1338;
wire n_1327;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_2565;
wire n_4201;
wire n_1636;
wire n_1687;
wire n_4584;
wire n_3184;
wire n_4155;
wire n_3890;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1680;
wire n_1195;
wire n_4304;
wire n_4821;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_3641;
wire n_4887;
wire n_3996;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_1841;
wire n_2685;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_3722;
wire n_3802;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_4806;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_1007;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_3765;
wire n_2216;
wire n_4259;
wire n_1620;
wire n_3518;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_2899;
wire n_3351;
wire n_2008;
wire n_2859;
wire n_2564;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_1764;
wire n_1019;
wire n_1250;
wire n_1190;
wire n_4598;
wire n_3259;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_2114;
wire n_1609;
wire n_3530;
wire n_1132;
wire n_4548;
wire n_1803;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_2660;
wire n_4604;
wire n_3467;
wire n_4240;
wire n_2219;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_2539;
wire n_1701;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4126;
wire n_4103;
wire n_4710;
wire n_3282;
wire n_1003;
wire n_2708;
wire n_2748;
wire n_2224;
wire n_2233;
wire n_2499;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_1553;
wire n_3542;
wire n_1090;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_3171;
wire n_1733;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_1189;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_4205;
wire n_3790;
wire n_2404;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_4504;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_2852;
wire n_2132;
wire n_1236;
wire n_3412;
wire n_1712;
wire n_4537;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_4184;
wire n_2468;
wire n_3248;
wire n_2606;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_4876;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_4747;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_2481;
wire n_4409;
wire n_1264;
wire n_2808;
wire n_3396;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_2977;
wire n_1682;
wire n_3599;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_4152;
wire n_1352;
wire n_2328;
wire n_4587;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_4500;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_2419;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_951;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_4496;
wire n_1528;
wire n_3840;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_1413;
wire n_2464;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_2414;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_3284;
wire n_2875;
wire n_1437;
wire n_2747;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_4316;
wire n_3328;
wire n_2763;
wire n_994;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_4306;
wire n_2997;
wire n_3735;
wire n_961;
wire n_2127;
wire n_3028;
wire n_3228;
wire n_3706;
wire n_1432;
wire n_3322;
wire n_996;
wire n_1174;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_2694;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_3960;
wire n_4007;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_982;
wire n_2180;
wire n_3376;
wire n_2617;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_2086;
wire n_4832;
wire n_3666;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2108;
wire n_2535;
wire n_2945;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_3773;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_1124;
wire n_2688;
wire n_3302;
wire n_1673;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_4340;
wire n_1476;
wire n_935;
wire n_1054;
wire n_2027;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_1642;
wire n_2447;
wire n_3358;
wire n_2894;
wire n_2587;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_3410;
wire n_975;
wire n_4900;
wire n_934;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_2299;
wire n_2078;
wire n_3709;
wire n_3011;
wire n_2315;
wire n_3623;
wire n_2157;
wire n_3446;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_4334;
wire n_2211;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_1501;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_2893;
wire n_2009;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_1005;
wire n_4581;
wire n_4618;
wire n_1105;
wire n_2898;
wire n_2519;
wire n_2231;
wire n_1000;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_4670;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_1939;
wire n_4053;
wire n_4279;
wire n_3937;
wire n_3303;
wire n_4555;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_1693;
wire n_2081;
wire n_2993;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_3989;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_4415;
wire n_3343;
wire n_3163;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_967;
wire n_4263;
wire n_3725;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_1336;
wire n_1358;
wire n_3318;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_3430;
wire n_1685;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_1074;
wire n_1462;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_1398;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_1692;
wire n_4796;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_3837;
wire n_4841;
wire n_3076;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2855;
wire n_2653;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_2331;
wire n_1600;
wire n_4701;
wire n_4088;
wire n_2136;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_1822;
wire n_1804;
wire n_1581;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_2262;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_4327;
wire n_2656;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_1016;
wire n_4465;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_983;
wire n_4224;
wire n_4868;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_4387;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_992;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_1080;
wire n_2290;
wire n_957;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_4668;
wire n_2383;
wire n_2640;
wire n_1492;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_2230;
wire n_3033;
wire n_2151;
wire n_4912;
wire n_1971;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_2571;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_989;
wire n_1668;
wire n_1681;
wire n_4031;
wire n_939;
wire n_4120;
wire n_3896;
wire n_3533;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_4311;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_1606;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_4650;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_979;
wire n_1999;
wire n_3810;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_2826;
wire n_2112;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_4671;
wire n_1326;
wire n_978;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_3618;
wire n_2727;
wire n_2719;
wire n_2213;
wire n_3521;
wire n_2723;
wire n_4054;
wire n_1569;
wire n_4012;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_2292;
wire n_3560;
wire n_1742;
wire n_1818;
wire n_3847;
wire n_2203;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_2646;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_4755;
wire n_3827;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_4136;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1360;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_1036;
wire n_1106;
wire n_4655;
wire n_1634;
wire n_1452;
wire n_4953;
wire n_4570;
wire n_3966;
wire n_4293;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_2819;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_3436;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_4527;
wire n_2877;
wire n_1996;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_4407;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_3680;
wire n_3624;
wire n_2467;
wire n_4292;
wire n_3145;
wire n_2662;
wire n_3872;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_1566;
wire n_1464;
wire n_944;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_4929;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_1009;
wire n_2160;
wire n_2991;
wire n_2699;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_4427;
wire n_3505;
wire n_4564;
wire n_2934;
wire n_942;
wire n_4042;
wire n_2525;
wire n_4624;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_4958;
wire n_4297;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_2095;
wire n_2486;
wire n_2521;
wire n_1574;
wire n_4764;
wire n_4899;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_2986;
wire n_2400;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_1357;
wire n_4566;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_2117;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_3638;
wire n_2106;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_964;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_4133;
wire n_3985;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_2745;
wire n_2110;
wire n_3747;
wire n_991;
wire n_1323;
wire n_3710;
wire n_1429;
wire n_3209;
wire n_2026;
wire n_3588;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_2105;
wire n_2187;
wire n_2642;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_4048;
wire n_4084;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_2849;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_4860;
wire n_4438;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_3047;
wire n_2610;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_4149;
wire n_3930;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_4383;
wire n_2709;
wire n_2244;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_2665;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_993;
wire n_2581;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_1406;
wire n_3591;
wire n_2137;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_3139;
wire n_4715;
wire n_4222;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_1167;
wire n_3231;
wire n_3138;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_3454;
wire n_4143;
wire n_4410;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_1513;
wire n_1788;
wire n_2348;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_2248;
wire n_958;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_3846;
wire n_4328;
wire n_1433;
wire n_1907;
wire n_3994;
wire n_2135;
wire n_1088;
wire n_1102;
wire n_4487;
wire n_1165;
wire n_4148;
wire n_3066;
wire n_2869;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_2667;
wire n_1565;
wire n_2325;
wire n_3346;
wire n_3391;
wire n_1542;
wire n_1547;
wire n_1362;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_3045;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_2021;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_2061;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_3042;
wire n_2561;
wire n_2491;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_4811;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_1759;
wire n_2096;
wire n_2296;
wire n_1911;
wire n_2870;
wire n_4869;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_1419;
wire n_4738;
wire n_980;
wire n_1193;
wire n_2928;
wire n_3557;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_4086;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_999;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_1499;
wire n_2155;
wire n_966;
wire n_3938;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_3053;
wire n_1039;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_1762;
wire n_940;
wire n_4944;
wire n_4468;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_1791;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_1164;
wire n_3749;
wire n_4452;
wire n_3691;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_4280;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_1665;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_1417;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_1410;
wire n_988;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_4662;
wire n_2658;

BUFx10_ASAP7_75t_L g933 ( 
.A(n_196),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_789),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_713),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_855),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_644),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_901),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_925),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_628),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_292),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_785),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_414),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_923),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_374),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_18),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_575),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_173),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_49),
.Y(n_949)
);

BUFx10_ASAP7_75t_L g950 ( 
.A(n_761),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_130),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_748),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_71),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_497),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_87),
.Y(n_955)
);

BUFx10_ASAP7_75t_L g956 ( 
.A(n_858),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_334),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_315),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_810),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_456),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_764),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_369),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_206),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_894),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_875),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_679),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_797),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_846),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_226),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_227),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_612),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_694),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_595),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_796),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_150),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_638),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_848),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_892),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_880),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_296),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_772),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_845),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_849),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_703),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_852),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_177),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_334),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_526),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_632),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_54),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_329),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_60),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_694),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_118),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_864),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_902),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_586),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_263),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_612),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_463),
.Y(n_1000)
);

BUFx5_ASAP7_75t_L g1001 ( 
.A(n_159),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_293),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_736),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_792),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_803),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_300),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_236),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_230),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_353),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_204),
.Y(n_1010)
);

BUFx5_ASAP7_75t_L g1011 ( 
.A(n_793),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_678),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_251),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_527),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_112),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_660),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_78),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_317),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_73),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_145),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_481),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_447),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_876),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_806),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_621),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_781),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_90),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_881),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_323),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_379),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_539),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_503),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_492),
.Y(n_1033)
);

BUFx10_ASAP7_75t_L g1034 ( 
.A(n_796),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_815),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_788),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_928),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_403),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_336),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_738),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_930),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_891),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_307),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_738),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_229),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_779),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_8),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_470),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_905),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_927),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_255),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_644),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_413),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_230),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_113),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_617),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_790),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_287),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_404),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_731),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_359),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_675),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_887),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_120),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_16),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_861),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_697),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_275),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_813),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_193),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_8),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_306),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_885),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_435),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_795),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_312),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_39),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_915),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_567),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_141),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_28),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_256),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_578),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_572),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_493),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_456),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_842),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_357),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_767),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_193),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_706),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_909),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_837),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_85),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_775),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_326),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_439),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_812),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_148),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_921),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_926),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_609),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_549),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_396),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_879),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_829),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_737),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_877),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_55),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_930),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_442),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_596),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_125),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_890),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_444),
.Y(n_1115)
);

BUFx10_ASAP7_75t_L g1116 ( 
.A(n_523),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_730),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_452),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_883),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_833),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_819),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_707),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_384),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_807),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_816),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_545),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_356),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_397),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_684),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_833),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_854),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_886),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_212),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_633),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_825),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_734),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_504),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_680),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_629),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_375),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_508),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_432),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_917),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_439),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_703),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_196),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_523),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_303),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_561),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_859),
.Y(n_1150)
);

BUFx8_ASAP7_75t_SL g1151 ( 
.A(n_875),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_717),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_515),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_868),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_231),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_924),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_358),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_518),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_102),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_869),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_382),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_530),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_363),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_200),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_831),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_282),
.Y(n_1166)
);

BUFx10_ASAP7_75t_L g1167 ( 
.A(n_910),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_322),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_229),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_705),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_777),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_4),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_217),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_371),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_350),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_280),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_699),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_335),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_837),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_789),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_927),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_736),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_293),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_402),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_720),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_13),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_799),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_294),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_846),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_659),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_514),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_883),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_325),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_44),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_919),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_774),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_755),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_741),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_382),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_233),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_50),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_473),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_53),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_438),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_709),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_199),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_161),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_811),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_839),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_494),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_65),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_29),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_596),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_605),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_863),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_12),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_917),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_59),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_754),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_408),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_567),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_178),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_253),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_821),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_97),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_646),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_866),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_824),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_853),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_914),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_5),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_904),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_258),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_186),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_34),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_371),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_907),
.Y(n_1237)
);

CKINVDCx14_ASAP7_75t_R g1238 ( 
.A(n_433),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_880),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_803),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_811),
.Y(n_1241)
);

INVxp33_ASAP7_75t_L g1242 ( 
.A(n_152),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_275),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_639),
.Y(n_1244)
);

INVxp67_ASAP7_75t_L g1245 ( 
.A(n_716),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_541),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_834),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_214),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_801),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_793),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_316),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_623),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_597),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_841),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_3),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_518),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_162),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_58),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_685),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_14),
.Y(n_1260)
);

BUFx10_ASAP7_75t_L g1261 ( 
.A(n_155),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_818),
.Y(n_1262)
);

CKINVDCx14_ASAP7_75t_R g1263 ( 
.A(n_830),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_350),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_859),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_102),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_532),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_0),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_827),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_143),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_908),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_446),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_477),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_553),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_380),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_895),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_160),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_72),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_157),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_504),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_812),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_828),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_298),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_860),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_244),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_780),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_870),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_873),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_314),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_158),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_835),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_483),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_447),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_882),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_838),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_168),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_47),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_556),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_897),
.Y(n_1299)
);

BUFx5_ASAP7_75t_L g1300 ( 
.A(n_862),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_733),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_90),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_10),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_663),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_896),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_663),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_798),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_309),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_802),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_298),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_808),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_804),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_367),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_475),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_722),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_794),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_840),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_920),
.Y(n_1318)
);

BUFx5_ASAP7_75t_L g1319 ( 
.A(n_627),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_916),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_547),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_570),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_297),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_305),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_884),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_129),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_872),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_820),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_861),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_410),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_647),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_222),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_342),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_781),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_352),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_617),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_135),
.Y(n_1337)
);

BUFx5_ASAP7_75t_L g1338 ( 
.A(n_670),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_899),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_274),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_351),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_911),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_860),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_69),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_851),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_109),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_465),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_543),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_419),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_304),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_889),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_814),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_15),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_0),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_902),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_306),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_763),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_795),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_374),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_315),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_577),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_669),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_621),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_922),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_684),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_384),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_513),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_822),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_761),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_344),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_87),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_533),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_542),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_820),
.Y(n_1374)
);

BUFx10_ASAP7_75t_L g1375 ( 
.A(n_692),
.Y(n_1375)
);

BUFx10_ASAP7_75t_L g1376 ( 
.A(n_73),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_826),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_484),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_135),
.Y(n_1379)
);

BUFx10_ASAP7_75t_L g1380 ( 
.A(n_13),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_353),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_867),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_410),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_931),
.Y(n_1384)
);

BUFx5_ASAP7_75t_L g1385 ( 
.A(n_403),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_759),
.Y(n_1386)
);

BUFx10_ASAP7_75t_L g1387 ( 
.A(n_241),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_666),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_839),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_620),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_857),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_202),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_805),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_429),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_705),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_900),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_0),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_779),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_844),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_891),
.Y(n_1400)
);

CKINVDCx16_ASAP7_75t_R g1401 ( 
.A(n_11),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_439),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_554),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_922),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_113),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_727),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_559),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_878),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_878),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_142),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_429),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_320),
.Y(n_1412)
);

CKINVDCx14_ASAP7_75t_R g1413 ( 
.A(n_412),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_850),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_858),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_838),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_847),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_198),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_413),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_906),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_836),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_913),
.Y(n_1422)
);

BUFx10_ASAP7_75t_L g1423 ( 
.A(n_342),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_871),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_11),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_910),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_932),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_633),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_117),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_315),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_19),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_865),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_398),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_929),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_770),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_671),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_618),
.Y(n_1437)
);

BUFx2_ASAP7_75t_SL g1438 ( 
.A(n_832),
.Y(n_1438)
);

BUFx10_ASAP7_75t_L g1439 ( 
.A(n_848),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_843),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_226),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_866),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_202),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_882),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_732),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_809),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_620),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_483),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_741),
.Y(n_1449)
);

BUFx10_ASAP7_75t_L g1450 ( 
.A(n_167),
.Y(n_1450)
);

BUFx10_ASAP7_75t_L g1451 ( 
.A(n_120),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_797),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_48),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_399),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_823),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_575),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_815),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_273),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_670),
.Y(n_1459)
);

BUFx8_ASAP7_75t_SL g1460 ( 
.A(n_27),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_123),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_157),
.Y(n_1462)
);

CKINVDCx16_ASAP7_75t_R g1463 ( 
.A(n_788),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_773),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_604),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_296),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_664),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_619),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_783),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_447),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_559),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_489),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_768),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_438),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_888),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_67),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_823),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_725),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_893),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_856),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_219),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_918),
.Y(n_1482)
);

BUFx8_ASAP7_75t_SL g1483 ( 
.A(n_484),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_742),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_561),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_258),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_822),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_800),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_480),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_807),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_594),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_3),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_746),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_134),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_269),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_280),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_250),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_449),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_449),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_544),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_182),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_885),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_893),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_903),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_370),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_648),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_619),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_137),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_740),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_271),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_817),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_403),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_6),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_856),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_237),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_293),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_336),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_97),
.Y(n_1518)
);

BUFx8_ASAP7_75t_SL g1519 ( 
.A(n_632),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_347),
.Y(n_1520)
);

CKINVDCx16_ASAP7_75t_R g1521 ( 
.A(n_912),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_898),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_58),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_874),
.Y(n_1524)
);

CKINVDCx16_ASAP7_75t_R g1525 ( 
.A(n_1401),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1011),
.Y(n_1526)
);

INVxp67_ASAP7_75t_SL g1527 ( 
.A(n_1045),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1004),
.B(n_1),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_989),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_989),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1238),
.Y(n_1531)
);

INVxp33_ASAP7_75t_L g1532 ( 
.A(n_1086),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1224),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1332),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1224),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1011),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1021),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1077),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1238),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1413),
.Y(n_1540)
);

BUFx2_ASAP7_75t_SL g1541 ( 
.A(n_957),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1003),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1413),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1006),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1115),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1460),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1162),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1045),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1483),
.Y(n_1549)
);

CKINVDCx16_ASAP7_75t_R g1550 ( 
.A(n_1336),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_987),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1002),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1003),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1242),
.B(n_1),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1188),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1022),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1500),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1053),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_943),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1263),
.Y(n_1560)
);

CKINVDCx16_ASAP7_75t_R g1561 ( 
.A(n_1463),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1095),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_945),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1263),
.Y(n_1564)
);

INVxp67_ASAP7_75t_SL g1565 ( 
.A(n_957),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_947),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_970),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1151),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1519),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_973),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1079),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1113),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_975),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_986),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_1199),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1009),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1018),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1233),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1019),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1020),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_1246),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1030),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1054),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_941),
.Y(n_1584)
);

INVxp67_ASAP7_75t_SL g1585 ( 
.A(n_1038),
.Y(n_1585)
);

BUFx2_ASAP7_75t_SL g1586 ( 
.A(n_1038),
.Y(n_1586)
);

CKINVDCx16_ASAP7_75t_R g1587 ( 
.A(n_1521),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1316),
.B(n_1067),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1374),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1083),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1064),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1477),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_1289),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1065),
.Y(n_1594)
);

CKINVDCx20_ASAP7_75t_R g1595 ( 
.A(n_1360),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1072),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_1379),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_1083),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1084),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1472),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_946),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1111),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1128),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1489),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_948),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1137),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_949),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_951),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1142),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_1497),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_942),
.B(n_2),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1510),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1157),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1178),
.Y(n_1614)
);

INVxp67_ASAP7_75t_SL g1615 ( 
.A(n_1088),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_959),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_953),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_954),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_955),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1186),
.Y(n_1620)
);

INVxp33_ASAP7_75t_L g1621 ( 
.A(n_944),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1191),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1200),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1207),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1210),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1211),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1218),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1220),
.Y(n_1628)
);

INVxp67_ASAP7_75t_SL g1629 ( 
.A(n_1088),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_971),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1222),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1323),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_958),
.Y(n_1633)
);

CKINVDCx20_ASAP7_75t_R g1634 ( 
.A(n_995),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_960),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_962),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1052),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_963),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1223),
.Y(n_1639)
);

NOR2xp67_ASAP7_75t_L g1640 ( 
.A(n_981),
.B(n_2),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1056),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_969),
.Y(n_1642)
);

INVxp33_ASAP7_75t_L g1643 ( 
.A(n_964),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1231),
.Y(n_1644)
);

CKINVDCx16_ASAP7_75t_R g1645 ( 
.A(n_933),
.Y(n_1645)
);

CKINVDCx20_ASAP7_75t_R g1646 ( 
.A(n_1073),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1323),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1235),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1089),
.Y(n_1649)
);

CKINVDCx20_ASAP7_75t_R g1650 ( 
.A(n_1132),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1236),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_988),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_990),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1253),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1255),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1565),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1565),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1585),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1544),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1534),
.B(n_1075),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1585),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1598),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1598),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1541),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1586),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1590),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1608),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1532),
.B(n_933),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1590),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1534),
.B(n_1116),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1632),
.Y(n_1671)
);

INVxp33_ASAP7_75t_SL g1672 ( 
.A(n_1531),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1632),
.B(n_991),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1542),
.Y(n_1674)
);

XOR2xp5_ASAP7_75t_L g1675 ( 
.A(n_1551),
.B(n_1136),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1584),
.Y(n_1676)
);

INVx4_ASAP7_75t_L g1677 ( 
.A(n_1645),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1601),
.Y(n_1678)
);

OA21x2_ASAP7_75t_L g1679 ( 
.A1(n_1526),
.A2(n_1061),
.B(n_1039),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1527),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1539),
.B(n_1001),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1544),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1615),
.B(n_1629),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1647),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1544),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1544),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1553),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1537),
.B(n_1245),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1538),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1605),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1562),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1536),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1545),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1548),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1529),
.Y(n_1695)
);

NAND3xp33_ASAP7_75t_L g1696 ( 
.A(n_1555),
.B(n_994),
.C(n_992),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1547),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1530),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1618),
.B(n_997),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1607),
.Y(n_1700)
);

NAND2x1_ASAP7_75t_L g1701 ( 
.A(n_1554),
.B(n_1039),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1533),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1535),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1559),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1560),
.B(n_1452),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1636),
.B(n_998),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1617),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1563),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1638),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1566),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1567),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1570),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1573),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1574),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1576),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1577),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1579),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1580),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1582),
.Y(n_1719)
);

AND2x6_ASAP7_75t_L g1720 ( 
.A(n_1557),
.B(n_1330),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1540),
.B(n_1001),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1589),
.B(n_1116),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1583),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1652),
.B(n_1154),
.Y(n_1724)
);

OA21x2_ASAP7_75t_L g1725 ( 
.A1(n_1591),
.A2(n_1164),
.B(n_1061),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1594),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1596),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1543),
.B(n_1000),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1599),
.Y(n_1729)
);

AND2x6_ASAP7_75t_L g1730 ( 
.A(n_1528),
.B(n_1330),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1602),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1603),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1619),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1606),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1609),
.B(n_1613),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1614),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1620),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1622),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1623),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1525),
.A2(n_1008),
.B1(n_1013),
.B2(n_1010),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1633),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_L g1742 ( 
.A(n_1624),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1625),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1626),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1627),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1628),
.Y(n_1746)
);

INVx3_ASAP7_75t_L g1747 ( 
.A(n_1631),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1639),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1644),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1648),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1651),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1654),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1655),
.Y(n_1753)
);

AND2x6_ASAP7_75t_L g1754 ( 
.A(n_1611),
.B(n_1381),
.Y(n_1754)
);

NAND2xp33_ASAP7_75t_L g1755 ( 
.A(n_1564),
.B(n_1001),
.Y(n_1755)
);

AND2x6_ASAP7_75t_L g1756 ( 
.A(n_1588),
.B(n_1381),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1640),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1592),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1635),
.B(n_1185),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1621),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1642),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1653),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1643),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1550),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1561),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1587),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1546),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1549),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1568),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1569),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1552),
.Y(n_1771)
);

INVx4_ASAP7_75t_L g1772 ( 
.A(n_1556),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1558),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1571),
.Y(n_1774)
);

BUFx8_ASAP7_75t_L g1775 ( 
.A(n_1572),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1575),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1578),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1581),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1593),
.B(n_1261),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1595),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1597),
.B(n_1261),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1600),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1604),
.B(n_1295),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1610),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1612),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1616),
.B(n_1427),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1630),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1634),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1637),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1641),
.A2(n_1196),
.B1(n_1239),
.B2(n_1180),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1646),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1649),
.B(n_1014),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1650),
.Y(n_1793)
);

BUFx8_ASAP7_75t_L g1794 ( 
.A(n_1555),
.Y(n_1794)
);

OA21x2_ASAP7_75t_L g1795 ( 
.A1(n_1526),
.A2(n_1176),
.B(n_1164),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1532),
.B(n_1376),
.Y(n_1796)
);

BUFx6f_ASAP7_75t_L g1797 ( 
.A(n_1544),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1542),
.Y(n_1798)
);

NAND2x1_ASAP7_75t_L g1799 ( 
.A(n_1554),
.B(n_1176),
.Y(n_1799)
);

INVx4_ASAP7_75t_L g1800 ( 
.A(n_1645),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1565),
.Y(n_1801)
);

OA21x2_ASAP7_75t_L g1802 ( 
.A1(n_1526),
.A2(n_1278),
.B(n_1202),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1565),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1544),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1542),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1565),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1542),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1532),
.B(n_1376),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1542),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1542),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1532),
.B(n_1380),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1565),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1542),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1532),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1565),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1590),
.B(n_1015),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1565),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1525),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1542),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1565),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1544),
.Y(n_1821)
);

OR2x6_ASAP7_75t_L g1822 ( 
.A(n_1534),
.B(n_1438),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1542),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1645),
.B(n_1001),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1590),
.B(n_1017),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1542),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1534),
.B(n_1095),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1534),
.B(n_1357),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1542),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1565),
.Y(n_1830)
);

INVx1_ASAP7_75t_SL g1831 ( 
.A(n_1532),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1565),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1532),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1544),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_L g1835 ( 
.A(n_1544),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1565),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1565),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1544),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1565),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1565),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1542),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1608),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1565),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1565),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1590),
.B(n_1029),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1565),
.Y(n_1846)
);

CKINVDCx20_ASAP7_75t_R g1847 ( 
.A(n_1551),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1534),
.B(n_1357),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1544),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1532),
.B(n_1380),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1565),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1590),
.B(n_1031),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1534),
.B(n_1404),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1565),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1532),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1565),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1565),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1565),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1565),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1542),
.Y(n_1860)
);

AND3x2_ASAP7_75t_L g1861 ( 
.A(n_1534),
.B(n_1278),
.C(n_1202),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1542),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1542),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1542),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1534),
.B(n_1404),
.Y(n_1865)
);

AND2x2_ASAP7_75t_R g1866 ( 
.A(n_1551),
.B(n_1240),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1534),
.B(n_1457),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1565),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1544),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1726),
.Y(n_1870)
);

BUFx2_ASAP7_75t_L g1871 ( 
.A(n_1831),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1745),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1747),
.Y(n_1873)
);

AND2x6_ASAP7_75t_L g1874 ( 
.A(n_1670),
.B(n_1392),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1763),
.B(n_1001),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1680),
.B(n_1032),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1728),
.B(n_1033),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1749),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1855),
.B(n_1353),
.Y(n_1879)
);

AND2x2_ASAP7_75t_SL g1880 ( 
.A(n_1677),
.B(n_1353),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1814),
.A2(n_1047),
.B1(n_1048),
.B2(n_1043),
.Y(n_1881)
);

INVx3_ASAP7_75t_L g1882 ( 
.A(n_1800),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1656),
.A2(n_1443),
.B1(n_1470),
.B2(n_1392),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1657),
.A2(n_1470),
.B1(n_1443),
.B2(n_1283),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_SL g1885 ( 
.A(n_1833),
.B(n_1051),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1673),
.B(n_1001),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1689),
.Y(n_1887)
);

NAND2xp33_ASAP7_75t_L g1888 ( 
.A(n_1720),
.B(n_1385),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1760),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1658),
.A2(n_1290),
.B1(n_1296),
.B2(n_1257),
.Y(n_1890)
);

OAI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1707),
.A2(n_1058),
.B1(n_1059),
.B2(n_1055),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1660),
.B(n_1068),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1725),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1670),
.A2(n_1071),
.B1(n_1074),
.B2(n_1070),
.Y(n_1894)
);

AND2x6_ASAP7_75t_L g1895 ( 
.A(n_1661),
.B(n_1359),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1691),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1693),
.Y(n_1897)
);

INVx4_ASAP7_75t_L g1898 ( 
.A(n_1720),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1679),
.Y(n_1899)
);

NAND2x1p5_ASAP7_75t_L g1900 ( 
.A(n_1668),
.B(n_980),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1668),
.A2(n_1080),
.B1(n_1082),
.B2(n_1076),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1691),
.Y(n_1902)
);

INVx3_ASAP7_75t_L g1903 ( 
.A(n_1694),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1795),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1808),
.B(n_1241),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1816),
.B(n_1385),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1684),
.B(n_1666),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1808),
.B(n_1811),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1697),
.Y(n_1909)
);

INVx6_ASAP7_75t_L g1910 ( 
.A(n_1761),
.Y(n_1910)
);

BUFx3_ASAP7_75t_L g1911 ( 
.A(n_1676),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1694),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1825),
.B(n_1385),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1845),
.B(n_1385),
.Y(n_1914)
);

CKINVDCx6p67_ASAP7_75t_R g1915 ( 
.A(n_1822),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1811),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1850),
.A2(n_1090),
.B1(n_1094),
.B2(n_1085),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1852),
.B(n_1385),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1802),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1829),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1662),
.A2(n_1801),
.B1(n_1803),
.B2(n_1663),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1702),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1702),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1695),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1805),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1708),
.Y(n_1926)
);

OAI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1758),
.A2(n_1097),
.B1(n_1099),
.B2(n_1096),
.Y(n_1927)
);

INVx5_ASAP7_75t_L g1928 ( 
.A(n_1720),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1806),
.A2(n_1104),
.B1(n_1109),
.B2(n_1103),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1669),
.B(n_1112),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1698),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1812),
.Y(n_1932)
);

INVx3_ASAP7_75t_L g1933 ( 
.A(n_1841),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1710),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1710),
.Y(n_1935)
);

INVxp67_ASAP7_75t_SL g1936 ( 
.A(n_1796),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1664),
.B(n_1118),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1815),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1817),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_L g1940 ( 
.A(n_1696),
.B(n_1126),
.C(n_1123),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1665),
.B(n_1127),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1667),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1713),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1820),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1830),
.A2(n_1308),
.B1(n_1313),
.B2(n_1297),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1832),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1678),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1774),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1683),
.B(n_1385),
.Y(n_1949)
);

AO22x1_ASAP7_75t_L g1950 ( 
.A1(n_1794),
.A2(n_1147),
.B1(n_1148),
.B2(n_1133),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1775),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1722),
.B(n_1149),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1827),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1671),
.B(n_1155),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1709),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1836),
.B(n_1161),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1837),
.Y(n_1957)
);

OAI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1822),
.A2(n_1166),
.B1(n_1168),
.B2(n_1163),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1839),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1840),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1699),
.B(n_1169),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1713),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1717),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1843),
.A2(n_1321),
.B1(n_1324),
.B2(n_1314),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1717),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1842),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1729),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1844),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1762),
.B(n_1172),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1729),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1846),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1731),
.Y(n_1972)
);

NAND3xp33_ASAP7_75t_L g1973 ( 
.A(n_1706),
.B(n_1174),
.C(n_1173),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1851),
.Y(n_1974)
);

INVxp67_ASAP7_75t_SL g1975 ( 
.A(n_1735),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1731),
.Y(n_1976)
);

NAND2xp33_ASAP7_75t_L g1977 ( 
.A(n_1754),
.B(n_1011),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1742),
.Y(n_1978)
);

OR2x6_ASAP7_75t_L g1979 ( 
.A(n_1772),
.B(n_1012),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1847),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1742),
.B(n_1175),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1854),
.Y(n_1982)
);

INVx5_ASAP7_75t_L g1983 ( 
.A(n_1860),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1690),
.Y(n_1984)
);

AND2x6_ASAP7_75t_L g1985 ( 
.A(n_1856),
.B(n_1006),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1857),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1761),
.Y(n_1987)
);

OR2x6_ASAP7_75t_L g1988 ( 
.A(n_1700),
.B(n_1012),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1701),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1799),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1674),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1687),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1724),
.B(n_1183),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1765),
.B(n_1244),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1792),
.B(n_1027),
.Y(n_1995)
);

XOR2x2_ASAP7_75t_L g1996 ( 
.A(n_1675),
.B(n_1773),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1858),
.B(n_1184),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1733),
.B(n_1387),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1766),
.B(n_1252),
.Y(n_1999)
);

INVx6_ASAP7_75t_L g2000 ( 
.A(n_1828),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1741),
.B(n_1387),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1859),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1868),
.B(n_1193),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1798),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1703),
.Y(n_2005)
);

AO21x2_ASAP7_75t_L g2006 ( 
.A1(n_1681),
.A2(n_1333),
.B(n_1326),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1715),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1704),
.B(n_1194),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1807),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1711),
.B(n_1201),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1824),
.B(n_1203),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1757),
.B(n_1712),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1718),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1779),
.B(n_1081),
.Y(n_2014)
);

NAND2xp33_ASAP7_75t_L g2015 ( 
.A(n_1754),
.B(n_1011),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1719),
.Y(n_2016)
);

OAI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1740),
.A2(n_1212),
.B1(n_1213),
.B2(n_1206),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1848),
.B(n_1423),
.Y(n_2018)
);

AND2x6_ASAP7_75t_L g2019 ( 
.A(n_1767),
.B(n_1006),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_1809),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1810),
.Y(n_2021)
);

INVx5_ASAP7_75t_L g2022 ( 
.A(n_1756),
.Y(n_2022)
);

AO22x2_ASAP7_75t_L g2023 ( 
.A1(n_1866),
.A2(n_1140),
.B1(n_1144),
.B2(n_1141),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1764),
.B(n_1276),
.Y(n_2024)
);

AND2x6_ASAP7_75t_L g2025 ( 
.A(n_1768),
.B(n_1006),
.Y(n_2025)
);

OAI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1714),
.A2(n_1513),
.B1(n_1515),
.B2(n_1512),
.Y(n_2026)
);

OR2x6_ASAP7_75t_L g2027 ( 
.A(n_1781),
.B(n_1063),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1723),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1727),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1752),
.Y(n_2030)
);

BUFx10_ASAP7_75t_L g2031 ( 
.A(n_1818),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1716),
.B(n_1523),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1732),
.B(n_1516),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1813),
.Y(n_2034)
);

INVx1_ASAP7_75t_SL g2035 ( 
.A(n_1853),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_1819),
.Y(n_2036)
);

BUFx2_ASAP7_75t_L g2037 ( 
.A(n_1756),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1823),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1770),
.B(n_1320),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_1759),
.B(n_1216),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1734),
.B(n_1518),
.Y(n_2041)
);

INVx5_ASAP7_75t_L g2042 ( 
.A(n_1756),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1736),
.B(n_1221),
.Y(n_2043)
);

BUFx10_ASAP7_75t_L g2044 ( 
.A(n_1783),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1737),
.B(n_1225),
.Y(n_2045)
);

INVx5_ASAP7_75t_L g2046 ( 
.A(n_1730),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1738),
.B(n_1234),
.Y(n_2047)
);

OAI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_1692),
.A2(n_1340),
.B(n_1335),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_1865),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1739),
.B(n_1243),
.Y(n_2050)
);

INVx3_ASAP7_75t_L g2051 ( 
.A(n_1826),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1743),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1744),
.B(n_1501),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1746),
.B(n_1508),
.Y(n_2054)
);

INVx6_ASAP7_75t_L g2055 ( 
.A(n_1867),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_SL g2056 ( 
.A(n_1672),
.B(n_1248),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1748),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1730),
.A2(n_1346),
.B1(n_1347),
.B2(n_1344),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1705),
.B(n_1251),
.Y(n_2059)
);

AOI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_1730),
.A2(n_1754),
.B1(n_1750),
.B2(n_1753),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1751),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1862),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1863),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1864),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1688),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1861),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1721),
.B(n_1755),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1786),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1769),
.A2(n_1349),
.B1(n_1366),
.B2(n_1348),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1659),
.Y(n_2070)
);

INVx2_ASAP7_75t_SL g2071 ( 
.A(n_1785),
.Y(n_2071)
);

AOI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_1776),
.A2(n_1258),
.B1(n_1260),
.B2(n_1256),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1785),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1771),
.B(n_1264),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_1787),
.B(n_1266),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1659),
.Y(n_2076)
);

BUFx4f_ASAP7_75t_L g2077 ( 
.A(n_1788),
.Y(n_2077)
);

INVx4_ASAP7_75t_L g2078 ( 
.A(n_1788),
.Y(n_2078)
);

OAI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_1777),
.A2(n_1268),
.B1(n_1270),
.B2(n_1267),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1789),
.B(n_1791),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1682),
.Y(n_2081)
);

BUFx3_ASAP7_75t_L g2082 ( 
.A(n_1789),
.Y(n_2082)
);

BUFx10_ASAP7_75t_L g2083 ( 
.A(n_1778),
.Y(n_2083)
);

BUFx2_ASAP7_75t_L g2084 ( 
.A(n_1780),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1782),
.B(n_1423),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1682),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1685),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1686),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1686),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_1793),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1784),
.B(n_1272),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1797),
.B(n_1273),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1797),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_1804),
.A2(n_1373),
.B1(n_1383),
.B2(n_1370),
.Y(n_2094)
);

INVx4_ASAP7_75t_L g2095 ( 
.A(n_1804),
.Y(n_2095)
);

NAND2xp33_ASAP7_75t_L g2096 ( 
.A(n_1821),
.B(n_1011),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1821),
.B(n_1274),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1834),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1834),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1835),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1835),
.B(n_1275),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1838),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_1790),
.B(n_1277),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1838),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1849),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1849),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1869),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_1869),
.B(n_1279),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_1831),
.B(n_1450),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1725),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_1656),
.A2(n_1402),
.B1(n_1403),
.B2(n_1394),
.Y(n_2111)
);

INVxp67_ASAP7_75t_SL g2112 ( 
.A(n_1814),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1725),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1726),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_L g2115 ( 
.A(n_1691),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_1831),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_1831),
.B(n_1411),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1763),
.B(n_1280),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1726),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1725),
.Y(n_2120)
);

BUFx3_ASAP7_75t_L g2121 ( 
.A(n_1831),
.Y(n_2121)
);

INVx2_ASAP7_75t_SL g2122 ( 
.A(n_1831),
.Y(n_2122)
);

AO22x2_ASAP7_75t_L g2123 ( 
.A1(n_1675),
.A2(n_1430),
.B1(n_1150),
.B2(n_1247),
.Y(n_2123)
);

XNOR2xp5_ASAP7_75t_L g2124 ( 
.A(n_1675),
.B(n_1522),
.Y(n_2124)
);

INVx3_ASAP7_75t_L g2125 ( 
.A(n_1831),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_1680),
.B(n_1292),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1725),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1726),
.Y(n_2128)
);

INVxp67_ASAP7_75t_SL g2129 ( 
.A(n_1814),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1831),
.B(n_1450),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1726),
.Y(n_2131)
);

OR2x6_ASAP7_75t_L g2132 ( 
.A(n_1677),
.B(n_1063),
.Y(n_2132)
);

INVxp67_ASAP7_75t_SL g2133 ( 
.A(n_1814),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1726),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1725),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1831),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_1680),
.B(n_1293),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1726),
.Y(n_2138)
);

BUFx3_ASAP7_75t_L g2139 ( 
.A(n_1831),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1725),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1726),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1763),
.B(n_1298),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1831),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_1763),
.B(n_1302),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1763),
.B(n_1303),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1725),
.Y(n_2146)
);

NAND2xp33_ASAP7_75t_L g2147 ( 
.A(n_1720),
.B(n_1011),
.Y(n_2147)
);

BUFx4f_ASAP7_75t_L g2148 ( 
.A(n_1761),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1726),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_1831),
.B(n_1310),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1726),
.Y(n_2151)
);

INVx1_ASAP7_75t_SL g2152 ( 
.A(n_1831),
.Y(n_2152)
);

INVxp67_ASAP7_75t_R g2153 ( 
.A(n_1814),
.Y(n_2153)
);

NAND2xp33_ASAP7_75t_L g2154 ( 
.A(n_1720),
.B(n_1300),
.Y(n_2154)
);

BUFx6f_ASAP7_75t_L g2155 ( 
.A(n_1691),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1726),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_1831),
.B(n_1451),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1726),
.Y(n_2158)
);

INVx3_ASAP7_75t_L g2159 ( 
.A(n_1831),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_SL g2160 ( 
.A(n_1763),
.B(n_1322),
.Y(n_2160)
);

CKINVDCx20_ASAP7_75t_R g2161 ( 
.A(n_1831),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1831),
.B(n_1451),
.Y(n_2162)
);

AND2x2_ASAP7_75t_SL g2163 ( 
.A(n_1871),
.B(n_1885),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1975),
.Y(n_2164)
);

OR2x6_ASAP7_75t_L g2165 ( 
.A(n_2121),
.B(n_1102),
.Y(n_2165)
);

INVxp67_ASAP7_75t_L g2166 ( 
.A(n_1871),
.Y(n_2166)
);

BUFx5_ASAP7_75t_L g2167 ( 
.A(n_1985),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1893),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1932),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_2152),
.B(n_1337),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1874),
.B(n_1341),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2110),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1938),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1874),
.B(n_1350),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1874),
.B(n_1354),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_2116),
.B(n_1367),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1939),
.Y(n_2177)
);

OR2x6_ASAP7_75t_L g2178 ( 
.A(n_2139),
.B(n_1102),
.Y(n_2178)
);

NOR2xp67_ASAP7_75t_SL g2179 ( 
.A(n_1928),
.B(n_1356),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2113),
.Y(n_2180)
);

AND3x1_ASAP7_75t_L g2181 ( 
.A(n_2056),
.B(n_1342),
.C(n_1325),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1961),
.B(n_1361),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1942),
.B(n_1382),
.Y(n_2183)
);

AO22x2_ASAP7_75t_L g2184 ( 
.A1(n_1947),
.A2(n_1281),
.B1(n_1364),
.B2(n_1050),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1944),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_2122),
.B(n_1397),
.Y(n_2186)
);

O2A1O1Ixp33_ASAP7_75t_L g2187 ( 
.A1(n_1908),
.A2(n_1410),
.B(n_1412),
.C(n_1405),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2136),
.B(n_2143),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2125),
.B(n_1395),
.Y(n_2189)
);

NOR2xp67_ASAP7_75t_SL g2190 ( 
.A(n_1928),
.B(n_1371),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2065),
.B(n_1372),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2159),
.B(n_1444),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_1955),
.B(n_1966),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1921),
.B(n_1378),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1946),
.Y(n_2195)
);

NAND2xp33_ASAP7_75t_SL g2196 ( 
.A(n_1898),
.B(n_1447),
.Y(n_2196)
);

BUFx6f_ASAP7_75t_L g2197 ( 
.A(n_1928),
.Y(n_2197)
);

INVxp67_ASAP7_75t_L g2198 ( 
.A(n_2117),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1895),
.B(n_1407),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_L g2200 ( 
.A(n_1916),
.B(n_1419),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_1936),
.B(n_1425),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1895),
.B(n_1894),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_2022),
.B(n_1441),
.Y(n_2203)
);

AOI22xp33_ASAP7_75t_L g2204 ( 
.A1(n_1895),
.A2(n_2003),
.B1(n_2126),
.B2(n_1876),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1957),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_2161),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_L g2207 ( 
.A1(n_2137),
.A2(n_1469),
.B1(n_1487),
.B2(n_1457),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1907),
.B(n_1429),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_1901),
.A2(n_1433),
.B1(n_1448),
.B2(n_1431),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1887),
.B(n_1453),
.Y(n_2210)
);

A2O1A1Ixp33_ASAP7_75t_L g2211 ( 
.A1(n_2048),
.A2(n_1487),
.B(n_1469),
.C(n_1418),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_1900),
.B(n_2112),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1959),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_2129),
.B(n_1454),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1960),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2153),
.B(n_1456),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2153),
.B(n_1458),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1968),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_2120),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1971),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1897),
.B(n_1909),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_2022),
.B(n_1471),
.Y(n_2222)
);

AO221x1_ASAP7_75t_L g2223 ( 
.A1(n_2123),
.A2(n_1153),
.B1(n_1158),
.B2(n_1146),
.C(n_1007),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1974),
.B(n_1461),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1982),
.B(n_1462),
.Y(n_2225)
);

NOR2xp67_ASAP7_75t_L g2226 ( 
.A(n_1951),
.B(n_2),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2127),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2133),
.B(n_1466),
.Y(n_2228)
);

CKINVDCx20_ASAP7_75t_R g2229 ( 
.A(n_1911),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_1917),
.A2(n_1481),
.B1(n_1485),
.B2(n_1474),
.Y(n_2230)
);

OAI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2060),
.A2(n_1486),
.B1(n_1494),
.B2(n_1492),
.Y(n_2231)
);

INVx3_ASAP7_75t_L g2232 ( 
.A(n_2036),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2135),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1986),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2002),
.B(n_1495),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2008),
.B(n_1496),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_1952),
.B(n_934),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2052),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_2042),
.B(n_935),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2010),
.B(n_1517),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2057),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_2042),
.B(n_936),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_1980),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2140),
.Y(n_2244)
);

AOI21xp5_ASAP7_75t_L g2245 ( 
.A1(n_1886),
.A2(n_1491),
.B(n_1476),
.Y(n_2245)
);

OAI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_1984),
.A2(n_938),
.B1(n_939),
.B2(n_937),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2061),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2109),
.B(n_950),
.Y(n_2248)
);

O2A1O1Ixp33_ASAP7_75t_L g2249 ( 
.A1(n_2014),
.A2(n_1499),
.B(n_1505),
.C(n_1498),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2005),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_2042),
.B(n_940),
.Y(n_2251)
);

INVxp67_ASAP7_75t_L g2252 ( 
.A(n_2150),
.Y(n_2252)
);

NOR3xp33_ASAP7_75t_L g2253 ( 
.A(n_1950),
.B(n_1511),
.C(n_1475),
.Y(n_2253)
);

INVxp67_ASAP7_75t_L g2254 ( 
.A(n_2162),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2007),
.Y(n_2255)
);

INVxp67_ASAP7_75t_L g2256 ( 
.A(n_2130),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_1995),
.B(n_1889),
.Y(n_2257)
);

OR2x2_ASAP7_75t_SL g2258 ( 
.A(n_2124),
.B(n_966),
.Y(n_2258)
);

NOR2xp67_ASAP7_75t_SL g2259 ( 
.A(n_2046),
.B(n_952),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2146),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_2046),
.B(n_961),
.Y(n_2261)
);

BUFx3_ASAP7_75t_L g2262 ( 
.A(n_1987),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1899),
.Y(n_2263)
);

NAND3xp33_ASAP7_75t_L g2264 ( 
.A(n_2059),
.B(n_967),
.C(n_965),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2013),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2016),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1904),
.Y(n_2267)
);

INVxp67_ASAP7_75t_L g2268 ( 
.A(n_2157),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_2085),
.B(n_968),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1919),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_L g2271 ( 
.A1(n_1930),
.A2(n_1520),
.B1(n_1146),
.B2(n_1153),
.Y(n_2271)
);

INVx8_ASAP7_75t_L g2272 ( 
.A(n_2132),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_1880),
.B(n_950),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2032),
.B(n_972),
.Y(n_2274)
);

INVxp67_ASAP7_75t_L g2275 ( 
.A(n_1988),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2043),
.B(n_974),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_1877),
.A2(n_976),
.B1(n_982),
.B2(n_978),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2050),
.B(n_985),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_1905),
.B(n_1399),
.Y(n_2279)
);

NAND3xp33_ASAP7_75t_L g2280 ( 
.A(n_1993),
.B(n_2040),
.C(n_1892),
.Y(n_2280)
);

A2O1A1Ixp33_ASAP7_75t_L g2281 ( 
.A1(n_1949),
.A2(n_1913),
.B(n_1914),
.C(n_1906),
.Y(n_2281)
);

AOI22xp33_ASAP7_75t_L g2282 ( 
.A1(n_2058),
.A2(n_1146),
.B1(n_1153),
.B2(n_1007),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2053),
.B(n_993),
.Y(n_2283)
);

AOI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2075),
.A2(n_1005),
.B1(n_1016),
.B2(n_999),
.Y(n_2284)
);

BUFx3_ASAP7_75t_L g2285 ( 
.A(n_1987),
.Y(n_2285)
);

BUFx3_ASAP7_75t_L g2286 ( 
.A(n_2082),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_2107),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_1937),
.B(n_977),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_1988),
.B(n_1998),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2028),
.Y(n_2290)
);

INVx2_ASAP7_75t_SL g2291 ( 
.A(n_2044),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2054),
.B(n_1023),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_1991),
.Y(n_2293)
);

AOI22xp33_ASAP7_75t_L g2294 ( 
.A1(n_1973),
.A2(n_1146),
.B1(n_1153),
.B2(n_1007),
.Y(n_2294)
);

AND3x1_ASAP7_75t_L g2295 ( 
.A(n_2103),
.B(n_983),
.C(n_979),
.Y(n_2295)
);

INVx3_ASAP7_75t_L g2296 ( 
.A(n_2036),
.Y(n_2296)
);

OAI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_1918),
.A2(n_996),
.B(n_984),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2029),
.Y(n_2298)
);

INVx2_ASAP7_75t_SL g2299 ( 
.A(n_2132),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2001),
.B(n_1024),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1929),
.B(n_1025),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_2046),
.B(n_1026),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2030),
.Y(n_2303)
);

NOR3xp33_ASAP7_75t_L g2304 ( 
.A(n_1958),
.B(n_1037),
.C(n_1036),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1924),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_SL g2306 ( 
.A(n_1891),
.B(n_1881),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2004),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1931),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_2037),
.B(n_1040),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_L g2310 ( 
.A(n_2000),
.B(n_1046),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_1927),
.B(n_1042),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2118),
.B(n_1049),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2009),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1875),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2026),
.B(n_1057),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2145),
.B(n_1060),
.Y(n_2316)
);

INVxp67_ASAP7_75t_SL g2317 ( 
.A(n_1882),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1870),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_R g2319 ( 
.A(n_1948),
.B(n_1066),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2017),
.B(n_1069),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_1902),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1872),
.Y(n_2322)
);

INVx2_ASAP7_75t_SL g2323 ( 
.A(n_2148),
.Y(n_2323)
);

INVxp67_ASAP7_75t_L g2324 ( 
.A(n_1994),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2027),
.B(n_956),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1873),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_1956),
.B(n_1087),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1878),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_1997),
.B(n_1093),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_1890),
.B(n_1098),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_L g2331 ( 
.A(n_2000),
.B(n_1100),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2027),
.B(n_956),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2114),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_1977),
.A2(n_1035),
.B(n_1028),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2119),
.Y(n_2335)
);

BUFx8_ASAP7_75t_L g2336 ( 
.A(n_2080),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_1989),
.B(n_1101),
.Y(n_2337)
);

INVx2_ASAP7_75t_SL g2338 ( 
.A(n_2077),
.Y(n_2338)
);

INVxp67_ASAP7_75t_L g2339 ( 
.A(n_1999),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_1989),
.B(n_1106),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_2055),
.B(n_1107),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_2107),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_1945),
.B(n_1108),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_1964),
.B(n_1114),
.Y(n_2344)
);

INVxp67_ASAP7_75t_L g2345 ( 
.A(n_2018),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2128),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_SL g2347 ( 
.A(n_1915),
.B(n_1119),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2111),
.B(n_1120),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_1990),
.B(n_1121),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1954),
.B(n_1122),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2069),
.B(n_1124),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_1990),
.B(n_1125),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_1884),
.B(n_1130),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_L g2354 ( 
.A(n_2055),
.B(n_1131),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2131),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2134),
.B(n_1135),
.Y(n_2356)
);

INVx4_ASAP7_75t_L g2357 ( 
.A(n_1910),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2138),
.Y(n_2358)
);

AOI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2072),
.A2(n_1143),
.B1(n_1152),
.B2(n_1138),
.Y(n_2359)
);

INVxp67_ASAP7_75t_SL g2360 ( 
.A(n_2039),
.Y(n_2360)
);

BUFx6f_ASAP7_75t_L g2361 ( 
.A(n_1985),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_1940),
.B(n_1156),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2021),
.Y(n_2363)
);

INVx1_ASAP7_75t_SL g2364 ( 
.A(n_2035),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2141),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2034),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2149),
.B(n_2151),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2038),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_2068),
.B(n_1160),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2079),
.A2(n_1171),
.B1(n_1177),
.B2(n_1170),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2156),
.B(n_1179),
.Y(n_2371)
);

BUFx12f_ASAP7_75t_L g2372 ( 
.A(n_2031),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_SL g2373 ( 
.A(n_2078),
.B(n_1181),
.Y(n_2373)
);

BUFx3_ASAP7_75t_L g2374 ( 
.A(n_1910),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2158),
.B(n_1187),
.Y(n_2375)
);

NOR3x1_ASAP7_75t_L g2376 ( 
.A(n_2084),
.B(n_1044),
.C(n_1041),
.Y(n_2376)
);

NOR2xp33_ASAP7_75t_L g2377 ( 
.A(n_1953),
.B(n_1192),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2064),
.Y(n_2378)
);

INVxp67_ASAP7_75t_SL g2379 ( 
.A(n_2073),
.Y(n_2379)
);

OAI22xp33_ASAP7_75t_L g2380 ( 
.A1(n_1979),
.A2(n_1493),
.B1(n_1502),
.B2(n_1484),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2062),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2011),
.B(n_1195),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_1883),
.B(n_1198),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_SL g2384 ( 
.A(n_2066),
.B(n_1205),
.Y(n_2384)
);

NAND3xp33_ASAP7_75t_L g2385 ( 
.A(n_2074),
.B(n_1209),
.C(n_1208),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2033),
.B(n_2041),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_1996),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2045),
.B(n_1214),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2063),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2012),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_2066),
.B(n_1215),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_SL g2392 ( 
.A(n_2091),
.B(n_1217),
.Y(n_2392)
);

AOI22xp33_ASAP7_75t_L g2393 ( 
.A1(n_2047),
.A2(n_1941),
.B1(n_1969),
.B2(n_2015),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_1902),
.B(n_1219),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2092),
.Y(n_2395)
);

NOR3xp33_ASAP7_75t_L g2396 ( 
.A(n_2024),
.B(n_1228),
.C(n_1227),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2097),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_1879),
.B(n_1229),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1992),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2115),
.B(n_1230),
.Y(n_2400)
);

AND2x4_ASAP7_75t_L g2401 ( 
.A(n_1983),
.B(n_1062),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2115),
.B(n_1232),
.Y(n_2402)
);

A2O1A1Ixp33_ASAP7_75t_L g2403 ( 
.A1(n_2067),
.A2(n_1078),
.B(n_1092),
.C(n_1091),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2155),
.B(n_1237),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_SL g2405 ( 
.A(n_2155),
.B(n_1250),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2049),
.B(n_1254),
.Y(n_2406)
);

NAND3xp33_ASAP7_75t_L g2407 ( 
.A(n_2147),
.B(n_1265),
.C(n_1259),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2142),
.B(n_1269),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2020),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_SL g2410 ( 
.A(n_2090),
.B(n_1271),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2144),
.B(n_2160),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_1981),
.B(n_1286),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2051),
.B(n_1287),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2101),
.Y(n_2414)
);

INVxp67_ASAP7_75t_L g2415 ( 
.A(n_1979),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_1926),
.Y(n_2416)
);

INVx8_ASAP7_75t_L g2417 ( 
.A(n_1983),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_2124),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_2108),
.B(n_1288),
.Y(n_2419)
);

AND2x6_ASAP7_75t_SL g2420 ( 
.A(n_2023),
.B(n_1117),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_1925),
.B(n_1291),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_2083),
.Y(n_2422)
);

BUFx3_ASAP7_75t_L g2423 ( 
.A(n_1920),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_1933),
.B(n_1294),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_1983),
.B(n_1888),
.Y(n_2425)
);

AND2x4_ASAP7_75t_SL g2426 ( 
.A(n_2071),
.B(n_1139),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2023),
.B(n_1034),
.Y(n_2427)
);

AOI22xp5_ASAP7_75t_L g2428 ( 
.A1(n_2154),
.A2(n_1301),
.B1(n_1304),
.B2(n_1299),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_1903),
.B(n_1305),
.Y(n_2429)
);

INVx2_ASAP7_75t_SL g2430 ( 
.A(n_1896),
.Y(n_2430)
);

NOR2xp33_ASAP7_75t_L g2431 ( 
.A(n_2006),
.B(n_1306),
.Y(n_2431)
);

INVx3_ASAP7_75t_L g2432 ( 
.A(n_1934),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1912),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_1935),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_SL g2435 ( 
.A(n_1943),
.B(n_1309),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2094),
.B(n_1311),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_1922),
.B(n_1312),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1923),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_1962),
.Y(n_2439)
);

INVx5_ASAP7_75t_L g2440 ( 
.A(n_1985),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_L g2441 ( 
.A1(n_1963),
.A2(n_1158),
.B1(n_1159),
.B2(n_1007),
.Y(n_2441)
);

INVxp67_ASAP7_75t_L g2442 ( 
.A(n_2123),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_1965),
.B(n_1315),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_1967),
.B(n_1317),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_1970),
.B(n_1318),
.Y(n_2445)
);

BUFx6f_ASAP7_75t_SL g2446 ( 
.A(n_2019),
.Y(n_2446)
);

INVx8_ASAP7_75t_L g2447 ( 
.A(n_2019),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_1972),
.B(n_1976),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_1978),
.B(n_1328),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2095),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_2025),
.B(n_1334),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2025),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2025),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_2070),
.B(n_1345),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2076),
.B(n_1343),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2081),
.B(n_1355),
.Y(n_2456)
);

OAI22xp33_ASAP7_75t_L g2457 ( 
.A1(n_2089),
.A2(n_1506),
.B1(n_1509),
.B2(n_1503),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2096),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2099),
.B(n_1358),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_L g2460 ( 
.A(n_2100),
.B(n_1365),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2104),
.B(n_1377),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2105),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2086),
.B(n_1384),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2087),
.Y(n_2464)
);

OAI221xp5_ASAP7_75t_L g2465 ( 
.A1(n_2088),
.A2(n_1393),
.B1(n_1400),
.B2(n_1391),
.C(n_1388),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2093),
.B(n_1406),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2098),
.B(n_1408),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2102),
.B(n_1034),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2106),
.B(n_1414),
.Y(n_2469)
);

NOR2xp33_ASAP7_75t_L g2470 ( 
.A(n_1908),
.B(n_1415),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_1975),
.B(n_1417),
.Y(n_2471)
);

INVxp67_ASAP7_75t_L g2472 ( 
.A(n_1871),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2152),
.B(n_1139),
.Y(n_2473)
);

INVx1_ASAP7_75t_SL g2474 ( 
.A(n_2152),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_1975),
.B(n_1420),
.Y(n_2475)
);

AND2x4_ASAP7_75t_L g2476 ( 
.A(n_2121),
.B(n_1129),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_1893),
.Y(n_2477)
);

NOR2xp67_ASAP7_75t_L g2478 ( 
.A(n_2116),
.B(n_3),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_1975),
.B(n_1421),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_1975),
.B(n_1422),
.Y(n_2480)
);

OR2x2_ASAP7_75t_L g2481 ( 
.A(n_2152),
.B(n_1426),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_1975),
.B(n_1434),
.Y(n_2482)
);

OAI22xp33_ASAP7_75t_L g2483 ( 
.A1(n_1885),
.A2(n_1478),
.B1(n_1479),
.B2(n_1468),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_1975),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_1975),
.B(n_1436),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_1975),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_1975),
.B(n_1440),
.Y(n_2487)
);

AOI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_1885),
.A2(n_1446),
.B1(n_1480),
.B2(n_1445),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_1893),
.Y(n_2489)
);

NAND3xp33_ASAP7_75t_L g2490 ( 
.A(n_1885),
.B(n_1514),
.C(n_1482),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_1975),
.B(n_1524),
.Y(n_2491)
);

AOI22xp5_ASAP7_75t_L g2492 ( 
.A1(n_1885),
.A2(n_1145),
.B1(n_1165),
.B2(n_1134),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_1975),
.B(n_1182),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_SL g2494 ( 
.A(n_1885),
.B(n_1158),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_1975),
.B(n_1197),
.Y(n_2495)
);

A2O1A1Ixp33_ASAP7_75t_L g2496 ( 
.A1(n_2048),
.A2(n_1249),
.B(n_1262),
.C(n_1226),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_1975),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_1885),
.B(n_1158),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_1975),
.B(n_1282),
.Y(n_2499)
);

AO22x2_ASAP7_75t_L g2500 ( 
.A1(n_2152),
.A2(n_1307),
.B1(n_1327),
.B2(n_1284),
.Y(n_2500)
);

NOR2x1p5_ASAP7_75t_L g2501 ( 
.A(n_1915),
.B(n_1329),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_L g2502 ( 
.A1(n_1895),
.A2(n_1204),
.B1(n_1285),
.B2(n_1159),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_1893),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_1975),
.B(n_1331),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_2161),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_1975),
.B(n_1339),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_1893),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_1885),
.B(n_1159),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_SL g2509 ( 
.A(n_2152),
.B(n_1167),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2152),
.B(n_1167),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_1975),
.B(n_1351),
.Y(n_2511)
);

OAI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_1975),
.A2(n_1362),
.B1(n_1363),
.B2(n_1352),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_1975),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_1975),
.Y(n_2514)
);

OAI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_1975),
.A2(n_1390),
.B1(n_1398),
.B2(n_1368),
.Y(n_2515)
);

NOR2xp33_ASAP7_75t_L g2516 ( 
.A(n_1908),
.B(n_1375),
.Y(n_2516)
);

INVxp33_ASAP7_75t_L g2517 ( 
.A(n_1871),
.Y(n_2517)
);

NOR2xp67_ASAP7_75t_L g2518 ( 
.A(n_2116),
.B(n_4),
.Y(n_2518)
);

OAI22x1_ASAP7_75t_SL g2519 ( 
.A1(n_1951),
.A2(n_1424),
.B1(n_1428),
.B2(n_1416),
.Y(n_2519)
);

INVx1_ASAP7_75t_SL g2520 ( 
.A(n_2152),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_1975),
.B(n_1432),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2152),
.B(n_1375),
.Y(n_2522)
);

BUFx6f_ASAP7_75t_L g2523 ( 
.A(n_1928),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_SL g2524 ( 
.A(n_1885),
.B(n_1159),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_1975),
.B(n_1435),
.Y(n_2525)
);

INVx2_ASAP7_75t_SL g2526 ( 
.A(n_2121),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_1975),
.B(n_1437),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_1975),
.B(n_1449),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_1975),
.B(n_1455),
.Y(n_2529)
);

OAI22xp5_ASAP7_75t_L g2530 ( 
.A1(n_1975),
.A2(n_1464),
.B1(n_1465),
.B2(n_1459),
.Y(n_2530)
);

AOI22xp33_ASAP7_75t_L g2531 ( 
.A1(n_1895),
.A2(n_1285),
.B1(n_1204),
.B2(n_1473),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_1975),
.B(n_1490),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2164),
.B(n_1507),
.Y(n_2533)
);

OAI21xp5_ASAP7_75t_L g2534 ( 
.A1(n_2281),
.A2(n_2245),
.B(n_2211),
.Y(n_2534)
);

AOI21xp5_ASAP7_75t_L g2535 ( 
.A1(n_2221),
.A2(n_1190),
.B(n_1189),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2484),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2486),
.Y(n_2537)
);

AOI21xp5_ASAP7_75t_L g2538 ( 
.A1(n_2263),
.A2(n_1190),
.B(n_1189),
.Y(n_2538)
);

BUFx3_ASAP7_75t_L g2539 ( 
.A(n_2229),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2497),
.B(n_2513),
.Y(n_2540)
);

AOI21xp5_ASAP7_75t_L g2541 ( 
.A1(n_2267),
.A2(n_1389),
.B(n_1386),
.Y(n_2541)
);

AOI21xp5_ASAP7_75t_L g2542 ( 
.A1(n_2270),
.A2(n_1389),
.B(n_1386),
.Y(n_2542)
);

INVxp67_ASAP7_75t_L g2543 ( 
.A(n_2474),
.Y(n_2543)
);

AOI21xp5_ASAP7_75t_L g2544 ( 
.A1(n_2168),
.A2(n_2180),
.B(n_2172),
.Y(n_2544)
);

AOI21xp5_ASAP7_75t_L g2545 ( 
.A1(n_2219),
.A2(n_1442),
.B(n_1396),
.Y(n_2545)
);

OAI22x1_ASAP7_75t_L g2546 ( 
.A1(n_2442),
.A2(n_1442),
.B1(n_1488),
.B2(n_1396),
.Y(n_2546)
);

AOI21xp5_ASAP7_75t_L g2547 ( 
.A1(n_2227),
.A2(n_1488),
.B(n_1285),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_2233),
.A2(n_1285),
.B(n_1204),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2514),
.B(n_1300),
.Y(n_2549)
);

O2A1O1Ixp33_ASAP7_75t_SL g2550 ( 
.A1(n_2494),
.A2(n_2498),
.B(n_2524),
.C(n_2508),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2257),
.B(n_1300),
.Y(n_2551)
);

AOI21xp5_ASAP7_75t_L g2552 ( 
.A1(n_2244),
.A2(n_2477),
.B(n_2260),
.Y(n_2552)
);

AOI21xp5_ASAP7_75t_L g2553 ( 
.A1(n_2489),
.A2(n_1110),
.B(n_1105),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2198),
.B(n_1300),
.Y(n_2554)
);

AOI21xp5_ASAP7_75t_L g2555 ( 
.A1(n_2503),
.A2(n_1110),
.B(n_1105),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2238),
.Y(n_2556)
);

AOI21xp5_ASAP7_75t_L g2557 ( 
.A1(n_2507),
.A2(n_1110),
.B(n_1105),
.Y(n_2557)
);

NOR2xp67_ASAP7_75t_L g2558 ( 
.A(n_2372),
.B(n_4),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2252),
.B(n_2254),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2169),
.B(n_1300),
.Y(n_2560)
);

NAND2x1p5_ASAP7_75t_L g2561 ( 
.A(n_2520),
.B(n_1369),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2173),
.B(n_2177),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2185),
.B(n_1319),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2195),
.B(n_1319),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2241),
.Y(n_2565)
);

AOI21xp5_ASAP7_75t_L g2566 ( 
.A1(n_2236),
.A2(n_2314),
.B(n_2240),
.Y(n_2566)
);

AOI21xp5_ASAP7_75t_L g2567 ( 
.A1(n_2210),
.A2(n_1409),
.B(n_1369),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2247),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2205),
.B(n_1319),
.Y(n_2569)
);

INVx4_ASAP7_75t_L g2570 ( 
.A(n_2272),
.Y(n_2570)
);

NOR2xp33_ASAP7_75t_L g2571 ( 
.A(n_2256),
.B(n_1439),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2213),
.B(n_1319),
.Y(n_2572)
);

AOI21xp5_ASAP7_75t_L g2573 ( 
.A1(n_2224),
.A2(n_1409),
.B(n_1369),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2215),
.B(n_1319),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2218),
.Y(n_2575)
);

AOI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2225),
.A2(n_1409),
.B(n_1369),
.Y(n_2576)
);

OAI21xp5_ASAP7_75t_L g2577 ( 
.A1(n_2334),
.A2(n_1338),
.B(n_1319),
.Y(n_2577)
);

INVx3_ASAP7_75t_L g2578 ( 
.A(n_2197),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2250),
.Y(n_2579)
);

NOR3xp33_ASAP7_75t_L g2580 ( 
.A(n_2280),
.B(n_1439),
.C(n_1338),
.Y(n_2580)
);

O2A1O1Ixp33_ASAP7_75t_L g2581 ( 
.A1(n_2403),
.A2(n_1338),
.B(n_7),
.C(n_5),
.Y(n_2581)
);

A2O1A1Ixp33_ASAP7_75t_L g2582 ( 
.A1(n_2249),
.A2(n_2187),
.B(n_2297),
.C(n_2204),
.Y(n_2582)
);

BUFx2_ASAP7_75t_L g2583 ( 
.A(n_2206),
.Y(n_2583)
);

INVx4_ASAP7_75t_L g2584 ( 
.A(n_2272),
.Y(n_2584)
);

OR2x2_ASAP7_75t_L g2585 ( 
.A(n_2183),
.B(n_5),
.Y(n_2585)
);

AOI21xp5_ASAP7_75t_L g2586 ( 
.A1(n_2235),
.A2(n_1467),
.B(n_1409),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2220),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2228),
.B(n_1338),
.Y(n_2588)
);

BUFx4f_ASAP7_75t_L g2589 ( 
.A(n_2163),
.Y(n_2589)
);

AOI21xp5_ASAP7_75t_L g2590 ( 
.A1(n_2386),
.A2(n_1504),
.B(n_1467),
.Y(n_2590)
);

BUFx6f_ASAP7_75t_L g2591 ( 
.A(n_2287),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2234),
.B(n_2193),
.Y(n_2592)
);

AOI21xp5_ASAP7_75t_L g2593 ( 
.A1(n_2367),
.A2(n_1504),
.B(n_1467),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2255),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2166),
.B(n_1338),
.Y(n_2595)
);

AOI21xp5_ASAP7_75t_L g2596 ( 
.A1(n_2274),
.A2(n_1504),
.B(n_1467),
.Y(n_2596)
);

O2A1O1Ixp33_ASAP7_75t_L g2597 ( 
.A1(n_2496),
.A2(n_1338),
.B(n_8),
.C(n_6),
.Y(n_2597)
);

AOI21xp5_ASAP7_75t_L g2598 ( 
.A1(n_2276),
.A2(n_1504),
.B(n_6),
.Y(n_2598)
);

BUFx4f_ASAP7_75t_L g2599 ( 
.A(n_2188),
.Y(n_2599)
);

O2A1O1Ixp33_ASAP7_75t_L g2600 ( 
.A1(n_2306),
.A2(n_10),
.B(n_7),
.C(n_9),
.Y(n_2600)
);

INVx8_ASAP7_75t_L g2601 ( 
.A(n_2417),
.Y(n_2601)
);

BUFx3_ASAP7_75t_L g2602 ( 
.A(n_2336),
.Y(n_2602)
);

AOI21x1_ASAP7_75t_L g2603 ( 
.A1(n_2425),
.A2(n_7),
.B(n_9),
.Y(n_2603)
);

AOI21xp5_ASAP7_75t_L g2604 ( 
.A1(n_2278),
.A2(n_9),
.B(n_10),
.Y(n_2604)
);

AOI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2283),
.A2(n_11),
.B(n_12),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2505),
.B(n_12),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2201),
.B(n_13),
.Y(n_2607)
);

O2A1O1Ixp33_ASAP7_75t_L g2608 ( 
.A1(n_2191),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_2608)
);

O2A1O1Ixp33_ASAP7_75t_L g2609 ( 
.A1(n_2427),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_2609)
);

OR2x2_ASAP7_75t_L g2610 ( 
.A(n_2472),
.B(n_17),
.Y(n_2610)
);

AOI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2292),
.A2(n_17),
.B(n_18),
.Y(n_2611)
);

OAI22xp5_ASAP7_75t_L g2612 ( 
.A1(n_2493),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_SL g2613 ( 
.A(n_2483),
.B(n_20),
.Y(n_2613)
);

INVxp67_ASAP7_75t_L g2614 ( 
.A(n_2212),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2526),
.B(n_20),
.Y(n_2615)
);

AOI21xp5_ASAP7_75t_L g2616 ( 
.A1(n_2327),
.A2(n_19),
.B(n_20),
.Y(n_2616)
);

AOI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2329),
.A2(n_21),
.B(n_22),
.Y(n_2617)
);

AOI21xp5_ASAP7_75t_L g2618 ( 
.A1(n_2350),
.A2(n_21),
.B(n_22),
.Y(n_2618)
);

HB1xp67_ASAP7_75t_L g2619 ( 
.A(n_2364),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_SL g2620 ( 
.A(n_2422),
.B(n_21),
.Y(n_2620)
);

AOI22xp5_ASAP7_75t_L g2621 ( 
.A1(n_2214),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_2621)
);

OAI21xp5_ASAP7_75t_L g2622 ( 
.A1(n_2431),
.A2(n_23),
.B(n_24),
.Y(n_2622)
);

INVx3_ASAP7_75t_L g2623 ( 
.A(n_2197),
.Y(n_2623)
);

AOI21xp5_ASAP7_75t_L g2624 ( 
.A1(n_2411),
.A2(n_23),
.B(n_24),
.Y(n_2624)
);

AOI21xp5_ASAP7_75t_L g2625 ( 
.A1(n_2312),
.A2(n_25),
.B(n_26),
.Y(n_2625)
);

O2A1O1Ixp33_ASAP7_75t_L g2626 ( 
.A1(n_2182),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_2626)
);

CKINVDCx6p67_ASAP7_75t_R g2627 ( 
.A(n_2165),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2316),
.A2(n_25),
.B(n_26),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2495),
.B(n_27),
.Y(n_2629)
);

AOI21xp5_ASAP7_75t_L g2630 ( 
.A1(n_2499),
.A2(n_28),
.B(n_29),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2265),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2504),
.B(n_28),
.Y(n_2632)
);

AOI21xp5_ASAP7_75t_L g2633 ( 
.A1(n_2506),
.A2(n_29),
.B(n_30),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2511),
.B(n_30),
.Y(n_2634)
);

AOI21xp5_ASAP7_75t_L g2635 ( 
.A1(n_2521),
.A2(n_30),
.B(n_31),
.Y(n_2635)
);

AOI21xp5_ASAP7_75t_L g2636 ( 
.A1(n_2525),
.A2(n_31),
.B(n_32),
.Y(n_2636)
);

A2O1A1Ixp33_ASAP7_75t_L g2637 ( 
.A1(n_2395),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_2637)
);

INVx1_ASAP7_75t_SL g2638 ( 
.A(n_2517),
.Y(n_2638)
);

OAI21xp5_ASAP7_75t_L g2639 ( 
.A1(n_2208),
.A2(n_32),
.B(n_33),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2527),
.B(n_33),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2528),
.B(n_2529),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2266),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2532),
.B(n_34),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_SL g2644 ( 
.A(n_2246),
.B(n_35),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2373),
.B(n_35),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2290),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2471),
.B(n_34),
.Y(n_2647)
);

O2A1O1Ixp33_ASAP7_75t_L g2648 ( 
.A1(n_2268),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_2648)
);

AO21x1_ASAP7_75t_L g2649 ( 
.A1(n_2202),
.A2(n_604),
.B(n_603),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2298),
.Y(n_2650)
);

A2O1A1Ixp33_ASAP7_75t_L g2651 ( 
.A1(n_2397),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_2651)
);

OAI22xp5_ASAP7_75t_L g2652 ( 
.A1(n_2303),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_2652)
);

AOI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_2392),
.A2(n_38),
.B(n_39),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2475),
.B(n_39),
.Y(n_2654)
);

AOI21xp5_ASAP7_75t_L g2655 ( 
.A1(n_2479),
.A2(n_40),
.B(n_41),
.Y(n_2655)
);

AOI21xp5_ASAP7_75t_L g2656 ( 
.A1(n_2480),
.A2(n_40),
.B(n_41),
.Y(n_2656)
);

BUFx6f_ASAP7_75t_L g2657 ( 
.A(n_2287),
.Y(n_2657)
);

OR2x2_ASAP7_75t_L g2658 ( 
.A(n_2258),
.B(n_40),
.Y(n_2658)
);

OAI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2305),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2659)
);

BUFx3_ASAP7_75t_L g2660 ( 
.A(n_2336),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2482),
.B(n_42),
.Y(n_2661)
);

OAI21xp5_ASAP7_75t_L g2662 ( 
.A1(n_2308),
.A2(n_2378),
.B(n_2389),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2318),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2345),
.B(n_42),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2322),
.Y(n_2665)
);

AOI21xp5_ASAP7_75t_L g2666 ( 
.A1(n_2485),
.A2(n_43),
.B(n_44),
.Y(n_2666)
);

OAI22xp5_ASAP7_75t_L g2667 ( 
.A1(n_2500),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2667)
);

AOI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2189),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2668)
);

AOI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2487),
.A2(n_45),
.B(n_46),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_SL g2670 ( 
.A(n_2287),
.B(n_47),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2491),
.B(n_46),
.Y(n_2671)
);

NOR2xp33_ASAP7_75t_L g2672 ( 
.A(n_2275),
.B(n_48),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2216),
.B(n_48),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_L g2674 ( 
.A(n_2289),
.B(n_49),
.Y(n_2674)
);

INVx4_ASAP7_75t_L g2675 ( 
.A(n_2417),
.Y(n_2675)
);

AOI21xp5_ASAP7_75t_L g2676 ( 
.A1(n_2356),
.A2(n_49),
.B(n_50),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_L g2677 ( 
.A(n_2324),
.B(n_50),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2326),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2217),
.B(n_51),
.Y(n_2679)
);

O2A1O1Ixp33_ASAP7_75t_L g2680 ( 
.A1(n_2339),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2328),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2415),
.B(n_51),
.Y(n_2682)
);

AOI21xp5_ASAP7_75t_L g2683 ( 
.A1(n_2371),
.A2(n_52),
.B(n_54),
.Y(n_2683)
);

A2O1A1Ixp33_ASAP7_75t_L g2684 ( 
.A1(n_2478),
.A2(n_55),
.B(n_52),
.C(n_54),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2248),
.B(n_55),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2194),
.B(n_56),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2200),
.B(n_56),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2512),
.B(n_2530),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_L g2689 ( 
.A(n_2360),
.B(n_56),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2333),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2335),
.Y(n_2691)
);

AOI21xp5_ASAP7_75t_L g2692 ( 
.A1(n_2375),
.A2(n_57),
.B(n_58),
.Y(n_2692)
);

OAI21x1_ASAP7_75t_L g2693 ( 
.A1(n_2452),
.A2(n_605),
.B(n_603),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2515),
.B(n_57),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2288),
.B(n_57),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2288),
.B(n_59),
.Y(n_2696)
);

OAI21xp33_ASAP7_75t_L g2697 ( 
.A1(n_2269),
.A2(n_59),
.B(n_60),
.Y(n_2697)
);

AOI21xp5_ASAP7_75t_L g2698 ( 
.A1(n_2382),
.A2(n_2448),
.B(n_2437),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_SL g2699 ( 
.A(n_2342),
.B(n_61),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2209),
.B(n_60),
.Y(n_2700)
);

INVx2_ASAP7_75t_SL g2701 ( 
.A(n_2262),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2342),
.B(n_62),
.Y(n_2702)
);

OAI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_2346),
.A2(n_2358),
.B(n_2355),
.Y(n_2703)
);

AOI21xp5_ASAP7_75t_L g2704 ( 
.A1(n_2455),
.A2(n_61),
.B(n_62),
.Y(n_2704)
);

AOI21xp33_ASAP7_75t_L g2705 ( 
.A1(n_2300),
.A2(n_61),
.B(n_62),
.Y(n_2705)
);

AOI22xp33_ASAP7_75t_L g2706 ( 
.A1(n_2396),
.A2(n_2304),
.B1(n_2273),
.B2(n_2196),
.Y(n_2706)
);

AOI21xp5_ASAP7_75t_L g2707 ( 
.A1(n_2456),
.A2(n_63),
.B(n_64),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2342),
.B(n_64),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2230),
.B(n_63),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2500),
.B(n_63),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2365),
.Y(n_2711)
);

BUFx6f_ASAP7_75t_L g2712 ( 
.A(n_2197),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2330),
.B(n_64),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2293),
.Y(n_2714)
);

AOI21xp5_ASAP7_75t_L g2715 ( 
.A1(n_2459),
.A2(n_2461),
.B(n_2438),
.Y(n_2715)
);

AOI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2433),
.A2(n_65),
.B(n_66),
.Y(n_2716)
);

CKINVDCx20_ASAP7_75t_R g2717 ( 
.A(n_2319),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2343),
.B(n_66),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2344),
.B(n_67),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2307),
.Y(n_2720)
);

INVx4_ASAP7_75t_L g2721 ( 
.A(n_2285),
.Y(n_2721)
);

NOR2xp33_ASAP7_75t_L g2722 ( 
.A(n_2279),
.B(n_67),
.Y(n_2722)
);

O2A1O1Ixp33_ASAP7_75t_L g2723 ( 
.A1(n_2348),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2184),
.B(n_68),
.Y(n_2724)
);

BUFx4f_ASAP7_75t_L g2725 ( 
.A(n_2165),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2351),
.B(n_68),
.Y(n_2726)
);

OAI21xp5_ASAP7_75t_L g2727 ( 
.A1(n_2271),
.A2(n_69),
.B(n_70),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2470),
.B(n_70),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2313),
.Y(n_2729)
);

AOI22xp5_ASAP7_75t_L g2730 ( 
.A1(n_2295),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_2730)
);

AO21x1_ASAP7_75t_L g2731 ( 
.A1(n_2223),
.A2(n_607),
.B(n_606),
.Y(n_2731)
);

HB1xp67_ASAP7_75t_L g2732 ( 
.A(n_2178),
.Y(n_2732)
);

OAI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2385),
.A2(n_74),
.B(n_75),
.Y(n_2733)
);

HB1xp67_ASAP7_75t_L g2734 ( 
.A(n_2178),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_SL g2735 ( 
.A(n_2380),
.B(n_75),
.Y(n_2735)
);

NOR3xp33_ASAP7_75t_L g2736 ( 
.A(n_2253),
.B(n_76),
.C(n_75),
.Y(n_2736)
);

AOI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2363),
.A2(n_2368),
.B(n_2366),
.Y(n_2737)
);

HB1xp67_ASAP7_75t_L g2738 ( 
.A(n_2192),
.Y(n_2738)
);

OAI22xp5_ASAP7_75t_L g2739 ( 
.A1(n_2393),
.A2(n_77),
.B1(n_74),
.B2(n_76),
.Y(n_2739)
);

BUFx6f_ASAP7_75t_L g2740 ( 
.A(n_2523),
.Y(n_2740)
);

OAI21xp5_ASAP7_75t_L g2741 ( 
.A1(n_2353),
.A2(n_77),
.B(n_78),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2381),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2492),
.B(n_77),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_SL g2744 ( 
.A(n_2347),
.B(n_2509),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2481),
.B(n_78),
.Y(n_2745)
);

AND2x6_ASAP7_75t_L g2746 ( 
.A(n_2523),
.B(n_79),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_SL g2747 ( 
.A(n_2490),
.B(n_80),
.Y(n_2747)
);

AOI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2416),
.A2(n_79),
.B(n_80),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2476),
.B(n_79),
.Y(n_2749)
);

INVx3_ASAP7_75t_L g2750 ( 
.A(n_2523),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2434),
.A2(n_81),
.B(n_82),
.Y(n_2751)
);

BUFx2_ASAP7_75t_L g2752 ( 
.A(n_2181),
.Y(n_2752)
);

BUFx4f_ASAP7_75t_L g2753 ( 
.A(n_2338),
.Y(n_2753)
);

AOI22xp5_ASAP7_75t_L g2754 ( 
.A1(n_2184),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2476),
.B(n_82),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2299),
.B(n_83),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2361),
.Y(n_2757)
);

AOI21xp5_ASAP7_75t_L g2758 ( 
.A1(n_2439),
.A2(n_83),
.B(n_84),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2390),
.B(n_84),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2473),
.B(n_2510),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2462),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2464),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2432),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2321),
.Y(n_2764)
);

O2A1O1Ixp33_ASAP7_75t_L g2765 ( 
.A1(n_2320),
.A2(n_2311),
.B(n_2315),
.C(n_2301),
.Y(n_2765)
);

AOI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2443),
.A2(n_84),
.B(n_85),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2522),
.B(n_85),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_SL g2768 ( 
.A(n_2457),
.B(n_87),
.Y(n_2768)
);

AOI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2444),
.A2(n_86),
.B(n_88),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2468),
.B(n_86),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2432),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2232),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2445),
.A2(n_86),
.B(n_88),
.Y(n_2773)
);

NOR3xp33_ASAP7_75t_L g2774 ( 
.A(n_2264),
.B(n_90),
.C(n_89),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2401),
.Y(n_2775)
);

OAI21xp5_ASAP7_75t_L g2776 ( 
.A1(n_2383),
.A2(n_88),
.B(n_89),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2231),
.B(n_2516),
.Y(n_2777)
);

AOI21xp5_ASAP7_75t_L g2778 ( 
.A1(n_2449),
.A2(n_2199),
.B(n_2463),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2176),
.B(n_89),
.Y(n_2779)
);

BUFx6f_ASAP7_75t_L g2780 ( 
.A(n_2361),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2414),
.B(n_91),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2376),
.B(n_91),
.Y(n_2782)
);

AOI22xp5_ASAP7_75t_L g2783 ( 
.A1(n_2488),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2401),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2399),
.B(n_92),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2186),
.B(n_92),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2232),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2466),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_SL g2789 ( 
.A(n_2243),
.B(n_93),
.Y(n_2789)
);

A2O1A1Ixp33_ASAP7_75t_L g2790 ( 
.A1(n_2518),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2277),
.B(n_94),
.Y(n_2791)
);

AOI21xp5_ASAP7_75t_L g2792 ( 
.A1(n_2469),
.A2(n_94),
.B(n_95),
.Y(n_2792)
);

AOI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2419),
.A2(n_95),
.B(n_96),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2237),
.B(n_96),
.Y(n_2794)
);

AOI21xp5_ASAP7_75t_L g2795 ( 
.A1(n_2171),
.A2(n_96),
.B(n_97),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2379),
.B(n_98),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_SL g2797 ( 
.A(n_2384),
.B(n_2446),
.Y(n_2797)
);

NOR2xp33_ASAP7_75t_SL g2798 ( 
.A(n_2446),
.B(n_98),
.Y(n_2798)
);

INVx3_ASAP7_75t_L g2799 ( 
.A(n_2321),
.Y(n_2799)
);

OAI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2174),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_2800)
);

INVx4_ASAP7_75t_L g2801 ( 
.A(n_2447),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_SL g2802 ( 
.A(n_2447),
.B(n_99),
.Y(n_2802)
);

O2A1O1Ixp33_ASAP7_75t_L g2803 ( 
.A1(n_2362),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2296),
.Y(n_2804)
);

A2O1A1Ixp33_ASAP7_75t_L g2805 ( 
.A1(n_2207),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2175),
.A2(n_2388),
.B(n_2421),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2369),
.B(n_101),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2408),
.B(n_103),
.Y(n_2808)
);

INVx1_ASAP7_75t_SL g2809 ( 
.A(n_2286),
.Y(n_2809)
);

AOI21xp5_ASAP7_75t_L g2810 ( 
.A1(n_2413),
.A2(n_103),
.B(n_104),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2317),
.B(n_103),
.Y(n_2811)
);

NOR2x2_ASAP7_75t_L g2812 ( 
.A(n_2418),
.B(n_104),
.Y(n_2812)
);

HB1xp67_ASAP7_75t_L g2813 ( 
.A(n_2291),
.Y(n_2813)
);

AOI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2458),
.A2(n_104),
.B(n_105),
.Y(n_2814)
);

AND2x2_ASAP7_75t_L g2815 ( 
.A(n_2370),
.B(n_105),
.Y(n_2815)
);

NAND2xp33_ASAP7_75t_SL g2816 ( 
.A(n_2179),
.B(n_105),
.Y(n_2816)
);

AO21x1_ASAP7_75t_L g2817 ( 
.A1(n_2453),
.A2(n_609),
.B(n_608),
.Y(n_2817)
);

AOI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2398),
.A2(n_2412),
.B(n_2410),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2325),
.B(n_106),
.Y(n_2819)
);

AND2x4_ASAP7_75t_L g2820 ( 
.A(n_2423),
.B(n_106),
.Y(n_2820)
);

OAI21xp5_ASAP7_75t_L g2821 ( 
.A1(n_2407),
.A2(n_106),
.B(n_107),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2284),
.B(n_107),
.Y(n_2822)
);

OAI21xp5_ASAP7_75t_L g2823 ( 
.A1(n_2282),
.A2(n_107),
.B(n_108),
.Y(n_2823)
);

AND2x4_ASAP7_75t_L g2824 ( 
.A(n_2409),
.B(n_108),
.Y(n_2824)
);

O2A1O1Ixp5_ASAP7_75t_L g2825 ( 
.A1(n_2203),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_2825)
);

AOI22xp5_ASAP7_75t_L g2826 ( 
.A1(n_2170),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_R g2827 ( 
.A(n_2387),
.B(n_111),
.Y(n_2827)
);

INVxp67_ASAP7_75t_L g2828 ( 
.A(n_2332),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2359),
.B(n_112),
.Y(n_2829)
);

O2A1O1Ixp33_ASAP7_75t_L g2830 ( 
.A1(n_2465),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_2830)
);

INVx3_ASAP7_75t_L g2831 ( 
.A(n_2296),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2436),
.B(n_114),
.Y(n_2832)
);

NOR2xp33_ASAP7_75t_L g2833 ( 
.A(n_2310),
.B(n_114),
.Y(n_2833)
);

AOI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2222),
.A2(n_115),
.B(n_116),
.Y(n_2834)
);

O2A1O1Ixp33_ASAP7_75t_L g2835 ( 
.A1(n_2337),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2424),
.B(n_2309),
.Y(n_2836)
);

NOR2xp33_ASAP7_75t_L g2837 ( 
.A(n_2331),
.B(n_116),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2377),
.B(n_117),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2406),
.B(n_118),
.Y(n_2839)
);

AOI22xp5_ASAP7_75t_L g2840 ( 
.A1(n_2451),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_2840)
);

AOI22xp5_ASAP7_75t_L g2841 ( 
.A1(n_2341),
.A2(n_2354),
.B1(n_2501),
.B2(n_2519),
.Y(n_2841)
);

BUFx6f_ASAP7_75t_L g2842 ( 
.A(n_2361),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2428),
.B(n_2454),
.Y(n_2843)
);

HB1xp67_ASAP7_75t_L g2844 ( 
.A(n_2374),
.Y(n_2844)
);

AOI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2429),
.A2(n_2242),
.B(n_2239),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2460),
.B(n_119),
.Y(n_2846)
);

O2A1O1Ixp33_ASAP7_75t_L g2847 ( 
.A1(n_2340),
.A2(n_122),
.B(n_119),
.C(n_121),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2394),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2400),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2402),
.Y(n_2850)
);

AOI21xp5_ASAP7_75t_L g2851 ( 
.A1(n_2251),
.A2(n_2302),
.B(n_2261),
.Y(n_2851)
);

AOI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2435),
.A2(n_121),
.B(n_122),
.Y(n_2852)
);

INVx3_ASAP7_75t_L g2853 ( 
.A(n_2440),
.Y(n_2853)
);

AOI22xp33_ASAP7_75t_L g2854 ( 
.A1(n_2349),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2352),
.B(n_123),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_SL g2856 ( 
.A(n_2440),
.B(n_125),
.Y(n_2856)
);

BUFx2_ASAP7_75t_L g2857 ( 
.A(n_2357),
.Y(n_2857)
);

BUFx8_ASAP7_75t_L g2858 ( 
.A(n_2323),
.Y(n_2858)
);

AOI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_2467),
.A2(n_124),
.B(n_125),
.Y(n_2859)
);

AO21x1_ASAP7_75t_L g2860 ( 
.A1(n_2420),
.A2(n_610),
.B(n_608),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2357),
.B(n_124),
.Y(n_2861)
);

INVx3_ASAP7_75t_L g2862 ( 
.A(n_2440),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2426),
.B(n_124),
.Y(n_2863)
);

AOI21xp5_ASAP7_75t_L g2864 ( 
.A1(n_2531),
.A2(n_126),
.B(n_127),
.Y(n_2864)
);

AND2x4_ASAP7_75t_L g2865 ( 
.A(n_2404),
.B(n_126),
.Y(n_2865)
);

NOR2x1_ASAP7_75t_L g2866 ( 
.A(n_2226),
.B(n_126),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_SL g2867 ( 
.A(n_2167),
.B(n_128),
.Y(n_2867)
);

OAI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2502),
.A2(n_2294),
.B1(n_2450),
.B2(n_2405),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2167),
.B(n_128),
.Y(n_2869)
);

INVx3_ASAP7_75t_L g2870 ( 
.A(n_2167),
.Y(n_2870)
);

INVx1_ASAP7_75t_SL g2871 ( 
.A(n_2391),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2430),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2190),
.B(n_127),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2259),
.B(n_127),
.Y(n_2874)
);

AOI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2441),
.A2(n_128),
.B(n_129),
.Y(n_2875)
);

NOR2xp33_ASAP7_75t_L g2876 ( 
.A(n_2167),
.B(n_129),
.Y(n_2876)
);

OAI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2221),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2281),
.A2(n_130),
.B(n_131),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2281),
.A2(n_131),
.B(n_132),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2164),
.B(n_132),
.Y(n_2880)
);

NOR2xp33_ASAP7_75t_L g2881 ( 
.A(n_2198),
.B(n_133),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2164),
.B(n_133),
.Y(n_2882)
);

AOI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2500),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_2883)
);

O2A1O1Ixp33_ASAP7_75t_L g2884 ( 
.A1(n_2403),
.A2(n_137),
.B(n_134),
.C(n_136),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2164),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2164),
.B(n_136),
.Y(n_2886)
);

NOR2xp33_ASAP7_75t_L g2887 ( 
.A(n_2198),
.B(n_136),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2164),
.B(n_137),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2164),
.B(n_138),
.Y(n_2889)
);

AND2x2_ASAP7_75t_L g2890 ( 
.A(n_2257),
.B(n_138),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2281),
.A2(n_138),
.B(n_139),
.Y(n_2891)
);

OAI21x1_ASAP7_75t_L g2892 ( 
.A1(n_2263),
.A2(n_611),
.B(n_610),
.Y(n_2892)
);

NAND2xp33_ASAP7_75t_L g2893 ( 
.A(n_2287),
.B(n_140),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2164),
.B(n_139),
.Y(n_2894)
);

AOI21xp5_ASAP7_75t_L g2895 ( 
.A1(n_2281),
.A2(n_139),
.B(n_140),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_SL g2896 ( 
.A(n_2163),
.B(n_141),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_L g2897 ( 
.A(n_2198),
.B(n_140),
.Y(n_2897)
);

OR2x2_ASAP7_75t_L g2898 ( 
.A(n_2474),
.B(n_141),
.Y(n_2898)
);

OAI21xp5_ASAP7_75t_L g2899 ( 
.A1(n_2281),
.A2(n_142),
.B(n_143),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2164),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2164),
.Y(n_2901)
);

OAI321xp33_ASAP7_75t_L g2902 ( 
.A1(n_2442),
.A2(n_144),
.A3(n_146),
.B1(n_142),
.B2(n_143),
.C(n_145),
.Y(n_2902)
);

A2O1A1Ixp33_ASAP7_75t_L g2903 ( 
.A1(n_2245),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_2903)
);

BUFx4f_ASAP7_75t_L g2904 ( 
.A(n_2372),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2164),
.Y(n_2905)
);

AOI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2281),
.A2(n_144),
.B(n_146),
.Y(n_2906)
);

AOI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2281),
.A2(n_147),
.B(n_148),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2198),
.B(n_147),
.Y(n_2908)
);

NAND2x1p5_ASAP7_75t_L g2909 ( 
.A(n_2474),
.B(n_147),
.Y(n_2909)
);

BUFx6f_ASAP7_75t_L g2910 ( 
.A(n_2287),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_SL g2911 ( 
.A(n_2163),
.B(n_148),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2164),
.Y(n_2912)
);

OAI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2281),
.A2(n_149),
.B(n_150),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2164),
.B(n_149),
.Y(n_2914)
);

INVx1_ASAP7_75t_SL g2915 ( 
.A(n_2474),
.Y(n_2915)
);

INVx4_ASAP7_75t_L g2916 ( 
.A(n_2272),
.Y(n_2916)
);

INVx3_ASAP7_75t_L g2917 ( 
.A(n_2197),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2164),
.B(n_149),
.Y(n_2918)
);

AOI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2281),
.A2(n_150),
.B(n_151),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2281),
.A2(n_151),
.B(n_152),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2281),
.A2(n_151),
.B(n_152),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2164),
.Y(n_2922)
);

CKINVDCx10_ASAP7_75t_R g2923 ( 
.A(n_2165),
.Y(n_2923)
);

AND2x2_ASAP7_75t_L g2924 ( 
.A(n_2257),
.B(n_153),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2257),
.B(n_153),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2164),
.Y(n_2926)
);

OAI21xp33_ASAP7_75t_L g2927 ( 
.A1(n_2257),
.A2(n_153),
.B(n_154),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2164),
.Y(n_2928)
);

INVx3_ASAP7_75t_L g2929 ( 
.A(n_2197),
.Y(n_2929)
);

OAI21xp5_ASAP7_75t_L g2930 ( 
.A1(n_2281),
.A2(n_154),
.B(n_155),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_SL g2931 ( 
.A(n_2163),
.B(n_155),
.Y(n_2931)
);

AOI22xp5_ASAP7_75t_L g2932 ( 
.A1(n_2500),
.A2(n_157),
.B1(n_154),
.B2(n_156),
.Y(n_2932)
);

INVxp67_ASAP7_75t_SL g2933 ( 
.A(n_2229),
.Y(n_2933)
);

AOI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_2281),
.A2(n_156),
.B(n_158),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2164),
.B(n_156),
.Y(n_2935)
);

CKINVDCx10_ASAP7_75t_R g2936 ( 
.A(n_2165),
.Y(n_2936)
);

BUFx4f_ASAP7_75t_L g2937 ( 
.A(n_2372),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_L g2938 ( 
.A(n_2198),
.B(n_158),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2164),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2164),
.B(n_159),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2281),
.A2(n_159),
.B(n_160),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_2372),
.Y(n_2942)
);

AOI21xp5_ASAP7_75t_L g2943 ( 
.A1(n_2281),
.A2(n_160),
.B(n_161),
.Y(n_2943)
);

A2O1A1Ixp33_ASAP7_75t_L g2944 ( 
.A1(n_2245),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_SL g2945 ( 
.A(n_2163),
.B(n_163),
.Y(n_2945)
);

NOR2xp33_ASAP7_75t_L g2946 ( 
.A(n_2198),
.B(n_162),
.Y(n_2946)
);

OAI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2221),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_2947)
);

O2A1O1Ixp5_ASAP7_75t_L g2948 ( 
.A1(n_2494),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_2948)
);

AOI21xp5_ASAP7_75t_L g2949 ( 
.A1(n_2281),
.A2(n_164),
.B(n_165),
.Y(n_2949)
);

AOI21x1_ASAP7_75t_L g2950 ( 
.A1(n_2263),
.A2(n_166),
.B(n_167),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_SL g2951 ( 
.A(n_2163),
.B(n_167),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2164),
.Y(n_2952)
);

AOI21x1_ASAP7_75t_L g2953 ( 
.A1(n_2263),
.A2(n_166),
.B(n_168),
.Y(n_2953)
);

AOI21xp5_ASAP7_75t_L g2954 ( 
.A1(n_2281),
.A2(n_168),
.B(n_169),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_2163),
.B(n_170),
.Y(n_2955)
);

INVxp67_ASAP7_75t_L g2956 ( 
.A(n_2474),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2164),
.Y(n_2957)
);

OAI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2281),
.A2(n_169),
.B(n_170),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2164),
.B(n_169),
.Y(n_2959)
);

OR2x2_ASAP7_75t_L g2960 ( 
.A(n_2474),
.B(n_170),
.Y(n_2960)
);

AOI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2281),
.A2(n_171),
.B(n_172),
.Y(n_2961)
);

AOI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2281),
.A2(n_171),
.B(n_172),
.Y(n_2962)
);

AOI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2281),
.A2(n_171),
.B(n_172),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2164),
.Y(n_2964)
);

OAI21xp5_ASAP7_75t_L g2965 ( 
.A1(n_2281),
.A2(n_173),
.B(n_174),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2164),
.B(n_173),
.Y(n_2966)
);

AOI21x1_ASAP7_75t_L g2967 ( 
.A1(n_2263),
.A2(n_174),
.B(n_175),
.Y(n_2967)
);

AOI21xp5_ASAP7_75t_L g2968 ( 
.A1(n_2281),
.A2(n_174),
.B(n_175),
.Y(n_2968)
);

AOI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2281),
.A2(n_175),
.B(n_176),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2164),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2164),
.B(n_176),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2257),
.B(n_176),
.Y(n_2972)
);

BUFx4f_ASAP7_75t_L g2973 ( 
.A(n_2372),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2164),
.Y(n_2974)
);

AOI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2500),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_2975)
);

O2A1O1Ixp33_ASAP7_75t_L g2976 ( 
.A1(n_2403),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_L g2977 ( 
.A(n_2198),
.B(n_179),
.Y(n_2977)
);

AOI22xp5_ASAP7_75t_L g2978 ( 
.A1(n_2500),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_2978)
);

INVx3_ASAP7_75t_L g2979 ( 
.A(n_2197),
.Y(n_2979)
);

NOR2xp33_ASAP7_75t_L g2980 ( 
.A(n_2198),
.B(n_180),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2164),
.B(n_180),
.Y(n_2981)
);

OAI22xp5_ASAP7_75t_L g2982 ( 
.A1(n_2221),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_2982)
);

INVx3_ASAP7_75t_L g2983 ( 
.A(n_2197),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2164),
.B(n_181),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2164),
.B(n_183),
.Y(n_2985)
);

OAI22xp5_ASAP7_75t_L g2986 ( 
.A1(n_2221),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2164),
.B(n_184),
.Y(n_2987)
);

NOR2x1_ASAP7_75t_L g2988 ( 
.A(n_2229),
.B(n_184),
.Y(n_2988)
);

A2O1A1Ixp33_ASAP7_75t_L g2989 ( 
.A1(n_2245),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2989)
);

O2A1O1Ixp33_ASAP7_75t_L g2990 ( 
.A1(n_2403),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2164),
.Y(n_2991)
);

A2O1A1Ixp33_ASAP7_75t_L g2992 ( 
.A1(n_2245),
.A2(n_189),
.B(n_187),
.C(n_188),
.Y(n_2992)
);

OAI21xp5_ASAP7_75t_L g2993 ( 
.A1(n_2281),
.A2(n_188),
.B(n_189),
.Y(n_2993)
);

NOR2xp33_ASAP7_75t_L g2994 ( 
.A(n_2198),
.B(n_188),
.Y(n_2994)
);

AOI21xp5_ASAP7_75t_L g2995 ( 
.A1(n_2281),
.A2(n_189),
.B(n_190),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2164),
.B(n_190),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2164),
.B(n_190),
.Y(n_2997)
);

BUFx12f_ASAP7_75t_L g2998 ( 
.A(n_2372),
.Y(n_2998)
);

AOI21xp5_ASAP7_75t_L g2999 ( 
.A1(n_2281),
.A2(n_191),
.B(n_192),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2164),
.B(n_191),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2164),
.Y(n_3001)
);

CKINVDCx5p33_ASAP7_75t_R g3002 ( 
.A(n_2372),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2164),
.B(n_191),
.Y(n_3003)
);

AOI21xp5_ASAP7_75t_L g3004 ( 
.A1(n_2281),
.A2(n_192),
.B(n_193),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2163),
.B(n_194),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2163),
.B(n_194),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2164),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2164),
.Y(n_3008)
);

AOI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2193),
.A2(n_195),
.B1(n_192),
.B2(n_194),
.Y(n_3009)
);

AOI21x1_ASAP7_75t_L g3010 ( 
.A1(n_2263),
.A2(n_195),
.B(n_196),
.Y(n_3010)
);

NAND2x1p5_ASAP7_75t_L g3011 ( 
.A(n_2474),
.B(n_195),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2164),
.B(n_197),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2164),
.B(n_197),
.Y(n_3013)
);

AOI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2193),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_3014)
);

AOI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2281),
.A2(n_198),
.B(n_199),
.Y(n_3015)
);

OAI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2281),
.A2(n_200),
.B(n_201),
.Y(n_3016)
);

AOI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_2281),
.A2(n_200),
.B(n_201),
.Y(n_3017)
);

INVx3_ASAP7_75t_L g3018 ( 
.A(n_2197),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2164),
.B(n_201),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2164),
.B(n_202),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2281),
.A2(n_203),
.B(n_204),
.Y(n_3021)
);

INVx4_ASAP7_75t_L g3022 ( 
.A(n_2272),
.Y(n_3022)
);

OAI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_2221),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2164),
.B(n_203),
.Y(n_3024)
);

A2O1A1Ixp33_ASAP7_75t_L g3025 ( 
.A1(n_2245),
.A2(n_207),
.B(n_205),
.C(n_206),
.Y(n_3025)
);

AO21x1_ASAP7_75t_L g3026 ( 
.A1(n_2263),
.A2(n_613),
.B(n_611),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2164),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2257),
.B(n_205),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2164),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2164),
.B(n_206),
.Y(n_3030)
);

OAI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_2281),
.A2(n_207),
.B(n_208),
.Y(n_3031)
);

INVxp67_ASAP7_75t_L g3032 ( 
.A(n_2474),
.Y(n_3032)
);

AOI21xp5_ASAP7_75t_L g3033 ( 
.A1(n_2281),
.A2(n_207),
.B(n_208),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_2474),
.B(n_208),
.Y(n_3034)
);

BUFx4f_ASAP7_75t_L g3035 ( 
.A(n_2372),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2164),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2164),
.B(n_209),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_L g3038 ( 
.A(n_2198),
.B(n_209),
.Y(n_3038)
);

O2A1O1Ixp33_ASAP7_75t_L g3039 ( 
.A1(n_2403),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_3039)
);

BUFx4f_ASAP7_75t_L g3040 ( 
.A(n_2372),
.Y(n_3040)
);

AOI21xp5_ASAP7_75t_L g3041 ( 
.A1(n_2281),
.A2(n_210),
.B(n_211),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2164),
.B(n_210),
.Y(n_3042)
);

AOI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2281),
.A2(n_211),
.B(n_212),
.Y(n_3043)
);

AOI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2281),
.A2(n_212),
.B(n_213),
.Y(n_3044)
);

OAI21xp5_ASAP7_75t_L g3045 ( 
.A1(n_2281),
.A2(n_213),
.B(n_214),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2198),
.B(n_213),
.Y(n_3046)
);

OAI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2281),
.A2(n_214),
.B(n_215),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2164),
.B(n_215),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2164),
.B(n_215),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2164),
.B(n_216),
.Y(n_3050)
);

AOI21x1_ASAP7_75t_L g3051 ( 
.A1(n_2263),
.A2(n_216),
.B(n_217),
.Y(n_3051)
);

NAND2xp33_ASAP7_75t_L g3052 ( 
.A(n_2287),
.B(n_219),
.Y(n_3052)
);

BUFx8_ASAP7_75t_L g3053 ( 
.A(n_2372),
.Y(n_3053)
);

NOR2xp67_ASAP7_75t_SL g3054 ( 
.A(n_2372),
.B(n_218),
.Y(n_3054)
);

AND2x4_ASAP7_75t_L g3055 ( 
.A(n_2164),
.B(n_218),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_SL g3056 ( 
.A(n_2163),
.B(n_220),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2164),
.B(n_219),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2164),
.B(n_220),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2164),
.Y(n_3059)
);

O2A1O1Ixp33_ASAP7_75t_L g3060 ( 
.A1(n_2403),
.A2(n_223),
.B(n_221),
.C(n_222),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2164),
.Y(n_3061)
);

AOI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_2281),
.A2(n_223),
.B(n_224),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2164),
.B(n_223),
.Y(n_3063)
);

NOR2xp33_ASAP7_75t_L g3064 ( 
.A(n_2198),
.B(n_224),
.Y(n_3064)
);

AOI21xp5_ASAP7_75t_L g3065 ( 
.A1(n_2281),
.A2(n_224),
.B(n_225),
.Y(n_3065)
);

BUFx6f_ASAP7_75t_L g3066 ( 
.A(n_2287),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_SL g3067 ( 
.A(n_2163),
.B(n_226),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_2163),
.B(n_227),
.Y(n_3068)
);

NOR2xp33_ASAP7_75t_L g3069 ( 
.A(n_2198),
.B(n_225),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2164),
.Y(n_3070)
);

AOI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2281),
.A2(n_225),
.B(n_227),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2164),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2164),
.B(n_228),
.Y(n_3073)
);

BUFx3_ASAP7_75t_L g3074 ( 
.A(n_2229),
.Y(n_3074)
);

INVx4_ASAP7_75t_L g3075 ( 
.A(n_2272),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2163),
.B(n_229),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_SL g3077 ( 
.A(n_2163),
.B(n_230),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2164),
.B(n_228),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2164),
.B(n_228),
.Y(n_3079)
);

HB1xp67_ASAP7_75t_L g3080 ( 
.A(n_2474),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2164),
.B(n_231),
.Y(n_3081)
);

NOR2xp33_ASAP7_75t_L g3082 ( 
.A(n_2198),
.B(n_231),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2281),
.A2(n_232),
.B(n_233),
.Y(n_3083)
);

BUFx2_ASAP7_75t_L g3084 ( 
.A(n_2229),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2281),
.A2(n_232),
.B(n_233),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2164),
.Y(n_3086)
);

BUFx8_ASAP7_75t_L g3087 ( 
.A(n_2372),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_SL g3088 ( 
.A(n_2163),
.B(n_235),
.Y(n_3088)
);

OAI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_2281),
.A2(n_234),
.B(n_235),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2164),
.Y(n_3090)
);

AOI21x1_ASAP7_75t_L g3091 ( 
.A1(n_2263),
.A2(n_234),
.B(n_235),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2164),
.Y(n_3092)
);

BUFx2_ASAP7_75t_L g3093 ( 
.A(n_2229),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2164),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2164),
.B(n_236),
.Y(n_3095)
);

OAI21xp5_ASAP7_75t_L g3096 ( 
.A1(n_2281),
.A2(n_236),
.B(n_237),
.Y(n_3096)
);

AOI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_2257),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_2198),
.B(n_238),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_SL g3099 ( 
.A(n_2163),
.B(n_239),
.Y(n_3099)
);

AOI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2281),
.A2(n_238),
.B(n_239),
.Y(n_3100)
);

AOI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_2281),
.A2(n_240),
.B(n_241),
.Y(n_3101)
);

AND2x6_ASAP7_75t_L g3102 ( 
.A(n_2164),
.B(n_240),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2164),
.B(n_240),
.Y(n_3103)
);

NOR2xp33_ASAP7_75t_L g3104 ( 
.A(n_2198),
.B(n_241),
.Y(n_3104)
);

NOR2xp33_ASAP7_75t_L g3105 ( 
.A(n_2198),
.B(n_242),
.Y(n_3105)
);

BUFx6f_ASAP7_75t_L g3106 ( 
.A(n_2287),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_2281),
.A2(n_242),
.B(n_243),
.Y(n_3107)
);

AOI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_2281),
.A2(n_242),
.B(n_243),
.Y(n_3108)
);

OAI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2281),
.A2(n_243),
.B(n_244),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2257),
.B(n_244),
.Y(n_3110)
);

NOR2xp33_ASAP7_75t_L g3111 ( 
.A(n_2198),
.B(n_245),
.Y(n_3111)
);

A2O1A1Ixp33_ASAP7_75t_L g3112 ( 
.A1(n_2245),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_2197),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2164),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2281),
.A2(n_246),
.B(n_247),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2164),
.Y(n_3116)
);

AOI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2281),
.A2(n_247),
.B(n_248),
.Y(n_3117)
);

A2O1A1Ixp33_ASAP7_75t_L g3118 ( 
.A1(n_2245),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_SL g3119 ( 
.A(n_2163),
.B(n_249),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_2198),
.B(n_248),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2164),
.B(n_249),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2287),
.Y(n_3122)
);

OR2x2_ASAP7_75t_L g3123 ( 
.A(n_2474),
.B(n_250),
.Y(n_3123)
);

AOI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2281),
.A2(n_251),
.B(n_252),
.Y(n_3124)
);

AOI21xp5_ASAP7_75t_L g3125 ( 
.A1(n_2281),
.A2(n_251),
.B(n_252),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2164),
.B(n_252),
.Y(n_3126)
);

AOI21xp5_ASAP7_75t_L g3127 ( 
.A1(n_2281),
.A2(n_253),
.B(n_254),
.Y(n_3127)
);

INVx4_ASAP7_75t_L g3128 ( 
.A(n_2272),
.Y(n_3128)
);

AOI21x1_ASAP7_75t_L g3129 ( 
.A1(n_2263),
.A2(n_253),
.B(n_254),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2164),
.Y(n_3130)
);

AOI21xp5_ASAP7_75t_L g3131 ( 
.A1(n_2281),
.A2(n_254),
.B(n_255),
.Y(n_3131)
);

HB1xp67_ASAP7_75t_L g3132 ( 
.A(n_2474),
.Y(n_3132)
);

AOI21xp5_ASAP7_75t_L g3133 ( 
.A1(n_2281),
.A2(n_256),
.B(n_257),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2164),
.B(n_257),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2164),
.B(n_258),
.Y(n_3135)
);

AND2x4_ASAP7_75t_L g3136 ( 
.A(n_2164),
.B(n_259),
.Y(n_3136)
);

O2A1O1Ixp33_ASAP7_75t_L g3137 ( 
.A1(n_2403),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_3137)
);

AOI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_2281),
.A2(n_260),
.B(n_261),
.Y(n_3138)
);

OAI21xp33_ASAP7_75t_L g3139 ( 
.A1(n_2257),
.A2(n_262),
.B(n_263),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2164),
.B(n_262),
.Y(n_3140)
);

AOI21xp5_ASAP7_75t_L g3141 ( 
.A1(n_2281),
.A2(n_262),
.B(n_263),
.Y(n_3141)
);

AOI21xp5_ASAP7_75t_L g3142 ( 
.A1(n_2281),
.A2(n_264),
.B(n_265),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2164),
.B(n_264),
.Y(n_3143)
);

NOR2xp67_ASAP7_75t_L g3144 ( 
.A(n_2372),
.B(n_264),
.Y(n_3144)
);

INVx2_ASAP7_75t_SL g3145 ( 
.A(n_2474),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2257),
.B(n_265),
.Y(n_3146)
);

AOI21xp5_ASAP7_75t_L g3147 ( 
.A1(n_2281),
.A2(n_265),
.B(n_266),
.Y(n_3147)
);

O2A1O1Ixp33_ASAP7_75t_L g3148 ( 
.A1(n_2403),
.A2(n_268),
.B(n_266),
.C(n_267),
.Y(n_3148)
);

OAI21xp5_ASAP7_75t_L g3149 ( 
.A1(n_2281),
.A2(n_266),
.B(n_267),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2164),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2164),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2164),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_SL g3153 ( 
.A(n_2163),
.B(n_269),
.Y(n_3153)
);

INVx4_ASAP7_75t_L g3154 ( 
.A(n_2272),
.Y(n_3154)
);

AOI21xp5_ASAP7_75t_L g3155 ( 
.A1(n_2281),
.A2(n_268),
.B(n_269),
.Y(n_3155)
);

NOR3xp33_ASAP7_75t_SL g3156 ( 
.A(n_2942),
.B(n_270),
.C(n_271),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2900),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2566),
.A2(n_2534),
.B(n_2698),
.Y(n_3158)
);

A2O1A1Ixp33_ASAP7_75t_L g3159 ( 
.A1(n_2899),
.A2(n_272),
.B(n_270),
.C(n_271),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2575),
.Y(n_3160)
);

NOR2xp67_ASAP7_75t_L g3161 ( 
.A(n_2675),
.B(n_270),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2901),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2715),
.A2(n_2778),
.B(n_2806),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2912),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2725),
.B(n_2911),
.Y(n_3165)
);

AOI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_2544),
.A2(n_272),
.B(n_273),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_SL g3167 ( 
.A(n_2725),
.B(n_613),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2922),
.Y(n_3168)
);

CKINVDCx5p33_ASAP7_75t_R g3169 ( 
.A(n_3053),
.Y(n_3169)
);

OAI22xp5_ASAP7_75t_L g3170 ( 
.A1(n_2641),
.A2(n_275),
.B1(n_272),
.B2(n_274),
.Y(n_3170)
);

CKINVDCx5p33_ASAP7_75t_R g3171 ( 
.A(n_3053),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_SL g3172 ( 
.A(n_2915),
.B(n_614),
.Y(n_3172)
);

O2A1O1Ixp5_ASAP7_75t_L g3173 ( 
.A1(n_2589),
.A2(n_277),
.B(n_274),
.C(n_276),
.Y(n_3173)
);

AOI21xp5_ASAP7_75t_L g3174 ( 
.A1(n_2552),
.A2(n_276),
.B(n_277),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2688),
.B(n_276),
.Y(n_3175)
);

BUFx3_ASAP7_75t_L g3176 ( 
.A(n_2601),
.Y(n_3176)
);

OAI22xp5_ASAP7_75t_L g3177 ( 
.A1(n_2589),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_3177)
);

AOI22xp33_ASAP7_75t_L g3178 ( 
.A1(n_3102),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_3178)
);

BUFx12f_ASAP7_75t_L g3179 ( 
.A(n_3087),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_R g3180 ( 
.A(n_2923),
.B(n_278),
.Y(n_3180)
);

NOR2xp33_ASAP7_75t_R g3181 ( 
.A(n_2923),
.B(n_279),
.Y(n_3181)
);

AO21x2_ASAP7_75t_L g3182 ( 
.A1(n_2913),
.A2(n_281),
.B(n_282),
.Y(n_3182)
);

AND2x4_ASAP7_75t_L g3183 ( 
.A(n_2675),
.B(n_281),
.Y(n_3183)
);

AOI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_2582),
.A2(n_281),
.B(n_282),
.Y(n_3184)
);

AOI22xp5_ASAP7_75t_L g3185 ( 
.A1(n_2559),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_3185)
);

CKINVDCx5p33_ASAP7_75t_R g3186 ( 
.A(n_3087),
.Y(n_3186)
);

A2O1A1Ixp33_ASAP7_75t_L g3187 ( 
.A1(n_2930),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_3187)
);

OAI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_2883),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_3188)
);

AND2x4_ASAP7_75t_L g3189 ( 
.A(n_2801),
.B(n_286),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_2737),
.A2(n_2596),
.B(n_2765),
.Y(n_3190)
);

NOR3xp33_ASAP7_75t_SL g3191 ( 
.A(n_3002),
.B(n_2744),
.C(n_2667),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_SL g3192 ( 
.A(n_2543),
.B(n_614),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_2567),
.A2(n_286),
.B(n_287),
.Y(n_3193)
);

AND2x4_ASAP7_75t_L g3194 ( 
.A(n_2801),
.B(n_286),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_SL g3195 ( 
.A(n_2956),
.B(n_615),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_2614),
.B(n_287),
.Y(n_3196)
);

INVx5_ASAP7_75t_L g3197 ( 
.A(n_2601),
.Y(n_3197)
);

INVx5_ASAP7_75t_L g3198 ( 
.A(n_2601),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_SL g3199 ( 
.A(n_3032),
.B(n_615),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2556),
.Y(n_3200)
);

OAI21xp33_ASAP7_75t_SL g3201 ( 
.A1(n_2883),
.A2(n_288),
.B(n_289),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2592),
.B(n_288),
.Y(n_3202)
);

AOI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_2573),
.A2(n_288),
.B(n_289),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_SL g3204 ( 
.A(n_3145),
.B(n_2802),
.Y(n_3204)
);

INVx5_ASAP7_75t_L g3205 ( 
.A(n_2746),
.Y(n_3205)
);

A2O1A1Ixp33_ASAP7_75t_SL g3206 ( 
.A1(n_2833),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_3206)
);

NOR3xp33_ASAP7_75t_SL g3207 ( 
.A(n_2896),
.B(n_290),
.C(n_291),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2565),
.Y(n_3208)
);

OAI22xp5_ASAP7_75t_SL g3209 ( 
.A1(n_2717),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2576),
.A2(n_292),
.B(n_294),
.Y(n_3210)
);

O2A1O1Ixp5_ASAP7_75t_L g3211 ( 
.A1(n_2577),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_3211)
);

NOR2xp33_ASAP7_75t_L g3212 ( 
.A(n_2828),
.B(n_295),
.Y(n_3212)
);

OAI21x1_ASAP7_75t_L g3213 ( 
.A1(n_2870),
.A2(n_295),
.B(n_297),
.Y(n_3213)
);

NOR2xp33_ASAP7_75t_L g3214 ( 
.A(n_2760),
.B(n_2777),
.Y(n_3214)
);

AOI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_2586),
.A2(n_297),
.B(n_298),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2568),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_2818),
.A2(n_299),
.B(n_300),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2926),
.Y(n_3218)
);

CKINVDCx5p33_ASAP7_75t_R g3219 ( 
.A(n_2998),
.Y(n_3219)
);

BUFx6f_ASAP7_75t_SL g3220 ( 
.A(n_2602),
.Y(n_3220)
);

OAI22xp5_ASAP7_75t_L g3221 ( 
.A1(n_2932),
.A2(n_2978),
.B1(n_2975),
.B2(n_3055),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_2548),
.A2(n_2843),
.B(n_2590),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2579),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2587),
.Y(n_3224)
);

INVx8_ASAP7_75t_L g3225 ( 
.A(n_2746),
.Y(n_3225)
);

OAI22xp5_ASAP7_75t_L g3226 ( 
.A1(n_2932),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3055),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3136),
.Y(n_3228)
);

OAI22xp5_ASAP7_75t_L g3229 ( 
.A1(n_2975),
.A2(n_302),
.B1(n_299),
.B2(n_301),
.Y(n_3229)
);

AOI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_2647),
.A2(n_301),
.B(n_302),
.Y(n_3230)
);

AND2x4_ASAP7_75t_L g3231 ( 
.A(n_2570),
.B(n_302),
.Y(n_3231)
);

BUFx12f_ASAP7_75t_L g3232 ( 
.A(n_2858),
.Y(n_3232)
);

AND2x4_ASAP7_75t_L g3233 ( 
.A(n_2570),
.B(n_303),
.Y(n_3233)
);

OAI21x1_ASAP7_75t_L g3234 ( 
.A1(n_2870),
.A2(n_303),
.B(n_304),
.Y(n_3234)
);

INVxp67_ASAP7_75t_SL g3235 ( 
.A(n_3080),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_R g3236 ( 
.A(n_2936),
.B(n_304),
.Y(n_3236)
);

OAI22xp5_ASAP7_75t_SL g3237 ( 
.A1(n_2752),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_2964),
.Y(n_3238)
);

A2O1A1Ixp33_ASAP7_75t_L g3239 ( 
.A1(n_2958),
.A2(n_308),
.B(n_305),
.C(n_307),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2841),
.B(n_308),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_2654),
.A2(n_308),
.B(n_309),
.Y(n_3241)
);

CKINVDCx14_ASAP7_75t_R g3242 ( 
.A(n_2904),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_2732),
.B(n_309),
.Y(n_3243)
);

OR2x6_ASAP7_75t_SL g3244 ( 
.A(n_2936),
.B(n_310),
.Y(n_3244)
);

OAI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_2978),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_3245)
);

AOI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_2661),
.A2(n_310),
.B(n_311),
.Y(n_3246)
);

INVxp67_ASAP7_75t_L g3247 ( 
.A(n_3132),
.Y(n_3247)
);

CKINVDCx20_ASAP7_75t_R g3248 ( 
.A(n_2904),
.Y(n_3248)
);

AOI22xp33_ASAP7_75t_SL g3249 ( 
.A1(n_2789),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_3249)
);

AOI21xp5_ASAP7_75t_L g3250 ( 
.A1(n_2671),
.A2(n_313),
.B(n_314),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_L g3251 ( 
.A(n_2734),
.B(n_313),
.Y(n_3251)
);

CKINVDCx5p33_ASAP7_75t_R g3252 ( 
.A(n_2937),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3136),
.Y(n_3253)
);

HB1xp67_ASAP7_75t_L g3254 ( 
.A(n_2619),
.Y(n_3254)
);

BUFx2_ASAP7_75t_L g3255 ( 
.A(n_2539),
.Y(n_3255)
);

BUFx3_ASAP7_75t_L g3256 ( 
.A(n_2937),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2594),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2890),
.B(n_314),
.Y(n_3258)
);

BUFx12f_ASAP7_75t_L g3259 ( 
.A(n_2858),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_2974),
.Y(n_3260)
);

AOI221xp5_ASAP7_75t_L g3261 ( 
.A1(n_2722),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.C(n_319),
.Y(n_3261)
);

O2A1O1Ixp33_ASAP7_75t_L g3262 ( 
.A1(n_2735),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_3262)
);

O2A1O1Ixp33_ASAP7_75t_L g3263 ( 
.A1(n_2644),
.A2(n_320),
.B(n_318),
.C(n_319),
.Y(n_3263)
);

AOI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_2551),
.A2(n_2593),
.B(n_2563),
.Y(n_3264)
);

AOI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_2560),
.A2(n_319),
.B(n_320),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2924),
.B(n_2925),
.Y(n_3266)
);

CKINVDCx5p33_ASAP7_75t_R g3267 ( 
.A(n_2973),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2646),
.Y(n_3268)
);

HB1xp67_ASAP7_75t_L g3269 ( 
.A(n_3074),
.Y(n_3269)
);

NAND3xp33_ASAP7_75t_L g3270 ( 
.A(n_2580),
.B(n_321),
.C(n_322),
.Y(n_3270)
);

BUFx6f_ASAP7_75t_L g3271 ( 
.A(n_2591),
.Y(n_3271)
);

AOI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_2564),
.A2(n_321),
.B(n_322),
.Y(n_3272)
);

BUFx6f_ASAP7_75t_L g3273 ( 
.A(n_2591),
.Y(n_3273)
);

INVx2_ASAP7_75t_L g3274 ( 
.A(n_3007),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_SL g3275 ( 
.A(n_2599),
.B(n_616),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_2972),
.B(n_321),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_3028),
.B(n_3110),
.Y(n_3277)
);

CKINVDCx20_ASAP7_75t_R g3278 ( 
.A(n_2973),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2631),
.Y(n_3279)
);

OAI21xp33_ASAP7_75t_SL g3280 ( 
.A1(n_2754),
.A2(n_323),
.B(n_324),
.Y(n_3280)
);

HB1xp67_ASAP7_75t_L g3281 ( 
.A(n_3084),
.Y(n_3281)
);

AOI21x1_ASAP7_75t_L g3282 ( 
.A1(n_2731),
.A2(n_323),
.B(n_324),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2642),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_2569),
.A2(n_2574),
.B(n_2572),
.Y(n_3284)
);

AOI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_2845),
.A2(n_324),
.B(n_325),
.Y(n_3285)
);

INVx3_ASAP7_75t_L g3286 ( 
.A(n_2712),
.Y(n_3286)
);

HB1xp67_ASAP7_75t_L g3287 ( 
.A(n_3093),
.Y(n_3287)
);

BUFx6f_ASAP7_75t_L g3288 ( 
.A(n_2591),
.Y(n_3288)
);

OAI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_2754),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_3289)
);

O2A1O1Ixp33_ASAP7_75t_L g3290 ( 
.A1(n_2768),
.A2(n_328),
.B(n_326),
.C(n_327),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2650),
.Y(n_3291)
);

HB1xp67_ASAP7_75t_L g3292 ( 
.A(n_2638),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_SL g3293 ( 
.A(n_2599),
.B(n_616),
.Y(n_3293)
);

AND2x2_ASAP7_75t_L g3294 ( 
.A(n_3146),
.B(n_327),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2536),
.Y(n_3295)
);

AOI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_2686),
.A2(n_328),
.B(n_329),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3008),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2537),
.Y(n_3298)
);

INVxp67_ASAP7_75t_L g3299 ( 
.A(n_2620),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_3036),
.Y(n_3300)
);

OAI22xp5_ASAP7_75t_L g3301 ( 
.A1(n_2730),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_3301)
);

INVx3_ASAP7_75t_L g3302 ( 
.A(n_2712),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2885),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2905),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_2928),
.B(n_330),
.Y(n_3305)
);

A2O1A1Ixp33_ASAP7_75t_SL g3306 ( 
.A1(n_2837),
.A2(n_2993),
.B(n_3016),
.C(n_2965),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2939),
.Y(n_3307)
);

O2A1O1Ixp33_ASAP7_75t_L g3308 ( 
.A1(n_2705),
.A2(n_332),
.B(n_330),
.C(n_331),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_SL g3309 ( 
.A(n_2561),
.B(n_2798),
.Y(n_3309)
);

HB1xp67_ASAP7_75t_L g3310 ( 
.A(n_2820),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_SL g3311 ( 
.A(n_2909),
.B(n_618),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_3059),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_2952),
.B(n_331),
.Y(n_3313)
);

OAI22xp5_ASAP7_75t_L g3314 ( 
.A1(n_2730),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3061),
.Y(n_3315)
);

OAI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_2840),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_3316)
);

AOI21xp5_ASAP7_75t_L g3317 ( 
.A1(n_2553),
.A2(n_333),
.B(n_335),
.Y(n_3317)
);

BUFx2_ASAP7_75t_L g3318 ( 
.A(n_2933),
.Y(n_3318)
);

CKINVDCx20_ASAP7_75t_R g3319 ( 
.A(n_3035),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2957),
.Y(n_3320)
);

BUFx3_ASAP7_75t_L g3321 ( 
.A(n_3035),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_2840),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_3322)
);

CKINVDCx5p33_ASAP7_75t_R g3323 ( 
.A(n_3040),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_2970),
.B(n_337),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2991),
.B(n_3001),
.Y(n_3325)
);

AND2x4_ASAP7_75t_L g3326 ( 
.A(n_2584),
.B(n_337),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3027),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3029),
.Y(n_3328)
);

OAI22xp5_ASAP7_75t_L g3329 ( 
.A1(n_2562),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3072),
.B(n_338),
.Y(n_3330)
);

O2A1O1Ixp33_ASAP7_75t_L g3331 ( 
.A1(n_2687),
.A2(n_340),
.B(n_338),
.C(n_339),
.Y(n_3331)
);

AND2x4_ASAP7_75t_L g3332 ( 
.A(n_2584),
.B(n_339),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_SL g3333 ( 
.A(n_3011),
.B(n_622),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3090),
.B(n_340),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3092),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_2555),
.A2(n_341),
.B(n_342),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3114),
.B(n_341),
.Y(n_3337)
);

OR2x6_ASAP7_75t_L g3338 ( 
.A(n_2916),
.B(n_341),
.Y(n_3338)
);

NOR2xp67_ASAP7_75t_L g3339 ( 
.A(n_2916),
.B(n_343),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3130),
.Y(n_3340)
);

BUFx2_ASAP7_75t_L g3341 ( 
.A(n_2746),
.Y(n_3341)
);

AOI21xp5_ASAP7_75t_L g3342 ( 
.A1(n_2557),
.A2(n_343),
.B(n_344),
.Y(n_3342)
);

AOI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_2549),
.A2(n_343),
.B(n_344),
.Y(n_3343)
);

NAND3xp33_ASAP7_75t_L g3344 ( 
.A(n_2774),
.B(n_345),
.C(n_346),
.Y(n_3344)
);

INVx4_ASAP7_75t_L g3345 ( 
.A(n_3040),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3070),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3151),
.Y(n_3347)
);

BUFx2_ASAP7_75t_L g3348 ( 
.A(n_2746),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3152),
.Y(n_3349)
);

BUFx6f_ASAP7_75t_L g3350 ( 
.A(n_2657),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2540),
.B(n_345),
.Y(n_3351)
);

NOR2xp33_ASAP7_75t_L g3352 ( 
.A(n_2738),
.B(n_345),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_SL g3353 ( 
.A(n_2820),
.B(n_622),
.Y(n_3353)
);

OAI22x1_ASAP7_75t_L g3354 ( 
.A1(n_2724),
.A2(n_2988),
.B1(n_3014),
.B2(n_3009),
.Y(n_3354)
);

OAI22xp5_ASAP7_75t_L g3355 ( 
.A1(n_2629),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_3355)
);

AND2x4_ASAP7_75t_L g3356 ( 
.A(n_3022),
.B(n_346),
.Y(n_3356)
);

INVxp67_ASAP7_75t_L g3357 ( 
.A(n_3102),
.Y(n_3357)
);

AOI21xp5_ASAP7_75t_L g3358 ( 
.A1(n_2632),
.A2(n_347),
.B(n_348),
.Y(n_3358)
);

AOI22xp5_ASAP7_75t_L g3359 ( 
.A1(n_2674),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_3359)
);

AOI21xp5_ASAP7_75t_L g3360 ( 
.A1(n_2634),
.A2(n_349),
.B(n_351),
.Y(n_3360)
);

O2A1O1Ixp33_ASAP7_75t_L g3361 ( 
.A1(n_2607),
.A2(n_352),
.B(n_349),
.C(n_351),
.Y(n_3361)
);

OAI21xp5_ASAP7_75t_L g3362 ( 
.A1(n_2640),
.A2(n_352),
.B(n_353),
.Y(n_3362)
);

BUFx6f_ASAP7_75t_L g3363 ( 
.A(n_2657),
.Y(n_3363)
);

A2O1A1Ixp33_ASAP7_75t_L g3364 ( 
.A1(n_3031),
.A2(n_356),
.B(n_354),
.C(n_355),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_3086),
.Y(n_3365)
);

NOR3xp33_ASAP7_75t_L g3366 ( 
.A(n_2609),
.B(n_354),
.C(n_355),
.Y(n_3366)
);

OAI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_2643),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_3367)
);

AOI21xp5_ASAP7_75t_L g3368 ( 
.A1(n_2878),
.A2(n_357),
.B(n_358),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_SL g3369 ( 
.A(n_2712),
.B(n_623),
.Y(n_3369)
);

OAI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_2627),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_3370)
);

HB1xp67_ASAP7_75t_L g3371 ( 
.A(n_2660),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_SL g3372 ( 
.A(n_2740),
.B(n_624),
.Y(n_3372)
);

OAI22xp5_ASAP7_75t_L g3373 ( 
.A1(n_2621),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3094),
.B(n_360),
.Y(n_3374)
);

AOI22xp5_ASAP7_75t_L g3375 ( 
.A1(n_3102),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_L g3376 ( 
.A(n_2706),
.B(n_361),
.Y(n_3376)
);

AOI21xp5_ASAP7_75t_L g3377 ( 
.A1(n_2879),
.A2(n_362),
.B(n_363),
.Y(n_3377)
);

INVx4_ASAP7_75t_L g3378 ( 
.A(n_3022),
.Y(n_3378)
);

BUFx6f_ASAP7_75t_L g3379 ( 
.A(n_2657),
.Y(n_3379)
);

AOI21xp5_ASAP7_75t_L g3380 ( 
.A1(n_2891),
.A2(n_362),
.B(n_363),
.Y(n_3380)
);

AOI22x1_ASAP7_75t_L g3381 ( 
.A1(n_2598),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_3381)
);

INVx3_ASAP7_75t_L g3382 ( 
.A(n_2740),
.Y(n_3382)
);

HB1xp67_ASAP7_75t_L g3383 ( 
.A(n_2583),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2665),
.Y(n_3384)
);

A2O1A1Ixp33_ASAP7_75t_L g3385 ( 
.A1(n_3045),
.A2(n_366),
.B(n_364),
.C(n_365),
.Y(n_3385)
);

AOI221xp5_ASAP7_75t_L g3386 ( 
.A1(n_2881),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.C(n_367),
.Y(n_3386)
);

NOR2xp33_ASAP7_75t_L g3387 ( 
.A(n_2836),
.B(n_367),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_2678),
.Y(n_3388)
);

AND2x4_ASAP7_75t_L g3389 ( 
.A(n_3075),
.B(n_368),
.Y(n_3389)
);

NAND2xp33_ASAP7_75t_R g3390 ( 
.A(n_2827),
.B(n_368),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_SL g3391 ( 
.A(n_2740),
.B(n_624),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3116),
.B(n_368),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3150),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_2663),
.B(n_369),
.Y(n_3394)
);

AND2x2_ASAP7_75t_L g3395 ( 
.A(n_2782),
.B(n_369),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_2871),
.B(n_370),
.Y(n_3396)
);

OR2x2_ASAP7_75t_L g3397 ( 
.A(n_2585),
.B(n_370),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_2681),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_2690),
.Y(n_3399)
);

INVx3_ASAP7_75t_L g3400 ( 
.A(n_2910),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_2691),
.B(n_371),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_2711),
.B(n_372),
.Y(n_3402)
);

INVxp67_ASAP7_75t_SL g3403 ( 
.A(n_2910),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_2788),
.B(n_2664),
.Y(n_3404)
);

BUFx6f_ASAP7_75t_L g3405 ( 
.A(n_2910),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_2815),
.B(n_372),
.Y(n_3406)
);

CKINVDCx20_ASAP7_75t_R g3407 ( 
.A(n_3075),
.Y(n_3407)
);

O2A1O1Ixp33_ASAP7_75t_L g3408 ( 
.A1(n_2838),
.A2(n_374),
.B(n_372),
.C(n_373),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_2694),
.B(n_373),
.Y(n_3409)
);

NAND2xp33_ASAP7_75t_L g3410 ( 
.A(n_3066),
.B(n_3106),
.Y(n_3410)
);

INVxp67_ASAP7_75t_L g3411 ( 
.A(n_3102),
.Y(n_3411)
);

BUFx6f_ASAP7_75t_L g3412 ( 
.A(n_3066),
.Y(n_3412)
);

HB1xp67_ASAP7_75t_L g3413 ( 
.A(n_2824),
.Y(n_3413)
);

A2O1A1Ixp33_ASAP7_75t_SL g3414 ( 
.A1(n_3047),
.A2(n_376),
.B(n_373),
.C(n_375),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_2775),
.B(n_2784),
.Y(n_3415)
);

AOI21xp5_ASAP7_75t_L g3416 ( 
.A1(n_2895),
.A2(n_375),
.B(n_376),
.Y(n_3416)
);

A2O1A1Ixp33_ASAP7_75t_SL g3417 ( 
.A1(n_3089),
.A2(n_378),
.B(n_376),
.C(n_377),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_2689),
.B(n_377),
.Y(n_3418)
);

AOI21xp5_ASAP7_75t_L g3419 ( 
.A1(n_2906),
.A2(n_377),
.B(n_378),
.Y(n_3419)
);

BUFx8_ASAP7_75t_SL g3420 ( 
.A(n_2753),
.Y(n_3420)
);

OAI21x1_ASAP7_75t_L g3421 ( 
.A1(n_2892),
.A2(n_378),
.B(n_379),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_3066),
.B(n_625),
.Y(n_3422)
);

INVx3_ASAP7_75t_L g3423 ( 
.A(n_3106),
.Y(n_3423)
);

INVx4_ASAP7_75t_L g3424 ( 
.A(n_3128),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_2658),
.B(n_379),
.Y(n_3425)
);

AND2x2_ASAP7_75t_SL g3426 ( 
.A(n_2797),
.B(n_380),
.Y(n_3426)
);

AOI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_2907),
.A2(n_380),
.B(n_381),
.Y(n_3427)
);

NOR2xp33_ASAP7_75t_L g3428 ( 
.A(n_2673),
.B(n_381),
.Y(n_3428)
);

BUFx4f_ASAP7_75t_L g3429 ( 
.A(n_2606),
.Y(n_3429)
);

NOR2x1_ASAP7_75t_SL g3430 ( 
.A(n_3106),
.B(n_381),
.Y(n_3430)
);

O2A1O1Ixp5_ASAP7_75t_L g3431 ( 
.A1(n_3096),
.A2(n_384),
.B(n_382),
.C(n_383),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_R g3432 ( 
.A(n_3128),
.B(n_383),
.Y(n_3432)
);

OAI21x1_ASAP7_75t_SL g3433 ( 
.A1(n_3109),
.A2(n_3149),
.B(n_2622),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_2919),
.A2(n_383),
.B(n_385),
.Y(n_3434)
);

A2O1A1Ixp33_ASAP7_75t_L g3435 ( 
.A1(n_3155),
.A2(n_387),
.B(n_385),
.C(n_386),
.Y(n_3435)
);

BUFx6f_ASAP7_75t_L g3436 ( 
.A(n_3122),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_2887),
.B(n_385),
.Y(n_3437)
);

A2O1A1Ixp33_ASAP7_75t_L g3438 ( 
.A1(n_2920),
.A2(n_388),
.B(n_386),
.C(n_387),
.Y(n_3438)
);

OAI22x1_ASAP7_75t_L g3439 ( 
.A1(n_2710),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_2880),
.Y(n_3440)
);

A2O1A1Ixp33_ASAP7_75t_L g3441 ( 
.A1(n_2921),
.A2(n_390),
.B(n_388),
.C(n_389),
.Y(n_3441)
);

O2A1O1Ixp33_ASAP7_75t_L g3442 ( 
.A1(n_2839),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_3442)
);

AO21x1_ASAP7_75t_L g3443 ( 
.A1(n_2816),
.A2(n_626),
.B(n_625),
.Y(n_3443)
);

XOR2xp5_ASAP7_75t_L g3444 ( 
.A(n_2813),
.B(n_390),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_2898),
.B(n_389),
.Y(n_3445)
);

BUFx4f_ASAP7_75t_SL g3446 ( 
.A(n_3154),
.Y(n_3446)
);

OAI22xp5_ASAP7_75t_L g3447 ( 
.A1(n_2668),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_SL g3448 ( 
.A(n_3122),
.B(n_626),
.Y(n_3448)
);

INVx4_ASAP7_75t_L g3449 ( 
.A(n_3154),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_2934),
.A2(n_391),
.B(n_392),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_2679),
.B(n_2571),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_2897),
.B(n_392),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_2882),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_2824),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_3454)
);

AOI21xp5_ASAP7_75t_L g3455 ( 
.A1(n_2941),
.A2(n_393),
.B(n_394),
.Y(n_3455)
);

INVxp67_ASAP7_75t_SL g3456 ( 
.A(n_3122),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_2886),
.Y(n_3457)
);

OAI221xp5_ASAP7_75t_L g3458 ( 
.A1(n_2736),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.C(n_397),
.Y(n_3458)
);

AOI22xp33_ASAP7_75t_L g3459 ( 
.A1(n_2908),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_3459)
);

BUFx12f_ASAP7_75t_L g3460 ( 
.A(n_2721),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_SL g3461 ( 
.A(n_2610),
.B(n_627),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2888),
.Y(n_3462)
);

A2O1A1Ixp33_ASAP7_75t_L g3463 ( 
.A1(n_2943),
.A2(n_400),
.B(n_398),
.C(n_399),
.Y(n_3463)
);

OAI21x1_ASAP7_75t_L g3464 ( 
.A1(n_2547),
.A2(n_398),
.B(n_399),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_2938),
.B(n_400),
.Y(n_3465)
);

O2A1O1Ixp33_ASAP7_75t_L g3466 ( 
.A1(n_2808),
.A2(n_402),
.B(n_400),
.C(n_401),
.Y(n_3466)
);

CKINVDCx5p33_ASAP7_75t_R g3467 ( 
.A(n_2753),
.Y(n_3467)
);

NOR2xp33_ASAP7_75t_L g3468 ( 
.A(n_2685),
.B(n_401),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_2889),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_2949),
.A2(n_401),
.B(n_402),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_2960),
.B(n_628),
.Y(n_3471)
);

BUFx2_ASAP7_75t_L g3472 ( 
.A(n_2809),
.Y(n_3472)
);

AO21x2_ASAP7_75t_L g3473 ( 
.A1(n_2776),
.A2(n_404),
.B(n_405),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_2954),
.A2(n_404),
.B(n_405),
.Y(n_3474)
);

OR2x4_ASAP7_75t_L g3475 ( 
.A(n_2863),
.B(n_405),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_2714),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_2894),
.Y(n_3477)
);

BUFx12f_ASAP7_75t_L g3478 ( 
.A(n_2721),
.Y(n_3478)
);

AND2x2_ASAP7_75t_SL g3479 ( 
.A(n_2893),
.B(n_406),
.Y(n_3479)
);

INVxp67_ASAP7_75t_SL g3480 ( 
.A(n_3052),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_2767),
.B(n_406),
.Y(n_3481)
);

AO32x1_ASAP7_75t_L g3482 ( 
.A1(n_2739),
.A2(n_408),
.A3(n_406),
.B1(n_407),
.B2(n_409),
.Y(n_3482)
);

OAI22xp5_ASAP7_75t_L g3483 ( 
.A1(n_2826),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_SL g3484 ( 
.A(n_3034),
.B(n_629),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_2914),
.Y(n_3485)
);

OAI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_2807),
.A2(n_407),
.B(n_409),
.Y(n_3486)
);

AND2x4_ASAP7_75t_L g3487 ( 
.A(n_2703),
.B(n_410),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_2918),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_2946),
.B(n_2977),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_2980),
.B(n_411),
.Y(n_3490)
);

A2O1A1Ixp33_ASAP7_75t_SL g3491 ( 
.A1(n_2876),
.A2(n_413),
.B(n_411),
.C(n_412),
.Y(n_3491)
);

AOI22xp33_ASAP7_75t_L g3492 ( 
.A1(n_2994),
.A2(n_414),
.B1(n_411),
.B2(n_412),
.Y(n_3492)
);

INVx2_ASAP7_75t_SL g3493 ( 
.A(n_2844),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_SL g3494 ( 
.A(n_3123),
.B(n_630),
.Y(n_3494)
);

INVxp67_ASAP7_75t_L g3495 ( 
.A(n_2672),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_L g3496 ( 
.A(n_3038),
.B(n_414),
.Y(n_3496)
);

OAI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_2826),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_3497)
);

OR2x6_ASAP7_75t_L g3498 ( 
.A(n_2558),
.B(n_415),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3046),
.B(n_415),
.Y(n_3499)
);

A2O1A1Ixp33_ASAP7_75t_SL g3500 ( 
.A1(n_2639),
.A2(n_418),
.B(n_416),
.C(n_417),
.Y(n_3500)
);

AND2x4_ASAP7_75t_L g3501 ( 
.A(n_2662),
.B(n_416),
.Y(n_3501)
);

OAI22xp5_ASAP7_75t_L g3502 ( 
.A1(n_3097),
.A2(n_419),
.B1(n_417),
.B2(n_418),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_2819),
.B(n_418),
.Y(n_3503)
);

INVx1_ASAP7_75t_SL g3504 ( 
.A(n_2857),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_SL g3505 ( 
.A(n_2757),
.B(n_630),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_2757),
.B(n_631),
.Y(n_3506)
);

AOI222xp33_ASAP7_75t_L g3507 ( 
.A1(n_3054),
.A2(n_421),
.B1(n_423),
.B2(n_419),
.C1(n_420),
.C2(n_422),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3064),
.B(n_420),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_SL g3509 ( 
.A(n_2757),
.B(n_631),
.Y(n_3509)
);

AOI21xp5_ASAP7_75t_L g3510 ( 
.A1(n_2961),
.A2(n_2963),
.B(n_2962),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3069),
.B(n_420),
.Y(n_3511)
);

OAI21xp33_ASAP7_75t_SL g3512 ( 
.A1(n_2931),
.A2(n_2951),
.B(n_2945),
.Y(n_3512)
);

O2A1O1Ixp5_ASAP7_75t_L g3513 ( 
.A1(n_2867),
.A2(n_423),
.B(n_421),
.C(n_422),
.Y(n_3513)
);

INVx6_ASAP7_75t_L g3514 ( 
.A(n_2865),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_2935),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_2940),
.Y(n_3516)
);

A2O1A1Ixp33_ASAP7_75t_L g3517 ( 
.A1(n_2968),
.A2(n_423),
.B(n_421),
.C(n_422),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_L g3518 ( 
.A(n_3082),
.B(n_3098),
.Y(n_3518)
);

AOI21xp5_ASAP7_75t_L g3519 ( 
.A1(n_2969),
.A2(n_424),
.B(n_425),
.Y(n_3519)
);

NOR2xp33_ASAP7_75t_L g3520 ( 
.A(n_3104),
.B(n_424),
.Y(n_3520)
);

NOR2xp33_ASAP7_75t_L g3521 ( 
.A(n_3105),
.B(n_424),
.Y(n_3521)
);

BUFx2_ASAP7_75t_L g3522 ( 
.A(n_2578),
.Y(n_3522)
);

INVx3_ASAP7_75t_L g3523 ( 
.A(n_2578),
.Y(n_3523)
);

NAND2x1_ASAP7_75t_L g3524 ( 
.A(n_2623),
.B(n_425),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3111),
.B(n_425),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_2720),
.Y(n_3526)
);

AOI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_2995),
.A2(n_426),
.B(n_427),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_2999),
.A2(n_426),
.B(n_427),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3120),
.B(n_426),
.Y(n_3529)
);

NOR2xp33_ASAP7_75t_L g3530 ( 
.A(n_2848),
.B(n_2849),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_SL g3531 ( 
.A(n_2780),
.B(n_634),
.Y(n_3531)
);

CKINVDCx5p33_ASAP7_75t_R g3532 ( 
.A(n_2546),
.Y(n_3532)
);

AND2x2_ASAP7_75t_L g3533 ( 
.A(n_2588),
.B(n_427),
.Y(n_3533)
);

NOR2xp33_ASAP7_75t_L g3534 ( 
.A(n_2850),
.B(n_428),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_2742),
.Y(n_3535)
);

OR2x2_ASAP7_75t_L g3536 ( 
.A(n_2749),
.B(n_2755),
.Y(n_3536)
);

BUFx8_ASAP7_75t_L g3537 ( 
.A(n_2865),
.Y(n_3537)
);

AOI21xp5_ASAP7_75t_L g3538 ( 
.A1(n_3004),
.A2(n_428),
.B(n_429),
.Y(n_3538)
);

OAI21x1_ASAP7_75t_L g3539 ( 
.A1(n_2950),
.A2(n_428),
.B(n_430),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_2959),
.Y(n_3540)
);

AND2x2_ASAP7_75t_L g3541 ( 
.A(n_2677),
.B(n_430),
.Y(n_3541)
);

AOI21xp5_ASAP7_75t_L g3542 ( 
.A1(n_3015),
.A2(n_3021),
.B(n_3017),
.Y(n_3542)
);

O2A1O1Ixp33_ASAP7_75t_L g3543 ( 
.A1(n_2794),
.A2(n_432),
.B(n_430),
.C(n_431),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_2953),
.Y(n_3544)
);

BUFx2_ASAP7_75t_L g3545 ( 
.A(n_2623),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_2682),
.B(n_431),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_2745),
.B(n_431),
.Y(n_3547)
);

CKINVDCx5p33_ASAP7_75t_R g3548 ( 
.A(n_2701),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_2533),
.B(n_432),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_2967),
.Y(n_3550)
);

CKINVDCx5p33_ASAP7_75t_R g3551 ( 
.A(n_2756),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_2695),
.B(n_433),
.Y(n_3552)
);

OAI22xp5_ASAP7_75t_L g3553 ( 
.A1(n_2783),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_SL g3554 ( 
.A(n_2780),
.B(n_634),
.Y(n_3554)
);

INVx4_ASAP7_75t_L g3555 ( 
.A(n_2780),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_2696),
.B(n_434),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_2966),
.Y(n_3557)
);

A2O1A1Ixp33_ASAP7_75t_L g3558 ( 
.A1(n_3033),
.A2(n_436),
.B(n_434),
.C(n_435),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_2791),
.B(n_436),
.Y(n_3559)
);

AND2x4_ASAP7_75t_L g3560 ( 
.A(n_2750),
.B(n_436),
.Y(n_3560)
);

OAI22xp5_ASAP7_75t_L g3561 ( 
.A1(n_2971),
.A2(n_440),
.B1(n_437),
.B2(n_438),
.Y(n_3561)
);

OAI22x1_ASAP7_75t_L g3562 ( 
.A1(n_2955),
.A2(n_441),
.B1(n_437),
.B2(n_440),
.Y(n_3562)
);

HB1xp67_ASAP7_75t_L g3563 ( 
.A(n_2729),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_2822),
.B(n_437),
.Y(n_3564)
);

AND2x4_ASAP7_75t_L g3565 ( 
.A(n_2750),
.B(n_440),
.Y(n_3565)
);

AOI22xp5_ASAP7_75t_L g3566 ( 
.A1(n_3005),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3010),
.Y(n_3567)
);

OAI22xp5_ASAP7_75t_L g3568 ( 
.A1(n_2981),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_3568)
);

OAI22xp5_ASAP7_75t_L g3569 ( 
.A1(n_2984),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_2985),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_3041),
.A2(n_444),
.B(n_445),
.Y(n_3571)
);

AOI22x1_ASAP7_75t_L g3572 ( 
.A1(n_3043),
.A2(n_448),
.B1(n_445),
.B2(n_446),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_SL g3573 ( 
.A(n_2842),
.B(n_635),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_2743),
.B(n_446),
.Y(n_3574)
);

A2O1A1Ixp33_ASAP7_75t_L g3575 ( 
.A1(n_3044),
.A2(n_450),
.B(n_448),
.C(n_449),
.Y(n_3575)
);

BUFx2_ASAP7_75t_L g3576 ( 
.A(n_2917),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_2728),
.B(n_448),
.Y(n_3577)
);

INVx8_ASAP7_75t_L g3578 ( 
.A(n_2842),
.Y(n_3578)
);

OAI22xp5_ASAP7_75t_L g3579 ( 
.A1(n_2987),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_2700),
.B(n_451),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_2709),
.B(n_453),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_2996),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3051),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_2997),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_3062),
.A2(n_453),
.B(n_454),
.Y(n_3585)
);

NOR2xp33_ASAP7_75t_L g3586 ( 
.A(n_3006),
.B(n_453),
.Y(n_3586)
);

CKINVDCx5p33_ASAP7_75t_R g3587 ( 
.A(n_2652),
.Y(n_3587)
);

AND2x4_ASAP7_75t_L g3588 ( 
.A(n_2917),
.B(n_454),
.Y(n_3588)
);

O2A1O1Ixp33_ASAP7_75t_L g3589 ( 
.A1(n_3056),
.A2(n_456),
.B(n_454),
.C(n_455),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3000),
.Y(n_3590)
);

AOI22xp5_ASAP7_75t_L g3591 ( 
.A1(n_3067),
.A2(n_458),
.B1(n_455),
.B2(n_457),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_2770),
.B(n_455),
.Y(n_3592)
);

BUFx8_ASAP7_75t_L g3593 ( 
.A(n_2872),
.Y(n_3593)
);

BUFx6f_ASAP7_75t_L g3594 ( 
.A(n_2842),
.Y(n_3594)
);

BUFx12f_ASAP7_75t_L g3595 ( 
.A(n_2595),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_2829),
.B(n_457),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_SL g3597 ( 
.A(n_2927),
.B(n_635),
.Y(n_3597)
);

BUFx3_ASAP7_75t_L g3598 ( 
.A(n_2929),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3003),
.Y(n_3599)
);

OAI22xp5_ASAP7_75t_L g3600 ( 
.A1(n_3012),
.A2(n_3013),
.B1(n_3020),
.B2(n_3019),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3024),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3030),
.Y(n_3602)
);

O2A1O1Ixp33_ASAP7_75t_L g3603 ( 
.A1(n_3068),
.A2(n_459),
.B(n_457),
.C(n_458),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3037),
.Y(n_3604)
);

OAI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_2846),
.A2(n_458),
.B(n_459),
.Y(n_3605)
);

BUFx3_ASAP7_75t_L g3606 ( 
.A(n_2929),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3042),
.B(n_459),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3048),
.B(n_460),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3049),
.B(n_460),
.Y(n_3609)
);

AOI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_3065),
.A2(n_460),
.B(n_461),
.Y(n_3610)
);

NAND2x1_ASAP7_75t_L g3611 ( 
.A(n_2979),
.B(n_461),
.Y(n_3611)
);

OAI22xp5_ASAP7_75t_L g3612 ( 
.A1(n_3050),
.A2(n_3057),
.B1(n_3063),
.B2(n_3058),
.Y(n_3612)
);

AOI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3071),
.A2(n_461),
.B(n_462),
.Y(n_3613)
);

NOR2xp33_ASAP7_75t_L g3614 ( 
.A(n_3153),
.B(n_462),
.Y(n_3614)
);

BUFx6f_ASAP7_75t_L g3615 ( 
.A(n_2979),
.Y(n_3615)
);

INVx4_ASAP7_75t_L g3616 ( 
.A(n_2983),
.Y(n_3616)
);

NOR2xp33_ASAP7_75t_L g3617 ( 
.A(n_3076),
.B(n_462),
.Y(n_3617)
);

AOI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_3083),
.A2(n_463),
.B(n_464),
.Y(n_3618)
);

AOI21x1_ASAP7_75t_L g3619 ( 
.A1(n_3091),
.A2(n_463),
.B(n_464),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_3129),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_3085),
.A2(n_464),
.B(n_465),
.Y(n_3621)
);

O2A1O1Ixp33_ASAP7_75t_L g3622 ( 
.A1(n_3077),
.A2(n_467),
.B(n_465),
.C(n_466),
.Y(n_3622)
);

O2A1O1Ixp33_ASAP7_75t_SL g3623 ( 
.A1(n_2869),
.A2(n_468),
.B(n_466),
.C(n_467),
.Y(n_3623)
);

NOR3xp33_ASAP7_75t_SL g3624 ( 
.A(n_3088),
.B(n_466),
.C(n_467),
.Y(n_3624)
);

OAI22xp5_ASAP7_75t_L g3625 ( 
.A1(n_3073),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3078),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3144),
.B(n_468),
.Y(n_3627)
);

INVx2_ASAP7_75t_SL g3628 ( 
.A(n_2861),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3079),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3081),
.B(n_469),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3095),
.B(n_471),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3103),
.B(n_471),
.Y(n_3632)
);

NOR2xp33_ASAP7_75t_L g3633 ( 
.A(n_3099),
.B(n_472),
.Y(n_3633)
);

OAI22xp5_ASAP7_75t_L g3634 ( 
.A1(n_3121),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_2779),
.B(n_474),
.Y(n_3635)
);

AO22x1_ASAP7_75t_L g3636 ( 
.A1(n_2866),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_3636)
);

NOR2xp33_ASAP7_75t_L g3637 ( 
.A(n_3119),
.B(n_475),
.Y(n_3637)
);

INVx6_ASAP7_75t_L g3638 ( 
.A(n_2812),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_2786),
.B(n_476),
.Y(n_3639)
);

NOR2x1_ASAP7_75t_L g3640 ( 
.A(n_2645),
.B(n_476),
.Y(n_3640)
);

NOR2xp33_ASAP7_75t_L g3641 ( 
.A(n_2796),
.B(n_477),
.Y(n_3641)
);

OAI22xp5_ASAP7_75t_L g3642 ( 
.A1(n_3126),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3100),
.A2(n_478),
.B(n_479),
.Y(n_3643)
);

AND2x4_ASAP7_75t_L g3644 ( 
.A(n_2983),
.B(n_478),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3134),
.Y(n_3645)
);

BUFx3_ASAP7_75t_L g3646 ( 
.A(n_3018),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3135),
.Y(n_3647)
);

AOI222xp33_ASAP7_75t_L g3648 ( 
.A1(n_2612),
.A2(n_481),
.B1(n_483),
.B2(n_479),
.C1(n_480),
.C2(n_482),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3140),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3143),
.Y(n_3650)
);

AOI21xp5_ASAP7_75t_L g3651 ( 
.A1(n_3101),
.A2(n_3108),
.B(n_3107),
.Y(n_3651)
);

CKINVDCx5p33_ASAP7_75t_R g3652 ( 
.A(n_2659),
.Y(n_3652)
);

AOI21x1_ASAP7_75t_L g3653 ( 
.A1(n_2603),
.A2(n_482),
.B(n_485),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_2761),
.Y(n_3654)
);

INVx2_ASAP7_75t_SL g3655 ( 
.A(n_3018),
.Y(n_3655)
);

INVx3_ASAP7_75t_L g3656 ( 
.A(n_3113),
.Y(n_3656)
);

AOI21xp5_ASAP7_75t_L g3657 ( 
.A1(n_3115),
.A2(n_485),
.B(n_486),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_2762),
.Y(n_3658)
);

AOI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_3117),
.A2(n_485),
.B(n_486),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_2693),
.Y(n_3660)
);

BUFx2_ASAP7_75t_L g3661 ( 
.A(n_3113),
.Y(n_3661)
);

CKINVDCx5p33_ASAP7_75t_R g3662 ( 
.A(n_2877),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_2948),
.Y(n_3663)
);

O2A1O1Ixp33_ASAP7_75t_L g3664 ( 
.A1(n_2684),
.A2(n_488),
.B(n_486),
.C(n_487),
.Y(n_3664)
);

OAI21xp33_ASAP7_75t_L g3665 ( 
.A1(n_2697),
.A2(n_487),
.B(n_488),
.Y(n_3665)
);

BUFx6f_ASAP7_75t_L g3666 ( 
.A(n_2853),
.Y(n_3666)
);

O2A1O1Ixp33_ASAP7_75t_L g3667 ( 
.A1(n_2790),
.A2(n_489),
.B(n_487),
.C(n_488),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_2713),
.B(n_489),
.Y(n_3668)
);

AOI21xp5_ASAP7_75t_L g3669 ( 
.A1(n_3124),
.A2(n_3127),
.B(n_3125),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_SL g3670 ( 
.A(n_3139),
.B(n_636),
.Y(n_3670)
);

AOI21xp5_ASAP7_75t_L g3671 ( 
.A1(n_3131),
.A2(n_490),
.B(n_491),
.Y(n_3671)
);

INVx3_ASAP7_75t_L g3672 ( 
.A(n_2853),
.Y(n_3672)
);

NAND3xp33_ASAP7_75t_L g3673 ( 
.A(n_2626),
.B(n_490),
.C(n_491),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_2785),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_2718),
.B(n_490),
.Y(n_3675)
);

CKINVDCx5p33_ASAP7_75t_R g3676 ( 
.A(n_2947),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_2825),
.Y(n_3677)
);

CKINVDCx5p33_ASAP7_75t_R g3678 ( 
.A(n_2982),
.Y(n_3678)
);

OAI21x1_ASAP7_75t_L g3679 ( 
.A1(n_2538),
.A2(n_491),
.B(n_492),
.Y(n_3679)
);

OAI22xp5_ASAP7_75t_L g3680 ( 
.A1(n_2719),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_3680)
);

NOR2xp33_ASAP7_75t_R g3681 ( 
.A(n_2862),
.B(n_493),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_2726),
.B(n_494),
.Y(n_3682)
);

INVxp67_ASAP7_75t_L g3683 ( 
.A(n_2855),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_2535),
.B(n_495),
.Y(n_3684)
);

AOI21xp5_ASAP7_75t_L g3685 ( 
.A1(n_3133),
.A2(n_495),
.B(n_496),
.Y(n_3685)
);

BUFx3_ASAP7_75t_L g3686 ( 
.A(n_3232),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3157),
.Y(n_3687)
);

OAI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_3518),
.A2(n_3141),
.B(n_3138),
.Y(n_3688)
);

A2O1A1Ixp33_ASAP7_75t_L g3689 ( 
.A1(n_3664),
.A2(n_2830),
.B(n_2581),
.C(n_2597),
.Y(n_3689)
);

AOI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_3158),
.A2(n_3147),
.B(n_3142),
.Y(n_3690)
);

OAI21xp5_ASAP7_75t_L g3691 ( 
.A1(n_3431),
.A2(n_2613),
.B(n_2605),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3295),
.Y(n_3692)
);

OAI22x1_ASAP7_75t_L g3693 ( 
.A1(n_3444),
.A2(n_2615),
.B1(n_2860),
.B2(n_2856),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3214),
.B(n_2630),
.Y(n_3694)
);

AOI21xp5_ASAP7_75t_L g3695 ( 
.A1(n_3163),
.A2(n_3542),
.B(n_3510),
.Y(n_3695)
);

AND2x2_ASAP7_75t_L g3696 ( 
.A(n_3503),
.B(n_2854),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3298),
.Y(n_3697)
);

OAI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_3184),
.A2(n_2611),
.B(n_2604),
.Y(n_3698)
);

OAI22xp5_ASAP7_75t_L g3699 ( 
.A1(n_3221),
.A2(n_2741),
.B1(n_2805),
.B2(n_2651),
.Y(n_3699)
);

AND2x4_ASAP7_75t_L g3700 ( 
.A(n_3197),
.B(n_2862),
.Y(n_3700)
);

CKINVDCx20_ASAP7_75t_R g3701 ( 
.A(n_3242),
.Y(n_3701)
);

OAI21x1_ASAP7_75t_L g3702 ( 
.A1(n_3660),
.A2(n_2542),
.B(n_2541),
.Y(n_3702)
);

NAND2x1_ASAP7_75t_L g3703 ( 
.A(n_3341),
.B(n_3348),
.Y(n_3703)
);

OAI22xp5_ASAP7_75t_L g3704 ( 
.A1(n_3205),
.A2(n_2637),
.B1(n_2733),
.B2(n_2903),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3587),
.B(n_2633),
.Y(n_3705)
);

AOI221xp5_ASAP7_75t_SL g3706 ( 
.A1(n_3458),
.A2(n_2680),
.B1(n_2648),
.B2(n_2618),
.C(n_2617),
.Y(n_3706)
);

A2O1A1Ixp33_ASAP7_75t_L g3707 ( 
.A1(n_3667),
.A2(n_2600),
.B(n_2976),
.C(n_2884),
.Y(n_3707)
);

BUFx2_ASAP7_75t_L g3708 ( 
.A(n_3407),
.Y(n_3708)
);

AO31x2_ASAP7_75t_L g3709 ( 
.A1(n_3544),
.A2(n_2649),
.A3(n_3026),
.B(n_2817),
.Y(n_3709)
);

BUFx3_ASAP7_75t_L g3710 ( 
.A(n_3259),
.Y(n_3710)
);

AOI22xp33_ASAP7_75t_L g3711 ( 
.A1(n_3366),
.A2(n_3354),
.B1(n_3676),
.B2(n_3662),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_SL g3712 ( 
.A(n_3205),
.B(n_2902),
.Y(n_3712)
);

INVx3_ASAP7_75t_L g3713 ( 
.A(n_3197),
.Y(n_3713)
);

O2A1O1Ixp33_ASAP7_75t_SL g3714 ( 
.A1(n_3309),
.A2(n_2989),
.B(n_2992),
.C(n_2944),
.Y(n_3714)
);

BUFx6f_ASAP7_75t_L g3715 ( 
.A(n_3197),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3162),
.Y(n_3716)
);

AOI22xp5_ASAP7_75t_L g3717 ( 
.A1(n_3678),
.A2(n_3023),
.B1(n_2986),
.B2(n_2800),
.Y(n_3717)
);

O2A1O1Ixp33_ASAP7_75t_SL g3718 ( 
.A1(n_3159),
.A2(n_3187),
.B(n_3364),
.C(n_3239),
.Y(n_3718)
);

CKINVDCx11_ASAP7_75t_R g3719 ( 
.A(n_3179),
.Y(n_3719)
);

AOI221xp5_ASAP7_75t_L g3720 ( 
.A1(n_3301),
.A2(n_3060),
.B1(n_3137),
.B2(n_3039),
.C(n_2990),
.Y(n_3720)
);

AOI21x1_ASAP7_75t_L g3721 ( 
.A1(n_3550),
.A2(n_3583),
.B(n_3567),
.Y(n_3721)
);

BUFx2_ASAP7_75t_R g3722 ( 
.A(n_3169),
.Y(n_3722)
);

AOI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_3651),
.A2(n_2550),
.B(n_2832),
.Y(n_3723)
);

OR2x2_ASAP7_75t_L g3724 ( 
.A(n_3397),
.B(n_2781),
.Y(n_3724)
);

CKINVDCx20_ASAP7_75t_R g3725 ( 
.A(n_3248),
.Y(n_3725)
);

OAI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_3600),
.A2(n_2616),
.B(n_2625),
.Y(n_3726)
);

OAI22xp5_ASAP7_75t_L g3727 ( 
.A1(n_3205),
.A2(n_3025),
.B1(n_3118),
.B2(n_3112),
.Y(n_3727)
);

AO31x2_ASAP7_75t_L g3728 ( 
.A1(n_3620),
.A2(n_3190),
.A3(n_3222),
.B(n_3669),
.Y(n_3728)
);

AOI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_3306),
.A2(n_2545),
.B(n_2670),
.Y(n_3729)
);

BUFx6f_ASAP7_75t_L g3730 ( 
.A(n_3198),
.Y(n_3730)
);

AOI31xp67_ASAP7_75t_L g3731 ( 
.A1(n_3677),
.A2(n_2699),
.A3(n_2708),
.B(n_2702),
.Y(n_3731)
);

CKINVDCx5p33_ASAP7_75t_R g3732 ( 
.A(n_3171),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3652),
.B(n_2635),
.Y(n_3733)
);

AOI22xp33_ASAP7_75t_L g3734 ( 
.A1(n_3537),
.A2(n_2747),
.B1(n_2628),
.B2(n_2656),
.Y(n_3734)
);

OAI21xp5_ASAP7_75t_L g3735 ( 
.A1(n_3612),
.A2(n_2653),
.B(n_2655),
.Y(n_3735)
);

AOI21xp5_ASAP7_75t_L g3736 ( 
.A1(n_3264),
.A2(n_2759),
.B(n_2868),
.Y(n_3736)
);

OAI21xp5_ASAP7_75t_L g3737 ( 
.A1(n_3512),
.A2(n_2669),
.B(n_2666),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3164),
.Y(n_3738)
);

OR2x2_ASAP7_75t_L g3739 ( 
.A(n_3235),
.B(n_2554),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3276),
.B(n_495),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3168),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_3284),
.A2(n_2821),
.B(n_2851),
.Y(n_3742)
);

OAI21xp5_ASAP7_75t_L g3743 ( 
.A1(n_3451),
.A2(n_3489),
.B(n_3673),
.Y(n_3743)
);

INVx4_ASAP7_75t_L g3744 ( 
.A(n_3198),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_3433),
.A2(n_2723),
.B(n_2608),
.Y(n_3745)
);

A2O1A1Ixp33_ASAP7_75t_L g3746 ( 
.A1(n_3201),
.A2(n_3148),
.B(n_2847),
.C(n_2835),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3303),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3218),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3404),
.B(n_2636),
.Y(n_3749)
);

OAI21x1_ASAP7_75t_L g3750 ( 
.A1(n_3421),
.A2(n_2751),
.B(n_2748),
.Y(n_3750)
);

OAI21x1_ASAP7_75t_SL g3751 ( 
.A1(n_3430),
.A2(n_2727),
.B(n_2823),
.Y(n_3751)
);

AO32x2_ASAP7_75t_L g3752 ( 
.A1(n_3237),
.A2(n_2803),
.A3(n_2624),
.B1(n_2814),
.B2(n_2810),
.Y(n_3752)
);

INVx2_ASAP7_75t_SL g3753 ( 
.A(n_3198),
.Y(n_3753)
);

INVx1_ASAP7_75t_SL g3754 ( 
.A(n_3446),
.Y(n_3754)
);

AOI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_3480),
.A2(n_2811),
.B(n_2771),
.Y(n_3755)
);

AND2x2_ASAP7_75t_SL g3756 ( 
.A(n_3426),
.B(n_2873),
.Y(n_3756)
);

BUFx12f_ASAP7_75t_L g3757 ( 
.A(n_3186),
.Y(n_3757)
);

INVxp67_ASAP7_75t_L g3758 ( 
.A(n_3254),
.Y(n_3758)
);

AOI21xp5_ASAP7_75t_L g3759 ( 
.A1(n_3410),
.A2(n_2763),
.B(n_2758),
.Y(n_3759)
);

AOI21xp5_ASAP7_75t_L g3760 ( 
.A1(n_3663),
.A2(n_2707),
.B(n_2704),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3294),
.B(n_496),
.Y(n_3761)
);

AOI21xp5_ASAP7_75t_L g3762 ( 
.A1(n_3414),
.A2(n_2683),
.B(n_2676),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3304),
.Y(n_3763)
);

O2A1O1Ixp33_ASAP7_75t_SL g3764 ( 
.A1(n_3385),
.A2(n_2874),
.B(n_2716),
.C(n_2795),
.Y(n_3764)
);

AOI21xp33_ASAP7_75t_L g3765 ( 
.A1(n_3206),
.A2(n_2787),
.B(n_2772),
.Y(n_3765)
);

BUFx6f_ASAP7_75t_L g3766 ( 
.A(n_3176),
.Y(n_3766)
);

AOI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_3417),
.A2(n_2692),
.B(n_2766),
.Y(n_3767)
);

OAI221xp5_ASAP7_75t_L g3768 ( 
.A1(n_3495),
.A2(n_3240),
.B1(n_3277),
.B2(n_3266),
.C(n_3376),
.Y(n_3768)
);

NOR3xp33_ASAP7_75t_L g3769 ( 
.A(n_3204),
.B(n_2793),
.C(n_2852),
.Y(n_3769)
);

BUFx2_ASAP7_75t_L g3770 ( 
.A(n_3460),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3307),
.Y(n_3771)
);

A2O1A1Ixp33_ASAP7_75t_L g3772 ( 
.A1(n_3290),
.A2(n_2769),
.B(n_2792),
.C(n_2773),
.Y(n_3772)
);

OAI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3211),
.A2(n_2864),
.B(n_2859),
.Y(n_3773)
);

BUFx6f_ASAP7_75t_SL g3774 ( 
.A(n_3256),
.Y(n_3774)
);

OAI22xp5_ASAP7_75t_L g3775 ( 
.A1(n_3479),
.A2(n_2834),
.B1(n_2875),
.B2(n_2799),
.Y(n_3775)
);

AOI21xp5_ASAP7_75t_L g3776 ( 
.A1(n_3175),
.A2(n_2804),
.B(n_2831),
.Y(n_3776)
);

AND2x2_ASAP7_75t_L g3777 ( 
.A(n_3563),
.B(n_496),
.Y(n_3777)
);

OAI21x1_ASAP7_75t_L g3778 ( 
.A1(n_3400),
.A2(n_2831),
.B(n_2799),
.Y(n_3778)
);

AOI21xp5_ASAP7_75t_L g3779 ( 
.A1(n_3500),
.A2(n_2764),
.B(n_497),
.Y(n_3779)
);

AND2x4_ASAP7_75t_L g3780 ( 
.A(n_3378),
.B(n_3424),
.Y(n_3780)
);

BUFx3_ASAP7_75t_L g3781 ( 
.A(n_3478),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3357),
.A2(n_2764),
.B(n_497),
.Y(n_3782)
);

OAI21xp5_ASAP7_75t_L g3783 ( 
.A1(n_3513),
.A2(n_498),
.B(n_499),
.Y(n_3783)
);

CKINVDCx20_ASAP7_75t_R g3784 ( 
.A(n_3278),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3200),
.B(n_3208),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3216),
.B(n_498),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3320),
.Y(n_3787)
);

BUFx4f_ASAP7_75t_SL g3788 ( 
.A(n_3319),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3327),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3328),
.Y(n_3790)
);

INVx1_ASAP7_75t_SL g3791 ( 
.A(n_3472),
.Y(n_3791)
);

NAND2xp33_ASAP7_75t_L g3792 ( 
.A(n_3225),
.B(n_498),
.Y(n_3792)
);

BUFx2_ASAP7_75t_L g3793 ( 
.A(n_3378),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3335),
.Y(n_3794)
);

INVx2_ASAP7_75t_L g3795 ( 
.A(n_3238),
.Y(n_3795)
);

A2O1A1Ixp33_ASAP7_75t_L g3796 ( 
.A1(n_3280),
.A2(n_501),
.B(n_499),
.C(n_500),
.Y(n_3796)
);

OAI21x1_ASAP7_75t_L g3797 ( 
.A1(n_3400),
.A2(n_501),
.B(n_500),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3395),
.B(n_499),
.Y(n_3798)
);

OAI22xp5_ASAP7_75t_L g3799 ( 
.A1(n_3225),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.Y(n_3799)
);

AOI21xp5_ASAP7_75t_L g3800 ( 
.A1(n_3411),
.A2(n_502),
.B(n_503),
.Y(n_3800)
);

INVx3_ASAP7_75t_L g3801 ( 
.A(n_3424),
.Y(n_3801)
);

AND2x4_ASAP7_75t_L g3802 ( 
.A(n_3449),
.B(n_502),
.Y(n_3802)
);

AOI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3597),
.A2(n_503),
.B(n_504),
.Y(n_3803)
);

OR2x2_ASAP7_75t_L g3804 ( 
.A(n_3504),
.B(n_3160),
.Y(n_3804)
);

A2O1A1Ixp33_ASAP7_75t_L g3805 ( 
.A1(n_3263),
.A2(n_507),
.B(n_505),
.C(n_506),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3340),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3223),
.B(n_505),
.Y(n_3807)
);

AOI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3670),
.A2(n_3456),
.B(n_3403),
.Y(n_3808)
);

O2A1O1Ixp33_ASAP7_75t_L g3809 ( 
.A1(n_3491),
.A2(n_507),
.B(n_505),
.C(n_506),
.Y(n_3809)
);

AO31x2_ASAP7_75t_L g3810 ( 
.A1(n_3443),
.A2(n_508),
.A3(n_506),
.B(n_507),
.Y(n_3810)
);

AOI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_3440),
.A2(n_508),
.B(n_509),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3224),
.B(n_509),
.Y(n_3812)
);

OAI21x1_ASAP7_75t_L g3813 ( 
.A1(n_3423),
.A2(n_511),
.B(n_510),
.Y(n_3813)
);

OAI21x1_ASAP7_75t_L g3814 ( 
.A1(n_3423),
.A2(n_511),
.B(n_510),
.Y(n_3814)
);

AND2x4_ASAP7_75t_L g3815 ( 
.A(n_3449),
.B(n_509),
.Y(n_3815)
);

A2O1A1Ixp33_ASAP7_75t_L g3816 ( 
.A1(n_3262),
.A2(n_512),
.B(n_510),
.C(n_511),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_SL g3817 ( 
.A(n_3501),
.B(n_512),
.Y(n_3817)
);

A2O1A1Ixp33_ASAP7_75t_L g3818 ( 
.A1(n_3466),
.A2(n_514),
.B(n_512),
.C(n_513),
.Y(n_3818)
);

OA21x2_ASAP7_75t_L g3819 ( 
.A1(n_3539),
.A2(n_513),
.B(n_514),
.Y(n_3819)
);

BUFx2_ASAP7_75t_L g3820 ( 
.A(n_3537),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3257),
.B(n_515),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3453),
.A2(n_515),
.B(n_516),
.Y(n_3822)
);

AOI221xp5_ASAP7_75t_SL g3823 ( 
.A1(n_3314),
.A2(n_3289),
.B1(n_3322),
.B2(n_3316),
.C(n_3370),
.Y(n_3823)
);

AO32x2_ASAP7_75t_L g3824 ( 
.A1(n_3209),
.A2(n_3226),
.A3(n_3245),
.B1(n_3229),
.B2(n_3188),
.Y(n_3824)
);

OR2x6_ASAP7_75t_L g3825 ( 
.A(n_3345),
.B(n_516),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3347),
.Y(n_3826)
);

AO31x2_ASAP7_75t_L g3827 ( 
.A1(n_3435),
.A2(n_518),
.A3(n_516),
.B(n_517),
.Y(n_3827)
);

OAI21x1_ASAP7_75t_L g3828 ( 
.A1(n_3619),
.A2(n_3302),
.B(n_3286),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3457),
.A2(n_517),
.B(n_519),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3349),
.Y(n_3830)
);

NOR2xp33_ASAP7_75t_SL g3831 ( 
.A(n_3345),
.B(n_517),
.Y(n_3831)
);

AOI221x1_ASAP7_75t_L g3832 ( 
.A1(n_3439),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.C(n_522),
.Y(n_3832)
);

AOI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3462),
.A2(n_519),
.B(n_520),
.Y(n_3833)
);

NAND2xp33_ASAP7_75t_L g3834 ( 
.A(n_3432),
.B(n_520),
.Y(n_3834)
);

INVx3_ASAP7_75t_SL g3835 ( 
.A(n_3252),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3268),
.B(n_521),
.Y(n_3836)
);

OAI21xp5_ASAP7_75t_L g3837 ( 
.A1(n_3641),
.A2(n_521),
.B(n_522),
.Y(n_3837)
);

BUFx3_ASAP7_75t_L g3838 ( 
.A(n_3321),
.Y(n_3838)
);

NOR2xp33_ASAP7_75t_L g3839 ( 
.A(n_3165),
.B(n_522),
.Y(n_3839)
);

BUFx6f_ASAP7_75t_L g3840 ( 
.A(n_3420),
.Y(n_3840)
);

NOR4xp25_ASAP7_75t_L g3841 ( 
.A(n_3177),
.B(n_525),
.C(n_523),
.D(n_524),
.Y(n_3841)
);

OR2x6_ASAP7_75t_L g3842 ( 
.A(n_3338),
.B(n_524),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3399),
.B(n_524),
.Y(n_3843)
);

O2A1O1Ixp5_ASAP7_75t_SL g3844 ( 
.A1(n_3311),
.A2(n_637),
.B(n_638),
.C(n_636),
.Y(n_3844)
);

AOI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_3469),
.A2(n_3485),
.B(n_3477),
.Y(n_3845)
);

NOR4xp25_ASAP7_75t_L g3846 ( 
.A(n_3454),
.B(n_3172),
.C(n_3361),
.D(n_3331),
.Y(n_3846)
);

OAI21xp5_ASAP7_75t_L g3847 ( 
.A1(n_3428),
.A2(n_525),
.B(n_526),
.Y(n_3847)
);

OAI21xp5_ASAP7_75t_L g3848 ( 
.A1(n_3468),
.A2(n_525),
.B(n_526),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3488),
.A2(n_527),
.B(n_528),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3260),
.Y(n_3850)
);

OAI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_3481),
.A2(n_527),
.B(n_528),
.Y(n_3851)
);

NOR2xp33_ASAP7_75t_L g3852 ( 
.A(n_3514),
.B(n_528),
.Y(n_3852)
);

OA21x2_ASAP7_75t_L g3853 ( 
.A1(n_3213),
.A2(n_529),
.B(n_530),
.Y(n_3853)
);

O2A1O1Ixp33_ASAP7_75t_SL g3854 ( 
.A1(n_3333),
.A2(n_531),
.B(n_529),
.C(n_530),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3398),
.Y(n_3855)
);

AOI21x1_ASAP7_75t_L g3856 ( 
.A1(n_3282),
.A2(n_639),
.B(n_637),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3445),
.B(n_529),
.Y(n_3857)
);

INVx3_ASAP7_75t_SL g3858 ( 
.A(n_3267),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3325),
.Y(n_3859)
);

AOI21xp5_ASAP7_75t_L g3860 ( 
.A1(n_3515),
.A2(n_531),
.B(n_532),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3387),
.B(n_531),
.Y(n_3861)
);

AOI21xp5_ASAP7_75t_L g3862 ( 
.A1(n_3516),
.A2(n_532),
.B(n_533),
.Y(n_3862)
);

NAND2x1p5_ASAP7_75t_L g3863 ( 
.A(n_3183),
.B(n_533),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3279),
.Y(n_3864)
);

BUFx10_ASAP7_75t_L g3865 ( 
.A(n_3323),
.Y(n_3865)
);

OAI22xp5_ASAP7_75t_L g3866 ( 
.A1(n_3487),
.A2(n_536),
.B1(n_534),
.B2(n_535),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3283),
.Y(n_3867)
);

OR2x2_ASAP7_75t_L g3868 ( 
.A(n_3291),
.B(n_534),
.Y(n_3868)
);

OAI21x1_ASAP7_75t_L g3869 ( 
.A1(n_3286),
.A2(n_536),
.B(n_535),
.Y(n_3869)
);

INVxp67_ASAP7_75t_SL g3870 ( 
.A(n_3413),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_3540),
.B(n_534),
.Y(n_3871)
);

AOI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3557),
.A2(n_535),
.B(n_536),
.Y(n_3872)
);

AO21x2_ASAP7_75t_L g3873 ( 
.A1(n_3665),
.A2(n_537),
.B(n_538),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3570),
.B(n_537),
.Y(n_3874)
);

NOR2xp33_ASAP7_75t_L g3875 ( 
.A(n_3514),
.B(n_3551),
.Y(n_3875)
);

OAI21x1_ASAP7_75t_L g3876 ( 
.A1(n_3302),
.A2(n_539),
.B(n_538),
.Y(n_3876)
);

OR2x6_ASAP7_75t_L g3877 ( 
.A(n_3338),
.B(n_537),
.Y(n_3877)
);

BUFx6f_ASAP7_75t_L g3878 ( 
.A(n_3271),
.Y(n_3878)
);

INVx1_ASAP7_75t_SL g3879 ( 
.A(n_3548),
.Y(n_3879)
);

AOI21xp5_ASAP7_75t_L g3880 ( 
.A1(n_3582),
.A2(n_538),
.B(n_539),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_3584),
.A2(n_540),
.B(n_541),
.Y(n_3881)
);

AOI22xp5_ASAP7_75t_L g3882 ( 
.A1(n_3390),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_3882)
);

INVx2_ASAP7_75t_L g3883 ( 
.A(n_3274),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3590),
.A2(n_540),
.B(n_542),
.Y(n_3884)
);

AO21x1_ASAP7_75t_L g3885 ( 
.A1(n_3487),
.A2(n_3501),
.B(n_3497),
.Y(n_3885)
);

AO31x2_ASAP7_75t_L g3886 ( 
.A1(n_3438),
.A2(n_545),
.A3(n_543),
.B(n_544),
.Y(n_3886)
);

BUFx2_ASAP7_75t_L g3887 ( 
.A(n_3593),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3384),
.Y(n_3888)
);

OAI21x1_ASAP7_75t_L g3889 ( 
.A1(n_3382),
.A2(n_545),
.B(n_544),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3297),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_3599),
.A2(n_543),
.B(n_546),
.Y(n_3891)
);

AOI21xp5_ASAP7_75t_L g3892 ( 
.A1(n_3601),
.A2(n_546),
.B(n_547),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3425),
.B(n_546),
.Y(n_3893)
);

O2A1O1Ixp33_ASAP7_75t_L g3894 ( 
.A1(n_3353),
.A2(n_3484),
.B(n_3494),
.C(n_3471),
.Y(n_3894)
);

HB1xp67_ASAP7_75t_L g3895 ( 
.A(n_3247),
.Y(n_3895)
);

OR2x2_ASAP7_75t_L g3896 ( 
.A(n_3388),
.B(n_547),
.Y(n_3896)
);

AOI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_3602),
.A2(n_548),
.B(n_549),
.Y(n_3897)
);

AO31x2_ASAP7_75t_L g3898 ( 
.A1(n_3441),
.A2(n_550),
.A3(n_548),
.B(n_549),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_3604),
.B(n_548),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_3300),
.Y(n_3900)
);

AO21x2_ASAP7_75t_L g3901 ( 
.A1(n_3653),
.A2(n_550),
.B(n_551),
.Y(n_3901)
);

O2A1O1Ixp33_ASAP7_75t_L g3902 ( 
.A1(n_3167),
.A2(n_552),
.B(n_550),
.C(n_551),
.Y(n_3902)
);

INVx4_ASAP7_75t_L g3903 ( 
.A(n_3219),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3626),
.B(n_551),
.Y(n_3904)
);

NOR2xp33_ASAP7_75t_L g3905 ( 
.A(n_3299),
.B(n_552),
.Y(n_3905)
);

OAI21x1_ASAP7_75t_L g3906 ( 
.A1(n_3382),
.A2(n_552),
.B(n_553),
.Y(n_3906)
);

A2O1A1Ixp33_ASAP7_75t_L g3907 ( 
.A1(n_3543),
.A2(n_555),
.B(n_553),
.C(n_554),
.Y(n_3907)
);

A2O1A1Ixp33_ASAP7_75t_L g3908 ( 
.A1(n_3408),
.A2(n_556),
.B(n_554),
.C(n_555),
.Y(n_3908)
);

BUFx6f_ASAP7_75t_L g3909 ( 
.A(n_3271),
.Y(n_3909)
);

OAI22x1_ASAP7_75t_L g3910 ( 
.A1(n_3183),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.Y(n_3910)
);

AOI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3496),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3629),
.B(n_557),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_3645),
.B(n_558),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3647),
.B(n_558),
.Y(n_3914)
);

INVx2_ASAP7_75t_L g3915 ( 
.A(n_3312),
.Y(n_3915)
);

BUFx12f_ASAP7_75t_L g3916 ( 
.A(n_3638),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3649),
.A2(n_560),
.B(n_561),
.Y(n_3917)
);

OAI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_3270),
.A2(n_560),
.B(n_562),
.Y(n_3918)
);

AOI21xp5_ASAP7_75t_L g3919 ( 
.A1(n_3650),
.A2(n_3674),
.B(n_3668),
.Y(n_3919)
);

OAI21x1_ASAP7_75t_L g3920 ( 
.A1(n_3234),
.A2(n_560),
.B(n_562),
.Y(n_3920)
);

INVx2_ASAP7_75t_L g3921 ( 
.A(n_3315),
.Y(n_3921)
);

AOI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_3675),
.A2(n_562),
.B(n_563),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3352),
.B(n_563),
.Y(n_3923)
);

AOI21xp5_ASAP7_75t_L g3924 ( 
.A1(n_3682),
.A2(n_563),
.B(n_564),
.Y(n_3924)
);

AO31x2_ASAP7_75t_L g3925 ( 
.A1(n_3463),
.A2(n_566),
.A3(n_564),
.B(n_565),
.Y(n_3925)
);

INVx2_ASAP7_75t_SL g3926 ( 
.A(n_3467),
.Y(n_3926)
);

AOI21xp5_ASAP7_75t_L g3927 ( 
.A1(n_3577),
.A2(n_564),
.B(n_565),
.Y(n_3927)
);

INVx4_ASAP7_75t_L g3928 ( 
.A(n_3220),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3196),
.B(n_565),
.Y(n_3929)
);

OA21x2_ASAP7_75t_L g3930 ( 
.A1(n_3679),
.A2(n_566),
.B(n_567),
.Y(n_3930)
);

A2O1A1Ixp33_ASAP7_75t_L g3931 ( 
.A1(n_3442),
.A2(n_3362),
.B(n_3603),
.C(n_3589),
.Y(n_3931)
);

AOI21xp5_ASAP7_75t_L g3932 ( 
.A1(n_3628),
.A2(n_566),
.B(n_568),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3202),
.B(n_568),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3658),
.Y(n_3934)
);

OAI21x1_ASAP7_75t_L g3935 ( 
.A1(n_3464),
.A2(n_569),
.B(n_570),
.Y(n_3935)
);

OAI21x1_ASAP7_75t_L g3936 ( 
.A1(n_3523),
.A2(n_569),
.B(n_570),
.Y(n_3936)
);

NOR2xp33_ASAP7_75t_SL g3937 ( 
.A(n_3638),
.B(n_569),
.Y(n_3937)
);

INVx2_ASAP7_75t_SL g3938 ( 
.A(n_3593),
.Y(n_3938)
);

NOR4xp25_ASAP7_75t_L g3939 ( 
.A(n_3192),
.B(n_573),
.C(n_571),
.D(n_572),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3346),
.Y(n_3940)
);

A2O1A1Ixp33_ASAP7_75t_L g3941 ( 
.A1(n_3622),
.A2(n_573),
.B(n_571),
.C(n_572),
.Y(n_3941)
);

BUFx2_ASAP7_75t_L g3942 ( 
.A(n_3681),
.Y(n_3942)
);

AOI22xp33_ASAP7_75t_L g3943 ( 
.A1(n_3520),
.A2(n_3521),
.B1(n_3429),
.B2(n_3447),
.Y(n_3943)
);

AO32x2_ASAP7_75t_L g3944 ( 
.A1(n_3483),
.A2(n_574),
.A3(n_571),
.B1(n_573),
.B2(n_575),
.Y(n_3944)
);

OAI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_3683),
.A2(n_3377),
.B(n_3368),
.Y(n_3945)
);

O2A1O1Ixp33_ASAP7_75t_L g3946 ( 
.A1(n_3437),
.A2(n_577),
.B(n_574),
.C(n_576),
.Y(n_3946)
);

BUFx3_ASAP7_75t_L g3947 ( 
.A(n_3371),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3365),
.Y(n_3948)
);

AOI211x1_ASAP7_75t_L g3949 ( 
.A1(n_3636),
.A2(n_577),
.B(n_574),
.C(n_576),
.Y(n_3949)
);

A2O1A1Ixp33_ASAP7_75t_L g3950 ( 
.A1(n_3486),
.A2(n_579),
.B(n_576),
.C(n_578),
.Y(n_3950)
);

AOI221xp5_ASAP7_75t_L g3951 ( 
.A1(n_3373),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.C(n_581),
.Y(n_3951)
);

OAI21xp5_ASAP7_75t_L g3952 ( 
.A1(n_3380),
.A2(n_579),
.B(n_580),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3393),
.Y(n_3953)
);

OA21x2_ASAP7_75t_L g3954 ( 
.A1(n_3217),
.A2(n_580),
.B(n_581),
.Y(n_3954)
);

OAI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3416),
.A2(n_581),
.B(n_582),
.Y(n_3955)
);

AOI221x1_ASAP7_75t_L g3956 ( 
.A1(n_3562),
.A2(n_584),
.B1(n_582),
.B2(n_583),
.C(n_585),
.Y(n_3956)
);

OAI21xp5_ASAP7_75t_L g3957 ( 
.A1(n_3419),
.A2(n_582),
.B(n_583),
.Y(n_3957)
);

OAI21x1_ASAP7_75t_L g3958 ( 
.A1(n_3523),
.A2(n_583),
.B(n_584),
.Y(n_3958)
);

A2O1A1Ixp33_ASAP7_75t_L g3959 ( 
.A1(n_3605),
.A2(n_3308),
.B(n_3161),
.C(n_3339),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3654),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3374),
.Y(n_3961)
);

OAI21x1_ASAP7_75t_L g3962 ( 
.A1(n_3656),
.A2(n_584),
.B(n_585),
.Y(n_3962)
);

CKINVDCx11_ASAP7_75t_R g3963 ( 
.A(n_3244),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3231),
.B(n_585),
.Y(n_3964)
);

AO31x2_ASAP7_75t_L g3965 ( 
.A1(n_3517),
.A2(n_588),
.A3(n_586),
.B(n_587),
.Y(n_3965)
);

NOR2x1_ASAP7_75t_SL g3966 ( 
.A(n_3498),
.B(n_586),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3476),
.Y(n_3967)
);

OAI21xp5_ASAP7_75t_L g3968 ( 
.A1(n_3427),
.A2(n_3450),
.B(n_3434),
.Y(n_3968)
);

AOI22xp5_ASAP7_75t_L g3969 ( 
.A1(n_3532),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_3969)
);

BUFx6f_ASAP7_75t_L g3970 ( 
.A(n_3271),
.Y(n_3970)
);

O2A1O1Ixp33_ASAP7_75t_L g3971 ( 
.A1(n_3452),
.A2(n_589),
.B(n_587),
.C(n_588),
.Y(n_3971)
);

INVx3_ASAP7_75t_L g3972 ( 
.A(n_3231),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3607),
.A2(n_589),
.B(n_590),
.Y(n_3973)
);

OAI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3455),
.A2(n_590),
.B(n_591),
.Y(n_3974)
);

AOI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_3608),
.A2(n_590),
.B(n_591),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3392),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3394),
.Y(n_3977)
);

OAI21x1_ASAP7_75t_SL g3978 ( 
.A1(n_3375),
.A2(n_591),
.B(n_592),
.Y(n_3978)
);

OAI21x1_ASAP7_75t_SL g3979 ( 
.A1(n_3178),
.A2(n_592),
.B(n_593),
.Y(n_3979)
);

OAI21xp5_ASAP7_75t_L g3980 ( 
.A1(n_3470),
.A2(n_592),
.B(n_593),
.Y(n_3980)
);

OAI21x1_ASAP7_75t_L g3981 ( 
.A1(n_3656),
.A2(n_593),
.B(n_594),
.Y(n_3981)
);

INVx3_ASAP7_75t_SL g3982 ( 
.A(n_3233),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_3609),
.A2(n_594),
.B(n_595),
.Y(n_3983)
);

A2O1A1Ixp33_ASAP7_75t_L g3984 ( 
.A1(n_3474),
.A2(n_597),
.B(n_595),
.C(n_596),
.Y(n_3984)
);

OA21x2_ASAP7_75t_L g3985 ( 
.A1(n_3173),
.A2(n_597),
.B(n_598),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3401),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3406),
.B(n_3409),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3402),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3227),
.B(n_598),
.Y(n_3989)
);

NOR2xp33_ASAP7_75t_L g3990 ( 
.A(n_3269),
.B(n_3475),
.Y(n_3990)
);

INVx2_ASAP7_75t_SL g3991 ( 
.A(n_3233),
.Y(n_3991)
);

OAI21x1_ASAP7_75t_L g3992 ( 
.A1(n_3572),
.A2(n_598),
.B(n_599),
.Y(n_3992)
);

A2O1A1Ixp33_ASAP7_75t_L g3993 ( 
.A1(n_3519),
.A2(n_601),
.B(n_599),
.C(n_600),
.Y(n_3993)
);

NAND3xp33_ASAP7_75t_L g3994 ( 
.A(n_3156),
.B(n_599),
.C(n_600),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3228),
.B(n_600),
.Y(n_3995)
);

OR2x6_ASAP7_75t_L g3996 ( 
.A(n_3498),
.B(n_601),
.Y(n_3996)
);

AO31x2_ASAP7_75t_L g3997 ( 
.A1(n_3558),
.A2(n_601),
.A3(n_602),
.B(n_640),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3326),
.B(n_602),
.Y(n_3998)
);

AOI21xp5_ASAP7_75t_L g3999 ( 
.A1(n_3630),
.A2(n_602),
.B(n_640),
.Y(n_3999)
);

OAI21x1_ASAP7_75t_L g4000 ( 
.A1(n_3524),
.A2(n_641),
.B(n_642),
.Y(n_4000)
);

AOI221x1_ASAP7_75t_L g4001 ( 
.A1(n_3344),
.A2(n_643),
.B1(n_641),
.B2(n_642),
.C(n_645),
.Y(n_4001)
);

OAI22x1_ASAP7_75t_L g4002 ( 
.A1(n_3326),
.A2(n_646),
.B1(n_643),
.B2(n_645),
.Y(n_4002)
);

AO31x2_ASAP7_75t_L g4003 ( 
.A1(n_3575),
.A2(n_649),
.A3(n_647),
.B(n_648),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3332),
.B(n_649),
.Y(n_4004)
);

NAND2x2_ASAP7_75t_L g4005 ( 
.A(n_3180),
.B(n_650),
.Y(n_4005)
);

OAI21x1_ASAP7_75t_L g4006 ( 
.A1(n_3611),
.A2(n_650),
.B(n_651),
.Y(n_4006)
);

INVx1_ASAP7_75t_SL g4007 ( 
.A(n_3181),
.Y(n_4007)
);

AOI21xp5_ASAP7_75t_L g4008 ( 
.A1(n_3631),
.A2(n_651),
.B(n_652),
.Y(n_4008)
);

AO31x2_ASAP7_75t_L g4009 ( 
.A1(n_3555),
.A2(n_654),
.A3(n_652),
.B(n_653),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3305),
.Y(n_4010)
);

AOI221xp5_ASAP7_75t_L g4011 ( 
.A1(n_3212),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.C(n_656),
.Y(n_4011)
);

OAI22xp33_ASAP7_75t_L g4012 ( 
.A1(n_3996),
.A2(n_3359),
.B1(n_3185),
.B2(n_3310),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3692),
.Y(n_4013)
);

INVx2_ASAP7_75t_L g4014 ( 
.A(n_3687),
.Y(n_4014)
);

OAI22xp5_ASAP7_75t_L g4015 ( 
.A1(n_3842),
.A2(n_3249),
.B1(n_3624),
.B2(n_3207),
.Y(n_4015)
);

INVx1_ASAP7_75t_SL g4016 ( 
.A(n_3770),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3697),
.Y(n_4017)
);

HB1xp67_ASAP7_75t_L g4018 ( 
.A(n_3804),
.Y(n_4018)
);

BUFx8_ASAP7_75t_L g4019 ( 
.A(n_3774),
.Y(n_4019)
);

AOI22xp33_ASAP7_75t_L g4020 ( 
.A1(n_3885),
.A2(n_3768),
.B1(n_3756),
.B2(n_3996),
.Y(n_4020)
);

BUFx12f_ASAP7_75t_L g4021 ( 
.A(n_3719),
.Y(n_4021)
);

INVxp67_ASAP7_75t_SL g4022 ( 
.A(n_3817),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3747),
.Y(n_4023)
);

BUFx3_ASAP7_75t_L g4024 ( 
.A(n_3781),
.Y(n_4024)
);

CKINVDCx6p67_ASAP7_75t_R g4025 ( 
.A(n_3701),
.Y(n_4025)
);

INVx4_ASAP7_75t_L g4026 ( 
.A(n_3780),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3763),
.Y(n_4027)
);

CKINVDCx16_ASAP7_75t_R g4028 ( 
.A(n_3725),
.Y(n_4028)
);

INVx3_ASAP7_75t_L g4029 ( 
.A(n_3801),
.Y(n_4029)
);

BUFx12f_ASAP7_75t_L g4030 ( 
.A(n_3963),
.Y(n_4030)
);

BUFx6f_ASAP7_75t_L g4031 ( 
.A(n_3766),
.Y(n_4031)
);

CKINVDCx5p33_ASAP7_75t_R g4032 ( 
.A(n_3757),
.Y(n_4032)
);

OAI21xp5_ASAP7_75t_SL g4033 ( 
.A1(n_3942),
.A2(n_3507),
.B(n_3648),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3771),
.Y(n_4034)
);

OAI22xp5_ASAP7_75t_L g4035 ( 
.A1(n_3842),
.A2(n_3191),
.B1(n_3591),
.B2(n_3566),
.Y(n_4035)
);

BUFx2_ASAP7_75t_L g4036 ( 
.A(n_3793),
.Y(n_4036)
);

INVx5_ASAP7_75t_L g4037 ( 
.A(n_3877),
.Y(n_4037)
);

BUFx4f_ASAP7_75t_L g4038 ( 
.A(n_3877),
.Y(n_4038)
);

OAI22xp33_ASAP7_75t_L g4039 ( 
.A1(n_3831),
.A2(n_3318),
.B1(n_3383),
.B2(n_3170),
.Y(n_4039)
);

BUFx6f_ASAP7_75t_L g4040 ( 
.A(n_3766),
.Y(n_4040)
);

INVx2_ASAP7_75t_L g4041 ( 
.A(n_3716),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3787),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3789),
.Y(n_4043)
);

BUFx4f_ASAP7_75t_SL g4044 ( 
.A(n_3686),
.Y(n_4044)
);

BUFx8_ASAP7_75t_L g4045 ( 
.A(n_3887),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_3738),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3790),
.Y(n_4047)
);

BUFx4f_ASAP7_75t_SL g4048 ( 
.A(n_3710),
.Y(n_4048)
);

OAI22xp5_ASAP7_75t_L g4049 ( 
.A1(n_3982),
.A2(n_3356),
.B1(n_3389),
.B2(n_3332),
.Y(n_4049)
);

BUFx6f_ASAP7_75t_L g4050 ( 
.A(n_3715),
.Y(n_4050)
);

BUFx12f_ASAP7_75t_L g4051 ( 
.A(n_3732),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3741),
.Y(n_4052)
);

CKINVDCx5p33_ASAP7_75t_R g4053 ( 
.A(n_3916),
.Y(n_4053)
);

INVx3_ASAP7_75t_SL g4054 ( 
.A(n_3754),
.Y(n_4054)
);

INVx2_ASAP7_75t_L g4055 ( 
.A(n_3748),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3859),
.B(n_3253),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3845),
.B(n_3292),
.Y(n_4057)
);

OAI22xp5_ASAP7_75t_L g4058 ( 
.A1(n_3711),
.A2(n_3389),
.B1(n_3356),
.B2(n_3640),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3794),
.B(n_3635),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3806),
.B(n_3639),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3795),
.Y(n_4061)
);

CKINVDCx11_ASAP7_75t_R g4062 ( 
.A(n_3784),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3826),
.B(n_3530),
.Y(n_4063)
);

AOI22xp33_ASAP7_75t_SL g4064 ( 
.A1(n_3966),
.A2(n_3236),
.B1(n_3189),
.B2(n_3194),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3830),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3785),
.Y(n_4066)
);

AOI22xp5_ASAP7_75t_L g4067 ( 
.A1(n_3834),
.A2(n_3586),
.B1(n_3617),
.B2(n_3614),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_3850),
.Y(n_4068)
);

INVx2_ASAP7_75t_L g4069 ( 
.A(n_3883),
.Y(n_4069)
);

CKINVDCx6p67_ASAP7_75t_R g4070 ( 
.A(n_3835),
.Y(n_4070)
);

OAI22xp33_ASAP7_75t_L g4071 ( 
.A1(n_3825),
.A2(n_3937),
.B1(n_4005),
.B2(n_3863),
.Y(n_4071)
);

INVx4_ASAP7_75t_SL g4072 ( 
.A(n_3825),
.Y(n_4072)
);

INVx4_ASAP7_75t_L g4073 ( 
.A(n_3788),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3864),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3867),
.Y(n_4075)
);

HB1xp67_ASAP7_75t_L g4076 ( 
.A(n_3758),
.Y(n_4076)
);

OAI22xp5_ASAP7_75t_L g4077 ( 
.A1(n_3943),
.A2(n_3492),
.B1(n_3459),
.B2(n_3194),
.Y(n_4077)
);

BUFx12f_ASAP7_75t_L g4078 ( 
.A(n_3840),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3740),
.B(n_3644),
.Y(n_4079)
);

BUFx12f_ASAP7_75t_L g4080 ( 
.A(n_3840),
.Y(n_4080)
);

INVx4_ASAP7_75t_L g4081 ( 
.A(n_3715),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_3890),
.Y(n_4082)
);

AOI22xp5_ASAP7_75t_L g4083 ( 
.A1(n_3792),
.A2(n_3633),
.B1(n_3637),
.B2(n_3396),
.Y(n_4083)
);

CKINVDCx20_ASAP7_75t_R g4084 ( 
.A(n_3708),
.Y(n_4084)
);

AOI22xp33_ASAP7_75t_L g4085 ( 
.A1(n_3720),
.A2(n_3553),
.B1(n_3261),
.B2(n_3502),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3900),
.Y(n_4086)
);

CKINVDCx6p67_ASAP7_75t_R g4087 ( 
.A(n_3858),
.Y(n_4087)
);

OAI22xp5_ASAP7_75t_L g4088 ( 
.A1(n_3717),
.A2(n_3189),
.B1(n_3565),
.B2(n_3560),
.Y(n_4088)
);

INVx3_ASAP7_75t_L g4089 ( 
.A(n_3730),
.Y(n_4089)
);

BUFx2_ASAP7_75t_L g4090 ( 
.A(n_3878),
.Y(n_4090)
);

AOI22xp33_ASAP7_75t_L g4091 ( 
.A1(n_3699),
.A2(n_3386),
.B1(n_3627),
.B2(n_3546),
.Y(n_4091)
);

AOI22xp33_ASAP7_75t_L g4092 ( 
.A1(n_3743),
.A2(n_3381),
.B1(n_3287),
.B2(n_3281),
.Y(n_4092)
);

INVx3_ASAP7_75t_L g4093 ( 
.A(n_3730),
.Y(n_4093)
);

HB1xp67_ASAP7_75t_L g4094 ( 
.A(n_3895),
.Y(n_4094)
);

INVx2_ASAP7_75t_SL g4095 ( 
.A(n_3865),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3888),
.Y(n_4096)
);

INVx2_ASAP7_75t_L g4097 ( 
.A(n_3915),
.Y(n_4097)
);

INVx8_ASAP7_75t_L g4098 ( 
.A(n_3802),
.Y(n_4098)
);

AOI22xp33_ASAP7_75t_L g4099 ( 
.A1(n_3978),
.A2(n_3541),
.B1(n_3329),
.B2(n_3251),
.Y(n_4099)
);

INVx2_ASAP7_75t_L g4100 ( 
.A(n_3921),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3855),
.Y(n_4101)
);

AOI22xp33_ASAP7_75t_L g4102 ( 
.A1(n_3696),
.A2(n_3243),
.B1(n_3367),
.B2(n_3355),
.Y(n_4102)
);

OAI22xp5_ASAP7_75t_L g4103 ( 
.A1(n_3796),
.A2(n_3565),
.B1(n_3588),
.B2(n_3560),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3934),
.Y(n_4104)
);

INVx6_ASAP7_75t_L g4105 ( 
.A(n_3744),
.Y(n_4105)
);

BUFx2_ASAP7_75t_L g4106 ( 
.A(n_3947),
.Y(n_4106)
);

BUFx4_ASAP7_75t_SL g4107 ( 
.A(n_3820),
.Y(n_4107)
);

AND2x2_ASAP7_75t_L g4108 ( 
.A(n_3761),
.B(n_3588),
.Y(n_4108)
);

INVx2_ASAP7_75t_SL g4109 ( 
.A(n_3838),
.Y(n_4109)
);

OAI22xp5_ASAP7_75t_L g4110 ( 
.A1(n_3959),
.A2(n_3644),
.B1(n_3293),
.B2(n_3275),
.Y(n_4110)
);

BUFx2_ASAP7_75t_L g4111 ( 
.A(n_3972),
.Y(n_4111)
);

CKINVDCx11_ASAP7_75t_R g4112 ( 
.A(n_3903),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_3940),
.Y(n_4113)
);

BUFx10_ASAP7_75t_L g4114 ( 
.A(n_3938),
.Y(n_4114)
);

OAI21xp33_ASAP7_75t_L g4115 ( 
.A1(n_3841),
.A2(n_3534),
.B(n_3258),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3948),
.Y(n_4116)
);

INVx6_ASAP7_75t_L g4117 ( 
.A(n_3928),
.Y(n_4117)
);

INVxp67_ASAP7_75t_SL g4118 ( 
.A(n_3870),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_3953),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3967),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3960),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3868),
.Y(n_4122)
);

BUFx8_ASAP7_75t_L g4123 ( 
.A(n_3926),
.Y(n_4123)
);

INVx6_ASAP7_75t_L g4124 ( 
.A(n_3700),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3896),
.Y(n_4125)
);

AOI22xp33_ASAP7_75t_L g4126 ( 
.A1(n_3693),
.A2(n_3705),
.B1(n_3733),
.B2(n_3951),
.Y(n_4126)
);

INVx2_ASAP7_75t_SL g4127 ( 
.A(n_3753),
.Y(n_4127)
);

BUFx10_ASAP7_75t_L g4128 ( 
.A(n_3815),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_3936),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_3958),
.Y(n_4130)
);

BUFx4f_ASAP7_75t_SL g4131 ( 
.A(n_3879),
.Y(n_4131)
);

OAI22xp5_ASAP7_75t_L g4132 ( 
.A1(n_3882),
.A2(n_3351),
.B1(n_3199),
.B2(n_3195),
.Y(n_4132)
);

AOI22xp5_ASAP7_75t_L g4133 ( 
.A1(n_3823),
.A2(n_3461),
.B1(n_3418),
.B2(n_3634),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3777),
.Y(n_4134)
);

OAI22xp33_ASAP7_75t_L g4135 ( 
.A1(n_3799),
.A2(n_3568),
.B1(n_3569),
.B2(n_3561),
.Y(n_4135)
);

AOI22xp33_ASAP7_75t_SL g4136 ( 
.A1(n_3991),
.A2(n_3182),
.B1(n_3473),
.B2(n_3672),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_3977),
.B(n_3415),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3786),
.Y(n_4138)
);

AOI22xp33_ASAP7_75t_L g4139 ( 
.A1(n_3694),
.A2(n_3680),
.B1(n_3533),
.B2(n_3465),
.Y(n_4139)
);

INVxp67_ASAP7_75t_L g4140 ( 
.A(n_3990),
.Y(n_4140)
);

CKINVDCx11_ASAP7_75t_R g4141 ( 
.A(n_4007),
.Y(n_4141)
);

INVx1_ASAP7_75t_SL g4142 ( 
.A(n_3791),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3807),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3812),
.Y(n_4144)
);

BUFx12f_ASAP7_75t_L g4145 ( 
.A(n_3722),
.Y(n_4145)
);

INVx3_ASAP7_75t_L g4146 ( 
.A(n_3713),
.Y(n_4146)
);

INVx6_ASAP7_75t_L g4147 ( 
.A(n_3878),
.Y(n_4147)
);

BUFx10_ASAP7_75t_L g4148 ( 
.A(n_3875),
.Y(n_4148)
);

HB1xp67_ASAP7_75t_L g4149 ( 
.A(n_3739),
.Y(n_4149)
);

AOI22xp33_ASAP7_75t_L g4150 ( 
.A1(n_3769),
.A2(n_3490),
.B1(n_3508),
.B2(n_3499),
.Y(n_4150)
);

AOI22xp33_ASAP7_75t_L g4151 ( 
.A1(n_3847),
.A2(n_3511),
.B1(n_3529),
.B2(n_3525),
.Y(n_4151)
);

BUFx6f_ASAP7_75t_L g4152 ( 
.A(n_3909),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_3964),
.B(n_3493),
.Y(n_4153)
);

CKINVDCx5p33_ASAP7_75t_R g4154 ( 
.A(n_3998),
.Y(n_4154)
);

BUFx2_ASAP7_75t_SL g4155 ( 
.A(n_4004),
.Y(n_4155)
);

INVx1_ASAP7_75t_SL g4156 ( 
.A(n_3857),
.Y(n_4156)
);

OAI22xp5_ASAP7_75t_L g4157 ( 
.A1(n_3950),
.A2(n_3536),
.B1(n_3625),
.B2(n_3579),
.Y(n_4157)
);

OAI22xp33_ASAP7_75t_L g4158 ( 
.A1(n_3910),
.A2(n_3642),
.B1(n_3574),
.B2(n_3549),
.Y(n_4158)
);

AOI22xp33_ASAP7_75t_L g4159 ( 
.A1(n_3848),
.A2(n_3684),
.B1(n_3559),
.B2(n_3564),
.Y(n_4159)
);

BUFx3_ASAP7_75t_L g4160 ( 
.A(n_3909),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3821),
.Y(n_4161)
);

OAI21xp5_ASAP7_75t_SL g4162 ( 
.A1(n_3837),
.A2(n_3360),
.B(n_3358),
.Y(n_4162)
);

INVx4_ASAP7_75t_L g4163 ( 
.A(n_3970),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_3986),
.B(n_3313),
.Y(n_4164)
);

BUFx3_ASAP7_75t_L g4165 ( 
.A(n_3970),
.Y(n_4165)
);

BUFx2_ASAP7_75t_SL g4166 ( 
.A(n_3893),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_SL g4167 ( 
.A(n_3939),
.B(n_3666),
.Y(n_4167)
);

BUFx3_ASAP7_75t_L g4168 ( 
.A(n_3798),
.Y(n_4168)
);

BUFx6f_ASAP7_75t_L g4169 ( 
.A(n_3703),
.Y(n_4169)
);

AOI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_3839),
.A2(n_3595),
.B1(n_3581),
.B2(n_3580),
.Y(n_4170)
);

AOI22xp33_ASAP7_75t_L g4171 ( 
.A1(n_3851),
.A2(n_3945),
.B1(n_3979),
.B2(n_3866),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3836),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_3843),
.Y(n_4173)
);

BUFx2_ASAP7_75t_SL g4174 ( 
.A(n_3712),
.Y(n_4174)
);

BUFx4_ASAP7_75t_SL g4175 ( 
.A(n_3994),
.Y(n_4175)
);

INVx6_ASAP7_75t_L g4176 ( 
.A(n_3929),
.Y(n_4176)
);

AOI22xp33_ASAP7_75t_SL g4177 ( 
.A1(n_3751),
.A2(n_3672),
.B1(n_3522),
.B2(n_3576),
.Y(n_4177)
);

OAI21xp5_ASAP7_75t_SL g4178 ( 
.A1(n_3956),
.A2(n_3241),
.B(n_3230),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3810),
.Y(n_4179)
);

INVx1_ASAP7_75t_SL g4180 ( 
.A(n_3871),
.Y(n_4180)
);

BUFx8_ASAP7_75t_L g4181 ( 
.A(n_3944),
.Y(n_4181)
);

BUFx8_ASAP7_75t_SL g4182 ( 
.A(n_3923),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3810),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_3962),
.Y(n_4184)
);

BUFx3_ASAP7_75t_L g4185 ( 
.A(n_3778),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3981),
.Y(n_4186)
);

INVx2_ASAP7_75t_SL g4187 ( 
.A(n_4002),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_3874),
.Y(n_4188)
);

AOI22xp33_ASAP7_75t_L g4189 ( 
.A1(n_3688),
.A2(n_3596),
.B1(n_3296),
.B2(n_3250),
.Y(n_4189)
);

INVx6_ASAP7_75t_L g4190 ( 
.A(n_3724),
.Y(n_4190)
);

AOI22xp33_ASAP7_75t_L g4191 ( 
.A1(n_3734),
.A2(n_3246),
.B1(n_3547),
.B2(n_3255),
.Y(n_4191)
);

INVx6_ASAP7_75t_L g4192 ( 
.A(n_3852),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_3899),
.Y(n_4193)
);

OAI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_3911),
.A2(n_3632),
.B1(n_3372),
.B2(n_3391),
.Y(n_4194)
);

BUFx12f_ASAP7_75t_L g4195 ( 
.A(n_3905),
.Y(n_4195)
);

INVx2_ASAP7_75t_SL g4196 ( 
.A(n_3904),
.Y(n_4196)
);

BUFx10_ASAP7_75t_L g4197 ( 
.A(n_3988),
.Y(n_4197)
);

BUFx12f_ASAP7_75t_L g4198 ( 
.A(n_3832),
.Y(n_4198)
);

CKINVDCx11_ASAP7_75t_R g4199 ( 
.A(n_4010),
.Y(n_4199)
);

AOI22xp33_ASAP7_75t_L g4200 ( 
.A1(n_3727),
.A2(n_3528),
.B1(n_3538),
.B2(n_3527),
.Y(n_4200)
);

AOI22xp33_ASAP7_75t_SL g4201 ( 
.A1(n_3704),
.A2(n_3661),
.B1(n_3545),
.B2(n_3666),
.Y(n_4201)
);

AND2x2_ASAP7_75t_L g4202 ( 
.A(n_3969),
.B(n_3526),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_3819),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3912),
.Y(n_4204)
);

INVx6_ASAP7_75t_L g4205 ( 
.A(n_3949),
.Y(n_4205)
);

BUFx3_ASAP7_75t_L g4206 ( 
.A(n_4000),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_3797),
.Y(n_4207)
);

OAI22xp5_ASAP7_75t_SL g4208 ( 
.A1(n_3846),
.A2(n_3330),
.B1(n_3334),
.B2(n_3324),
.Y(n_4208)
);

INVx3_ASAP7_75t_L g4209 ( 
.A(n_4006),
.Y(n_4209)
);

AOI22xp33_ASAP7_75t_L g4210 ( 
.A1(n_3861),
.A2(n_3585),
.B1(n_3610),
.B2(n_3571),
.Y(n_4210)
);

AND2x2_ASAP7_75t_L g4211 ( 
.A(n_3913),
.B(n_3535),
.Y(n_4211)
);

INVx3_ASAP7_75t_L g4212 ( 
.A(n_3813),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_3914),
.Y(n_4213)
);

AOI22xp33_ASAP7_75t_L g4214 ( 
.A1(n_3952),
.A2(n_3613),
.B1(n_3621),
.B2(n_3618),
.Y(n_4214)
);

AOI22xp33_ASAP7_75t_SL g4215 ( 
.A1(n_3918),
.A2(n_3666),
.B1(n_3616),
.B2(n_3598),
.Y(n_4215)
);

OAI22x1_ASAP7_75t_L g4216 ( 
.A1(n_3853),
.A2(n_3369),
.B1(n_3616),
.B2(n_3448),
.Y(n_4216)
);

BUFx3_ASAP7_75t_L g4217 ( 
.A(n_3814),
.Y(n_4217)
);

BUFx3_ASAP7_75t_L g4218 ( 
.A(n_3869),
.Y(n_4218)
);

OAI22xp33_ASAP7_75t_L g4219 ( 
.A1(n_3955),
.A2(n_3337),
.B1(n_3556),
.B2(n_3552),
.Y(n_4219)
);

BUFx10_ASAP7_75t_L g4220 ( 
.A(n_3961),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_4014),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4013),
.Y(n_4222)
);

OR2x2_ASAP7_75t_L g4223 ( 
.A(n_4149),
.B(n_3976),
.Y(n_4223)
);

CKINVDCx20_ASAP7_75t_R g4224 ( 
.A(n_4044),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4017),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_4156),
.B(n_4009),
.Y(n_4226)
);

AOI21x1_ASAP7_75t_L g4227 ( 
.A1(n_4216),
.A2(n_3695),
.B(n_3721),
.Y(n_4227)
);

INVx6_ASAP7_75t_L g4228 ( 
.A(n_4026),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4023),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4027),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4034),
.Y(n_4231)
);

AND2x2_ASAP7_75t_L g4232 ( 
.A(n_4168),
.B(n_4009),
.Y(n_4232)
);

INVx2_ASAP7_75t_L g4233 ( 
.A(n_4041),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4042),
.Y(n_4234)
);

INVx2_ASAP7_75t_SL g4235 ( 
.A(n_4107),
.Y(n_4235)
);

HB1xp67_ASAP7_75t_L g4236 ( 
.A(n_4036),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_4046),
.Y(n_4237)
);

BUFx3_ASAP7_75t_L g4238 ( 
.A(n_4024),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_4052),
.Y(n_4239)
);

OAI21xp33_ASAP7_75t_SL g4240 ( 
.A1(n_4020),
.A2(n_3889),
.B(n_3876),
.Y(n_4240)
);

INVxp33_ASAP7_75t_L g4241 ( 
.A(n_4038),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_4079),
.B(n_3944),
.Y(n_4242)
);

INVx2_ASAP7_75t_L g4243 ( 
.A(n_4055),
.Y(n_4243)
);

OAI21x1_ASAP7_75t_L g4244 ( 
.A1(n_4209),
.A2(n_3828),
.B(n_3736),
.Y(n_4244)
);

OAI21x1_ASAP7_75t_L g4245 ( 
.A1(n_4212),
.A2(n_3723),
.B(n_3690),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4043),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4047),
.Y(n_4247)
);

INVx1_ASAP7_75t_SL g4248 ( 
.A(n_4106),
.Y(n_4248)
);

BUFx3_ASAP7_75t_L g4249 ( 
.A(n_4048),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4061),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_4108),
.B(n_3997),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4065),
.Y(n_4252)
);

CKINVDCx12_ASAP7_75t_R g4253 ( 
.A(n_4019),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4074),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4075),
.Y(n_4255)
);

INVx2_ASAP7_75t_L g4256 ( 
.A(n_4068),
.Y(n_4256)
);

INVx2_ASAP7_75t_L g4257 ( 
.A(n_4069),
.Y(n_4257)
);

INVx2_ASAP7_75t_L g4258 ( 
.A(n_4082),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_4086),
.Y(n_4259)
);

BUFx6f_ASAP7_75t_L g4260 ( 
.A(n_4050),
.Y(n_4260)
);

INVxp67_ASAP7_75t_L g4261 ( 
.A(n_4166),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4096),
.Y(n_4262)
);

OA21x2_ASAP7_75t_L g4263 ( 
.A1(n_4179),
.A2(n_4001),
.B(n_3742),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_4097),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4183),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_4101),
.Y(n_4266)
);

AND2x2_ASAP7_75t_L g4267 ( 
.A(n_4036),
.B(n_3997),
.Y(n_4267)
);

INVx2_ASAP7_75t_L g4268 ( 
.A(n_4100),
.Y(n_4268)
);

OAI21x1_ASAP7_75t_L g4269 ( 
.A1(n_4207),
.A2(n_3702),
.B(n_3808),
.Y(n_4269)
);

AND2x2_ASAP7_75t_L g4270 ( 
.A(n_4153),
.B(n_3827),
.Y(n_4270)
);

BUFx3_ASAP7_75t_L g4271 ( 
.A(n_4031),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4104),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_4066),
.B(n_3919),
.Y(n_4273)
);

AOI22xp5_ASAP7_75t_L g4274 ( 
.A1(n_4015),
.A2(n_3706),
.B1(n_3987),
.B2(n_4011),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4121),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_4018),
.B(n_3827),
.Y(n_4276)
);

INVxp67_ASAP7_75t_SL g4277 ( 
.A(n_4118),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4094),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4076),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_4113),
.Y(n_4280)
);

OAI21x1_ASAP7_75t_L g4281 ( 
.A1(n_4129),
.A2(n_3760),
.B(n_3759),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_4134),
.B(n_3886),
.Y(n_4282)
);

INVx2_ASAP7_75t_L g4283 ( 
.A(n_4116),
.Y(n_4283)
);

BUFx2_ASAP7_75t_L g4284 ( 
.A(n_4169),
.Y(n_4284)
);

BUFx3_ASAP7_75t_L g4285 ( 
.A(n_4031),
.Y(n_4285)
);

AND2x4_ASAP7_75t_L g4286 ( 
.A(n_4072),
.B(n_3728),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_4119),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4120),
.Y(n_4288)
);

INVx2_ASAP7_75t_L g4289 ( 
.A(n_4056),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4063),
.Y(n_4290)
);

OAI21xp5_ASAP7_75t_L g4291 ( 
.A1(n_4033),
.A2(n_3745),
.B(n_3844),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4122),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4125),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4203),
.Y(n_4294)
);

INVx2_ASAP7_75t_L g4295 ( 
.A(n_4090),
.Y(n_4295)
);

BUFx3_ASAP7_75t_L g4296 ( 
.A(n_4040),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4057),
.Y(n_4297)
);

OR2x2_ASAP7_75t_L g4298 ( 
.A(n_4142),
.B(n_3989),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4197),
.Y(n_4299)
);

OAI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_4064),
.A2(n_4071),
.B(n_4039),
.Y(n_4300)
);

OAI21x1_ASAP7_75t_L g4301 ( 
.A1(n_4130),
.A2(n_3750),
.B(n_3856),
.Y(n_4301)
);

AO21x2_ASAP7_75t_L g4302 ( 
.A1(n_4167),
.A2(n_3901),
.B(n_3729),
.Y(n_4302)
);

BUFx6f_ASAP7_75t_L g4303 ( 
.A(n_4050),
.Y(n_4303)
);

BUFx6f_ASAP7_75t_L g4304 ( 
.A(n_4105),
.Y(n_4304)
);

BUFx6f_ASAP7_75t_L g4305 ( 
.A(n_4105),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4220),
.Y(n_4306)
);

AND2x2_ASAP7_75t_L g4307 ( 
.A(n_4176),
.B(n_3886),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_4090),
.Y(n_4308)
);

OAI21x1_ASAP7_75t_L g4309 ( 
.A1(n_4184),
.A2(n_3920),
.B(n_3992),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4190),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4186),
.Y(n_4311)
);

INVx3_ASAP7_75t_SL g4312 ( 
.A(n_4070),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_4211),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_4152),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4190),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4059),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4060),
.Y(n_4317)
);

INVx4_ASAP7_75t_L g4318 ( 
.A(n_4037),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4188),
.Y(n_4319)
);

OAI21x1_ASAP7_75t_L g4320 ( 
.A1(n_4110),
.A2(n_3755),
.B(n_3906),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4152),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_4160),
.Y(n_4322)
);

BUFx2_ASAP7_75t_L g4323 ( 
.A(n_4169),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_4165),
.Y(n_4324)
);

INVx3_ASAP7_75t_L g4325 ( 
.A(n_4029),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_4193),
.B(n_3749),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4204),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_4147),
.Y(n_4328)
);

BUFx6f_ASAP7_75t_L g4329 ( 
.A(n_4040),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4213),
.Y(n_4330)
);

INVx1_ASAP7_75t_SL g4331 ( 
.A(n_4054),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4138),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4147),
.Y(n_4333)
);

INVx3_ASAP7_75t_L g4334 ( 
.A(n_4163),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4111),
.Y(n_4335)
);

BUFx3_ASAP7_75t_L g4336 ( 
.A(n_4045),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4176),
.B(n_4155),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4143),
.Y(n_4338)
);

INVx2_ASAP7_75t_SL g4339 ( 
.A(n_4114),
.Y(n_4339)
);

AND2x4_ASAP7_75t_L g4340 ( 
.A(n_4072),
.B(n_3728),
.Y(n_4340)
);

INVx2_ASAP7_75t_L g4341 ( 
.A(n_4144),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4161),
.Y(n_4342)
);

INVx3_ASAP7_75t_L g4343 ( 
.A(n_4081),
.Y(n_4343)
);

OAI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_4126),
.A2(n_3809),
.B(n_4008),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4172),
.Y(n_4345)
);

BUFx6f_ASAP7_75t_L g4346 ( 
.A(n_4124),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4173),
.Y(n_4347)
);

HB1xp67_ASAP7_75t_L g4348 ( 
.A(n_4127),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4187),
.Y(n_4349)
);

CKINVDCx6p67_ASAP7_75t_R g4350 ( 
.A(n_4021),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4137),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4164),
.Y(n_4352)
);

OA21x2_ASAP7_75t_L g4353 ( 
.A1(n_4092),
.A2(n_3737),
.B(n_3726),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4196),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_L g4355 ( 
.A(n_4180),
.B(n_3933),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4022),
.Y(n_4356)
);

BUFx6f_ASAP7_75t_L g4357 ( 
.A(n_4124),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4217),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4140),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4181),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4146),
.Y(n_4361)
);

BUFx2_ASAP7_75t_L g4362 ( 
.A(n_4185),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4206),
.Y(n_4363)
);

O2A1O1Ixp33_ASAP7_75t_L g4364 ( 
.A1(n_4300),
.A2(n_4012),
.B(n_4035),
.C(n_4049),
.Y(n_4364)
);

BUFx3_ASAP7_75t_L g4365 ( 
.A(n_4224),
.Y(n_4365)
);

OA21x2_ASAP7_75t_L g4366 ( 
.A1(n_4244),
.A2(n_4178),
.B(n_4171),
.Y(n_4366)
);

OAI21x1_ASAP7_75t_L g4367 ( 
.A1(n_4227),
.A2(n_4245),
.B(n_4301),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4222),
.Y(n_4368)
);

NOR2xp33_ASAP7_75t_L g4369 ( 
.A(n_4331),
.B(n_4241),
.Y(n_4369)
);

NOR2xp33_ASAP7_75t_L g4370 ( 
.A(n_4238),
.B(n_4199),
.Y(n_4370)
);

AND2x4_ASAP7_75t_L g4371 ( 
.A(n_4235),
.B(n_4037),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4225),
.Y(n_4372)
);

OAI21xp5_ASAP7_75t_L g4373 ( 
.A1(n_4291),
.A2(n_4037),
.B(n_4088),
.Y(n_4373)
);

A2O1A1Ixp33_ASAP7_75t_L g4374 ( 
.A1(n_4261),
.A2(n_4098),
.B(n_4058),
.C(n_4109),
.Y(n_4374)
);

INVx4_ASAP7_75t_SL g4375 ( 
.A(n_4312),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4229),
.Y(n_4376)
);

OAI21x1_ASAP7_75t_L g4377 ( 
.A1(n_4227),
.A2(n_4103),
.B(n_3935),
.Y(n_4377)
);

OA21x2_ASAP7_75t_L g4378 ( 
.A1(n_4281),
.A2(n_4150),
.B(n_4162),
.Y(n_4378)
);

OR2x2_ASAP7_75t_L g4379 ( 
.A(n_4297),
.B(n_4016),
.Y(n_4379)
);

AND2x4_ASAP7_75t_L g4380 ( 
.A(n_4277),
.B(n_4089),
.Y(n_4380)
);

AND2x4_ASAP7_75t_L g4381 ( 
.A(n_4248),
.B(n_4093),
.Y(n_4381)
);

AND2x4_ASAP7_75t_L g4382 ( 
.A(n_4337),
.B(n_4084),
.Y(n_4382)
);

OR2x2_ASAP7_75t_L g4383 ( 
.A(n_4313),
.B(n_4174),
.Y(n_4383)
);

AND2x4_ASAP7_75t_L g4384 ( 
.A(n_4343),
.B(n_4095),
.Y(n_4384)
);

O2A1O1Ixp33_ASAP7_75t_SL g4385 ( 
.A1(n_4360),
.A2(n_4158),
.B(n_4135),
.C(n_4145),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4221),
.Y(n_4386)
);

OR2x6_ASAP7_75t_L g4387 ( 
.A(n_4228),
.B(n_4098),
.Y(n_4387)
);

OAI22xp33_ASAP7_75t_L g4388 ( 
.A1(n_4228),
.A2(n_4198),
.B1(n_4131),
.B2(n_4083),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_4310),
.B(n_4192),
.Y(n_4389)
);

NOR2xp33_ASAP7_75t_L g4390 ( 
.A(n_4339),
.B(n_4182),
.Y(n_4390)
);

INVx4_ASAP7_75t_L g4391 ( 
.A(n_4249),
.Y(n_4391)
);

AND2x2_ASAP7_75t_L g4392 ( 
.A(n_4315),
.B(n_4192),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4233),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_L g4394 ( 
.A(n_4316),
.B(n_4115),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4230),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4349),
.B(n_4154),
.Y(n_4396)
);

A2O1A1Ixp33_ASAP7_75t_L g4397 ( 
.A1(n_4343),
.A2(n_3946),
.B(n_3971),
.C(n_3894),
.Y(n_4397)
);

INVx2_ASAP7_75t_L g4398 ( 
.A(n_4237),
.Y(n_4398)
);

AOI22xp5_ASAP7_75t_L g4399 ( 
.A1(n_4274),
.A2(n_4208),
.B1(n_4170),
.B2(n_4077),
.Y(n_4399)
);

BUFx3_ASAP7_75t_L g4400 ( 
.A(n_4336),
.Y(n_4400)
);

INVx3_ASAP7_75t_L g4401 ( 
.A(n_4304),
.Y(n_4401)
);

OAI21xp5_ASAP7_75t_L g4402 ( 
.A1(n_4344),
.A2(n_4215),
.B(n_4136),
.Y(n_4402)
);

OAI22xp5_ASAP7_75t_SL g4403 ( 
.A1(n_4253),
.A2(n_4030),
.B1(n_4028),
.B2(n_4078),
.Y(n_4403)
);

AND2x2_ASAP7_75t_L g4404 ( 
.A(n_4278),
.B(n_4148),
.Y(n_4404)
);

INVx2_ASAP7_75t_L g4405 ( 
.A(n_4239),
.Y(n_4405)
);

OA21x2_ASAP7_75t_L g4406 ( 
.A1(n_4269),
.A2(n_4189),
.B(n_3735),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_4279),
.B(n_4128),
.Y(n_4407)
);

OR2x2_ASAP7_75t_L g4408 ( 
.A(n_4236),
.B(n_3709),
.Y(n_4408)
);

AND2x4_ASAP7_75t_L g4409 ( 
.A(n_4334),
.B(n_4073),
.Y(n_4409)
);

INVx4_ASAP7_75t_L g4410 ( 
.A(n_4304),
.Y(n_4410)
);

NAND4xp25_ASAP7_75t_SL g4411 ( 
.A(n_4240),
.B(n_4201),
.C(n_4067),
.D(n_4099),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4231),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4234),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4335),
.B(n_4218),
.Y(n_4414)
);

INVx3_ASAP7_75t_L g4415 ( 
.A(n_4304),
.Y(n_4415)
);

AND2x4_ASAP7_75t_L g4416 ( 
.A(n_4334),
.B(n_4053),
.Y(n_4416)
);

AND2x4_ASAP7_75t_L g4417 ( 
.A(n_4305),
.B(n_4032),
.Y(n_4417)
);

INVx2_ASAP7_75t_SL g4418 ( 
.A(n_4305),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4246),
.Y(n_4419)
);

AND2x4_ASAP7_75t_L g4420 ( 
.A(n_4305),
.B(n_4202),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_4243),
.Y(n_4421)
);

INVx2_ASAP7_75t_L g4422 ( 
.A(n_4250),
.Y(n_4422)
);

INVx3_ASAP7_75t_L g4423 ( 
.A(n_4271),
.Y(n_4423)
);

AND2x2_ASAP7_75t_L g4424 ( 
.A(n_4354),
.B(n_4195),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_4256),
.Y(n_4425)
);

NOR2x1_ASAP7_75t_SL g4426 ( 
.A(n_4318),
.B(n_4080),
.Y(n_4426)
);

A2O1A1Ixp33_ASAP7_75t_L g4427 ( 
.A1(n_4325),
.A2(n_3902),
.B(n_3932),
.C(n_4133),
.Y(n_4427)
);

AO21x1_ASAP7_75t_L g4428 ( 
.A1(n_4273),
.A2(n_4219),
.B(n_4132),
.Y(n_4428)
);

INVx2_ASAP7_75t_L g4429 ( 
.A(n_4257),
.Y(n_4429)
);

OAI21xp5_ASAP7_75t_L g4430 ( 
.A1(n_4320),
.A2(n_3907),
.B(n_3818),
.Y(n_4430)
);

AOI22xp5_ASAP7_75t_L g4431 ( 
.A1(n_4251),
.A2(n_4205),
.B1(n_4091),
.B2(n_4102),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4317),
.B(n_4177),
.Y(n_4432)
);

A2O1A1Ixp33_ASAP7_75t_L g4433 ( 
.A1(n_4325),
.A2(n_3974),
.B(n_3980),
.C(n_3957),
.Y(n_4433)
);

OAI21xp5_ASAP7_75t_L g4434 ( 
.A1(n_4355),
.A2(n_4356),
.B(n_3908),
.Y(n_4434)
);

AND2x4_ASAP7_75t_L g4435 ( 
.A(n_4348),
.B(n_3606),
.Y(n_4435)
);

OR2x2_ASAP7_75t_L g4436 ( 
.A(n_4223),
.B(n_3709),
.Y(n_4436)
);

HB1xp67_ASAP7_75t_L g4437 ( 
.A(n_4258),
.Y(n_4437)
);

OR2x2_ASAP7_75t_L g4438 ( 
.A(n_4290),
.B(n_4292),
.Y(n_4438)
);

NOR2xp33_ASAP7_75t_L g4439 ( 
.A(n_4299),
.B(n_4117),
.Y(n_4439)
);

AND2x2_ASAP7_75t_L g4440 ( 
.A(n_4293),
.B(n_4205),
.Y(n_4440)
);

OAI21xp33_ASAP7_75t_L g4441 ( 
.A1(n_4359),
.A2(n_4191),
.B(n_4151),
.Y(n_4441)
);

AND2x2_ASAP7_75t_L g4442 ( 
.A(n_4295),
.B(n_4087),
.Y(n_4442)
);

AND2x2_ASAP7_75t_L g4443 ( 
.A(n_4308),
.B(n_4117),
.Y(n_4443)
);

AND2x2_ASAP7_75t_L g4444 ( 
.A(n_4270),
.B(n_3930),
.Y(n_4444)
);

AND2x4_ASAP7_75t_L g4445 ( 
.A(n_4284),
.B(n_3646),
.Y(n_4445)
);

CKINVDCx5p33_ASAP7_75t_R g4446 ( 
.A(n_4350),
.Y(n_4446)
);

O2A1O1Ixp33_ASAP7_75t_L g4447 ( 
.A1(n_4306),
.A2(n_4157),
.B(n_3931),
.C(n_3941),
.Y(n_4447)
);

AND2x2_ASAP7_75t_L g4448 ( 
.A(n_4226),
.B(n_4139),
.Y(n_4448)
);

AND2x4_ASAP7_75t_L g4449 ( 
.A(n_4284),
.B(n_3555),
.Y(n_4449)
);

OAI21xp5_ASAP7_75t_L g4450 ( 
.A1(n_4232),
.A2(n_3924),
.B(n_3922),
.Y(n_4450)
);

AND2x4_ASAP7_75t_L g4451 ( 
.A(n_4323),
.B(n_3615),
.Y(n_4451)
);

HB1xp67_ASAP7_75t_L g4452 ( 
.A(n_4437),
.Y(n_4452)
);

AND2x2_ASAP7_75t_L g4453 ( 
.A(n_4389),
.B(n_4276),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4392),
.B(n_4267),
.Y(n_4454)
);

AND2x2_ASAP7_75t_L g4455 ( 
.A(n_4448),
.B(n_4307),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_4414),
.B(n_4442),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_4394),
.B(n_4352),
.Y(n_4457)
);

AND2x2_ASAP7_75t_SL g4458 ( 
.A(n_4371),
.B(n_4410),
.Y(n_4458)
);

INVx2_ASAP7_75t_L g4459 ( 
.A(n_4386),
.Y(n_4459)
);

HB1xp67_ASAP7_75t_L g4460 ( 
.A(n_4379),
.Y(n_4460)
);

AND2x4_ASAP7_75t_SL g4461 ( 
.A(n_4387),
.B(n_4025),
.Y(n_4461)
);

INVx6_ASAP7_75t_L g4462 ( 
.A(n_4375),
.Y(n_4462)
);

INVxp67_ASAP7_75t_R g4463 ( 
.A(n_4403),
.Y(n_4463)
);

INVx2_ASAP7_75t_L g4464 ( 
.A(n_4393),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4438),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4438),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4368),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4443),
.B(n_4286),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_4372),
.Y(n_4469)
);

AND2x2_ASAP7_75t_L g4470 ( 
.A(n_4404),
.B(n_4407),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_4379),
.B(n_4286),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4382),
.B(n_4340),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_4440),
.B(n_4340),
.Y(n_4473)
);

INVx1_ASAP7_75t_SL g4474 ( 
.A(n_4400),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4376),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4395),
.Y(n_4476)
);

AND2x2_ASAP7_75t_L g4477 ( 
.A(n_4444),
.B(n_4351),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4436),
.B(n_4432),
.Y(n_4478)
);

AND2x2_ASAP7_75t_L g4479 ( 
.A(n_4396),
.B(n_4380),
.Y(n_4479)
);

AND2x2_ASAP7_75t_L g4480 ( 
.A(n_4381),
.B(n_4323),
.Y(n_4480)
);

AND2x2_ASAP7_75t_L g4481 ( 
.A(n_4424),
.B(n_4247),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4412),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4413),
.Y(n_4483)
);

AOI22xp5_ASAP7_75t_L g4484 ( 
.A1(n_4411),
.A2(n_4242),
.B1(n_4282),
.B2(n_4326),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_4436),
.B(n_4341),
.Y(n_4485)
);

AOI22xp5_ASAP7_75t_L g4486 ( 
.A1(n_4399),
.A2(n_4353),
.B1(n_4318),
.B2(n_4289),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_4398),
.Y(n_4487)
);

AND2x4_ASAP7_75t_L g4488 ( 
.A(n_4375),
.B(n_4363),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4383),
.B(n_4252),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_4419),
.B(n_4319),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4405),
.Y(n_4491)
);

NOR2x1_ASAP7_75t_L g4492 ( 
.A(n_4387),
.B(n_4285),
.Y(n_4492)
);

AND2x2_ASAP7_75t_L g4493 ( 
.A(n_4383),
.B(n_4254),
.Y(n_4493)
);

INVx1_ASAP7_75t_L g4494 ( 
.A(n_4421),
.Y(n_4494)
);

AND2x2_ASAP7_75t_L g4495 ( 
.A(n_4422),
.B(n_4255),
.Y(n_4495)
);

AND2x2_ASAP7_75t_L g4496 ( 
.A(n_4425),
.B(n_4429),
.Y(n_4496)
);

AND2x4_ASAP7_75t_L g4497 ( 
.A(n_4408),
.B(n_4362),
.Y(n_4497)
);

OAI22xp5_ASAP7_75t_L g4498 ( 
.A1(n_4374),
.A2(n_4322),
.B1(n_4324),
.B2(n_4346),
.Y(n_4498)
);

INVx2_ASAP7_75t_L g4499 ( 
.A(n_4408),
.Y(n_4499)
);

OR2x2_ASAP7_75t_L g4500 ( 
.A(n_4423),
.B(n_4262),
.Y(n_4500)
);

INVx3_ASAP7_75t_L g4501 ( 
.A(n_4384),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4420),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4434),
.Y(n_4503)
);

AND2x4_ASAP7_75t_L g4504 ( 
.A(n_4418),
.B(n_4362),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4366),
.Y(n_4505)
);

NAND2x1_ASAP7_75t_SL g4506 ( 
.A(n_4391),
.B(n_4361),
.Y(n_4506)
);

AND2x4_ASAP7_75t_L g4507 ( 
.A(n_4401),
.B(n_4358),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4428),
.Y(n_4508)
);

HB1xp67_ASAP7_75t_L g4509 ( 
.A(n_4435),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_4415),
.Y(n_4510)
);

AND2x2_ASAP7_75t_L g4511 ( 
.A(n_4439),
.B(n_4327),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_4428),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_SL g4513 ( 
.A(n_4388),
.B(n_4329),
.Y(n_4513)
);

INVx2_ASAP7_75t_L g4514 ( 
.A(n_4378),
.Y(n_4514)
);

BUFx2_ASAP7_75t_L g4515 ( 
.A(n_4409),
.Y(n_4515)
);

AOI22xp33_ASAP7_75t_L g4516 ( 
.A1(n_4402),
.A2(n_4353),
.B1(n_4358),
.B2(n_4302),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_4366),
.Y(n_4517)
);

AND2x4_ASAP7_75t_L g4518 ( 
.A(n_4426),
.B(n_4265),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4378),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4406),
.Y(n_4520)
);

AND2x4_ASAP7_75t_L g4521 ( 
.A(n_4445),
.B(n_4265),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4369),
.B(n_4330),
.Y(n_4522)
);

AND2x2_ASAP7_75t_L g4523 ( 
.A(n_4416),
.B(n_4332),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4499),
.Y(n_4524)
);

INVx2_ASAP7_75t_SL g4525 ( 
.A(n_4462),
.Y(n_4525)
);

OR2x2_ASAP7_75t_L g4526 ( 
.A(n_4452),
.B(n_4338),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_4508),
.B(n_4342),
.Y(n_4527)
);

NOR2x1p5_ASAP7_75t_L g4528 ( 
.A(n_4512),
.B(n_4446),
.Y(n_4528)
);

AND2x2_ASAP7_75t_L g4529 ( 
.A(n_4471),
.B(n_4345),
.Y(n_4529)
);

OR2x2_ASAP7_75t_L g4530 ( 
.A(n_4460),
.B(n_4347),
.Y(n_4530)
);

BUFx3_ASAP7_75t_L g4531 ( 
.A(n_4462),
.Y(n_4531)
);

AOI22xp5_ASAP7_75t_L g4532 ( 
.A1(n_4484),
.A2(n_4385),
.B1(n_4441),
.B2(n_4431),
.Y(n_4532)
);

OR2x6_ASAP7_75t_L g4533 ( 
.A(n_4506),
.B(n_4370),
.Y(n_4533)
);

INVx2_ASAP7_75t_L g4534 ( 
.A(n_4496),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4480),
.B(n_4406),
.Y(n_4535)
);

OR2x2_ASAP7_75t_L g4536 ( 
.A(n_4485),
.B(n_4266),
.Y(n_4536)
);

AND2x2_ASAP7_75t_L g4537 ( 
.A(n_4456),
.B(n_4373),
.Y(n_4537)
);

INVx4_ASAP7_75t_L g4538 ( 
.A(n_4461),
.Y(n_4538)
);

AND4x1_ASAP7_75t_L g4539 ( 
.A(n_4492),
.B(n_4364),
.C(n_4390),
.D(n_4447),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4491),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4465),
.Y(n_4541)
);

OAI221xp5_ASAP7_75t_SL g4542 ( 
.A1(n_4486),
.A2(n_4397),
.B1(n_4433),
.B2(n_4427),
.C(n_4298),
.Y(n_4542)
);

HB1xp67_ASAP7_75t_L g4543 ( 
.A(n_4515),
.Y(n_4543)
);

OAI22xp5_ASAP7_75t_L g4544 ( 
.A1(n_4458),
.A2(n_4417),
.B1(n_4296),
.B2(n_4357),
.Y(n_4544)
);

INVx2_ASAP7_75t_SL g4545 ( 
.A(n_4474),
.Y(n_4545)
);

NOR3xp33_ASAP7_75t_L g4546 ( 
.A(n_4503),
.B(n_4430),
.C(n_4450),
.Y(n_4546)
);

NAND2xp5_ASAP7_75t_L g4547 ( 
.A(n_4465),
.B(n_4272),
.Y(n_4547)
);

INVx2_ASAP7_75t_L g4548 ( 
.A(n_4459),
.Y(n_4548)
);

HB1xp67_ASAP7_75t_L g4549 ( 
.A(n_4464),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4475),
.Y(n_4550)
);

AND2x4_ASAP7_75t_L g4551 ( 
.A(n_4518),
.B(n_4275),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_4468),
.B(n_4451),
.Y(n_4552)
);

AOI221xp5_ASAP7_75t_L g4553 ( 
.A1(n_4516),
.A2(n_3854),
.B1(n_4194),
.B2(n_3927),
.C(n_3975),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4473),
.B(n_4449),
.Y(n_4554)
);

NOR2xp33_ASAP7_75t_L g4555 ( 
.A(n_4509),
.B(n_4365),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_L g4556 ( 
.A(n_4466),
.B(n_4288),
.Y(n_4556)
);

AOI22xp33_ASAP7_75t_L g4557 ( 
.A1(n_4478),
.A2(n_4477),
.B1(n_4502),
.B2(n_4501),
.Y(n_4557)
);

OAI211xp5_ASAP7_75t_L g4558 ( 
.A1(n_4513),
.A2(n_4141),
.B(n_4062),
.C(n_4112),
.Y(n_4558)
);

AND2x2_ASAP7_75t_L g4559 ( 
.A(n_4472),
.B(n_4263),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4475),
.Y(n_4560)
);

AND2x4_ASAP7_75t_L g4561 ( 
.A(n_4518),
.B(n_4259),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4476),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4491),
.Y(n_4563)
);

INVx2_ASAP7_75t_SL g4564 ( 
.A(n_4501),
.Y(n_4564)
);

INVx2_ASAP7_75t_L g4565 ( 
.A(n_4487),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4457),
.B(n_4264),
.Y(n_4566)
);

HB1xp67_ASAP7_75t_L g4567 ( 
.A(n_4494),
.Y(n_4567)
);

BUFx3_ASAP7_75t_L g4568 ( 
.A(n_4488),
.Y(n_4568)
);

OR2x2_ASAP7_75t_L g4569 ( 
.A(n_4494),
.B(n_4294),
.Y(n_4569)
);

INVx2_ASAP7_75t_L g4570 ( 
.A(n_4497),
.Y(n_4570)
);

AOI22xp5_ASAP7_75t_L g4571 ( 
.A1(n_4463),
.A2(n_4333),
.B1(n_4328),
.B2(n_4346),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4497),
.Y(n_4572)
);

INVx2_ASAP7_75t_SL g4573 ( 
.A(n_4488),
.Y(n_4573)
);

AOI31xp33_ASAP7_75t_L g4574 ( 
.A1(n_4498),
.A2(n_4123),
.A3(n_4175),
.B(n_4085),
.Y(n_4574)
);

AND2x2_ASAP7_75t_L g4575 ( 
.A(n_4454),
.B(n_4263),
.Y(n_4575)
);

BUFx2_ASAP7_75t_L g4576 ( 
.A(n_4504),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4476),
.Y(n_4577)
);

AND2x2_ASAP7_75t_L g4578 ( 
.A(n_4453),
.B(n_4268),
.Y(n_4578)
);

AND2x2_ASAP7_75t_L g4579 ( 
.A(n_4455),
.B(n_4489),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_L g4580 ( 
.A(n_4495),
.B(n_4280),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4467),
.Y(n_4581)
);

CKINVDCx5p33_ASAP7_75t_R g4582 ( 
.A(n_4470),
.Y(n_4582)
);

AND2x2_ASAP7_75t_L g4583 ( 
.A(n_4493),
.B(n_4283),
.Y(n_4583)
);

OR2x2_ASAP7_75t_L g4584 ( 
.A(n_4490),
.B(n_4287),
.Y(n_4584)
);

AO21x2_ASAP7_75t_L g4585 ( 
.A1(n_4505),
.A2(n_4367),
.B(n_4377),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4576),
.B(n_4479),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4549),
.Y(n_4587)
);

AND2x2_ASAP7_75t_L g4588 ( 
.A(n_4559),
.B(n_4523),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4546),
.B(n_4469),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4577),
.Y(n_4590)
);

BUFx3_ASAP7_75t_L g4591 ( 
.A(n_4538),
.Y(n_4591)
);

OR2x2_ASAP7_75t_L g4592 ( 
.A(n_4543),
.B(n_4500),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4537),
.B(n_4522),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4535),
.B(n_4511),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4551),
.B(n_4481),
.Y(n_4595)
);

OR2x2_ASAP7_75t_L g4596 ( 
.A(n_4536),
.B(n_4519),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4577),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_4541),
.B(n_4482),
.Y(n_4598)
);

NAND2xp33_ASAP7_75t_SL g4599 ( 
.A(n_4528),
.B(n_4521),
.Y(n_4599)
);

OR2x2_ASAP7_75t_L g4600 ( 
.A(n_4567),
.B(n_4519),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4551),
.B(n_4504),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4527),
.B(n_4483),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4575),
.B(n_4521),
.Y(n_4603)
);

NAND2x1p5_ASAP7_75t_L g4604 ( 
.A(n_4538),
.B(n_4260),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4581),
.Y(n_4605)
);

NAND2x1_ASAP7_75t_L g4606 ( 
.A(n_4533),
.B(n_4507),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4581),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4550),
.B(n_4560),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4562),
.Y(n_4609)
);

AND2x2_ASAP7_75t_L g4610 ( 
.A(n_4573),
.B(n_4514),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4570),
.B(n_4510),
.Y(n_4611)
);

INVx3_ASAP7_75t_L g4612 ( 
.A(n_4533),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_4540),
.B(n_4505),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4526),
.Y(n_4614)
);

AND2x2_ASAP7_75t_L g4615 ( 
.A(n_4572),
.B(n_4507),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4568),
.B(n_4517),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4530),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4584),
.Y(n_4618)
);

INVx2_ASAP7_75t_SL g4619 ( 
.A(n_4545),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_4540),
.B(n_4517),
.Y(n_4620)
);

INVx2_ASAP7_75t_L g4621 ( 
.A(n_4561),
.Y(n_4621)
);

AND2x4_ASAP7_75t_L g4622 ( 
.A(n_4591),
.B(n_4531),
.Y(n_4622)
);

OR2x2_ASAP7_75t_L g4623 ( 
.A(n_4589),
.B(n_4566),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4589),
.B(n_4532),
.Y(n_4624)
);

INVxp67_ASAP7_75t_L g4625 ( 
.A(n_4619),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4598),
.Y(n_4626)
);

INVx2_ASAP7_75t_SL g4627 ( 
.A(n_4604),
.Y(n_4627)
);

OR2x2_ASAP7_75t_L g4628 ( 
.A(n_4596),
.B(n_4580),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4598),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4612),
.B(n_4525),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4612),
.B(n_4571),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4608),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4608),
.Y(n_4633)
);

NAND2xp5_ASAP7_75t_L g4634 ( 
.A(n_4617),
.B(n_4614),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4618),
.Y(n_4635)
);

INVx1_ASAP7_75t_SL g4636 ( 
.A(n_4604),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4593),
.B(n_4557),
.Y(n_4637)
);

NAND2xp5_ASAP7_75t_SL g4638 ( 
.A(n_4599),
.B(n_4544),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4602),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4602),
.Y(n_4640)
);

INVxp67_ASAP7_75t_L g4641 ( 
.A(n_4592),
.Y(n_4641)
);

INVxp67_ASAP7_75t_L g4642 ( 
.A(n_4586),
.Y(n_4642)
);

HB1xp67_ASAP7_75t_L g4643 ( 
.A(n_4587),
.Y(n_4643)
);

AND2x4_ASAP7_75t_L g4644 ( 
.A(n_4606),
.B(n_4555),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_4600),
.Y(n_4645)
);

INVx1_ASAP7_75t_SL g4646 ( 
.A(n_4599),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_4603),
.B(n_4564),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4613),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_4616),
.Y(n_4649)
);

OR2x2_ASAP7_75t_L g4650 ( 
.A(n_4613),
.B(n_4620),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4620),
.Y(n_4651)
);

NAND2x1p5_ASAP7_75t_L g4652 ( 
.A(n_4601),
.B(n_4561),
.Y(n_4652)
);

INVxp67_ASAP7_75t_SL g4653 ( 
.A(n_4621),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_4605),
.Y(n_4654)
);

NAND3xp33_ASAP7_75t_L g4655 ( 
.A(n_4607),
.B(n_4542),
.C(n_4539),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4609),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4590),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4594),
.B(n_4579),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4597),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4610),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4595),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4588),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4611),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_4615),
.Y(n_4664)
);

INVx3_ASAP7_75t_L g4665 ( 
.A(n_4606),
.Y(n_4665)
);

AND2x2_ASAP7_75t_L g4666 ( 
.A(n_4612),
.B(n_4552),
.Y(n_4666)
);

AND2x2_ASAP7_75t_L g4667 ( 
.A(n_4612),
.B(n_4554),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4613),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4630),
.B(n_4529),
.Y(n_4669)
);

AND2x2_ASAP7_75t_L g4670 ( 
.A(n_4644),
.B(n_4578),
.Y(n_4670)
);

INVx1_ASAP7_75t_SL g4671 ( 
.A(n_4622),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4639),
.B(n_4547),
.Y(n_4672)
);

OR2x6_ASAP7_75t_L g4673 ( 
.A(n_4622),
.B(n_4558),
.Y(n_4673)
);

AND2x2_ASAP7_75t_L g4674 ( 
.A(n_4644),
.B(n_4582),
.Y(n_4674)
);

AND2x2_ASAP7_75t_L g4675 ( 
.A(n_4631),
.B(n_4534),
.Y(n_4675)
);

NOR2xp33_ASAP7_75t_L g4676 ( 
.A(n_4625),
.B(n_4624),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4641),
.Y(n_4677)
);

INVx2_ASAP7_75t_L g4678 ( 
.A(n_4645),
.Y(n_4678)
);

INVx2_ASAP7_75t_L g4679 ( 
.A(n_4643),
.Y(n_4679)
);

OAI31xp33_ASAP7_75t_SL g4680 ( 
.A1(n_4646),
.A2(n_4574),
.A3(n_4553),
.B(n_4520),
.Y(n_4680)
);

AND2x2_ASAP7_75t_L g4681 ( 
.A(n_4667),
.B(n_4666),
.Y(n_4681)
);

INVx1_ASAP7_75t_SL g4682 ( 
.A(n_4636),
.Y(n_4682)
);

INVxp67_ASAP7_75t_L g4683 ( 
.A(n_4655),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4652),
.B(n_4583),
.Y(n_4684)
);

AND2x2_ASAP7_75t_L g4685 ( 
.A(n_4642),
.B(n_4524),
.Y(n_4685)
);

NOR3xp33_ASAP7_75t_L g4686 ( 
.A(n_4638),
.B(n_3816),
.C(n_3805),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4640),
.B(n_4520),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4654),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4668),
.Y(n_4689)
);

NOR3xp33_ASAP7_75t_L g4690 ( 
.A(n_4665),
.B(n_3993),
.C(n_3984),
.Y(n_4690)
);

NAND3xp33_ASAP7_75t_L g4691 ( 
.A(n_4668),
.B(n_4563),
.C(n_4556),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4648),
.Y(n_4692)
);

INVx2_ASAP7_75t_SL g4693 ( 
.A(n_4665),
.Y(n_4693)
);

NOR2xp33_ASAP7_75t_L g4694 ( 
.A(n_4637),
.B(n_4051),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4634),
.Y(n_4695)
);

AND2x2_ASAP7_75t_L g4696 ( 
.A(n_4660),
.B(n_4524),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4626),
.Y(n_4697)
);

AND2x4_ASAP7_75t_L g4698 ( 
.A(n_4627),
.B(n_4653),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4629),
.Y(n_4699)
);

NAND2x1_ASAP7_75t_SL g4700 ( 
.A(n_4632),
.B(n_4563),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4651),
.Y(n_4701)
);

INVx3_ASAP7_75t_SL g4702 ( 
.A(n_4623),
.Y(n_4702)
);

OR2x2_ASAP7_75t_L g4703 ( 
.A(n_4650),
.B(n_4569),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4658),
.B(n_4662),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4647),
.B(n_4585),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4633),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4635),
.Y(n_4707)
);

NOR2xp33_ASAP7_75t_L g4708 ( 
.A(n_4661),
.B(n_4548),
.Y(n_4708)
);

NOR2xp33_ASAP7_75t_L g4709 ( 
.A(n_4664),
.B(n_4663),
.Y(n_4709)
);

AND2x2_ASAP7_75t_L g4710 ( 
.A(n_4664),
.B(n_4565),
.Y(n_4710)
);

AND2x2_ASAP7_75t_L g4711 ( 
.A(n_4649),
.B(n_4346),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4656),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4657),
.Y(n_4713)
);

OR2x2_ASAP7_75t_L g4714 ( 
.A(n_4628),
.B(n_4311),
.Y(n_4714)
);

INVx2_ASAP7_75t_L g4715 ( 
.A(n_4659),
.Y(n_4715)
);

OR2x2_ASAP7_75t_L g4716 ( 
.A(n_4650),
.B(n_4311),
.Y(n_4716)
);

HB1xp67_ASAP7_75t_L g4717 ( 
.A(n_4643),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4630),
.B(n_4357),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4683),
.B(n_4159),
.Y(n_4719)
);

OAI32xp33_ASAP7_75t_L g4720 ( 
.A1(n_4671),
.A2(n_4682),
.A3(n_4693),
.B1(n_4676),
.B2(n_4717),
.Y(n_4720)
);

O2A1O1Ixp33_ASAP7_75t_L g4721 ( 
.A1(n_4702),
.A2(n_3983),
.B(n_3973),
.C(n_3999),
.Y(n_4721)
);

A2O1A1Ixp33_ASAP7_75t_L g4722 ( 
.A1(n_4680),
.A2(n_3811),
.B(n_3829),
.C(n_3822),
.Y(n_4722)
);

OAI32xp33_ASAP7_75t_L g4723 ( 
.A1(n_4677),
.A2(n_4321),
.A3(n_4314),
.B1(n_3995),
.B2(n_4200),
.Y(n_4723)
);

AOI221xp5_ASAP7_75t_L g4724 ( 
.A1(n_4695),
.A2(n_3718),
.B1(n_3714),
.B2(n_3849),
.C(n_3833),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4679),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4685),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4678),
.Y(n_4727)
);

NAND2xp33_ASAP7_75t_SL g4728 ( 
.A(n_4700),
.B(n_4357),
.Y(n_4728)
);

AND2x2_ASAP7_75t_L g4729 ( 
.A(n_4673),
.B(n_4329),
.Y(n_4729)
);

NAND2x1p5_ASAP7_75t_L g4730 ( 
.A(n_4674),
.B(n_4329),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4673),
.B(n_4260),
.Y(n_4731)
);

O2A1O1Ixp33_ASAP7_75t_SL g4732 ( 
.A1(n_4694),
.A2(n_3746),
.B(n_3689),
.C(n_3800),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4681),
.B(n_4698),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4709),
.Y(n_4734)
);

AOI22xp5_ASAP7_75t_L g4735 ( 
.A1(n_4698),
.A2(n_4214),
.B1(n_4210),
.B2(n_3775),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4710),
.Y(n_4736)
);

AND2x2_ASAP7_75t_L g4737 ( 
.A(n_4670),
.B(n_4260),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4672),
.Y(n_4738)
);

NOR2xp33_ASAP7_75t_L g4739 ( 
.A(n_4706),
.B(n_4303),
.Y(n_4739)
);

OAI22xp5_ASAP7_75t_L g4740 ( 
.A1(n_4703),
.A2(n_4303),
.B1(n_3707),
.B2(n_3772),
.Y(n_4740)
);

AND2x4_ASAP7_75t_L g4741 ( 
.A(n_4704),
.B(n_4303),
.Y(n_4741)
);

OAI221xp5_ASAP7_75t_L g4742 ( 
.A1(n_4686),
.A2(n_4697),
.B1(n_4699),
.B2(n_4690),
.C(n_4707),
.Y(n_4742)
);

OAI21xp33_ASAP7_75t_L g4743 ( 
.A1(n_4705),
.A2(n_4701),
.B(n_4692),
.Y(n_4743)
);

INVx2_ASAP7_75t_L g4744 ( 
.A(n_4696),
.Y(n_4744)
);

INVx1_ASAP7_75t_L g4745 ( 
.A(n_4715),
.Y(n_4745)
);

OAI21xp33_ASAP7_75t_L g4746 ( 
.A1(n_4692),
.A2(n_3698),
.B(n_3783),
.Y(n_4746)
);

NOR3xp33_ASAP7_75t_L g4747 ( 
.A(n_4720),
.B(n_4742),
.C(n_4725),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4727),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4733),
.B(n_4712),
.Y(n_4749)
);

AOI221xp5_ASAP7_75t_L g4750 ( 
.A1(n_4734),
.A2(n_4701),
.B1(n_4689),
.B2(n_4713),
.C(n_4688),
.Y(n_4750)
);

OR2x2_ASAP7_75t_L g4751 ( 
.A(n_4719),
.B(n_4738),
.Y(n_4751)
);

AND2x2_ASAP7_75t_L g4752 ( 
.A(n_4729),
.B(n_4731),
.Y(n_4752)
);

OR2x2_ASAP7_75t_L g4753 ( 
.A(n_4726),
.B(n_4687),
.Y(n_4753)
);

OAI32xp33_ASAP7_75t_L g4754 ( 
.A1(n_4743),
.A2(n_4689),
.A3(n_4688),
.B1(n_4718),
.B2(n_4708),
.Y(n_4754)
);

OAI33xp33_ASAP7_75t_L g4755 ( 
.A1(n_4745),
.A2(n_4691),
.A3(n_4716),
.B1(n_4714),
.B2(n_3592),
.B3(n_3422),
.Y(n_4755)
);

HB1xp67_ASAP7_75t_L g4756 ( 
.A(n_4736),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4730),
.B(n_4741),
.Y(n_4757)
);

AOI21xp5_ASAP7_75t_L g4758 ( 
.A1(n_4739),
.A2(n_4669),
.B(n_4675),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_SL g4759 ( 
.A(n_4728),
.B(n_4711),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4744),
.B(n_4684),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4740),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4721),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4732),
.B(n_655),
.Y(n_4763)
);

NAND2xp5_ASAP7_75t_L g4764 ( 
.A(n_4741),
.B(n_656),
.Y(n_4764)
);

AOI22xp5_ASAP7_75t_L g4765 ( 
.A1(n_4735),
.A2(n_3873),
.B1(n_3954),
.B2(n_3860),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4737),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4722),
.B(n_657),
.Y(n_4767)
);

OAI221xp5_ASAP7_75t_SL g4768 ( 
.A1(n_4746),
.A2(n_3872),
.B1(n_3881),
.B2(n_3880),
.C(n_3862),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4723),
.Y(n_4769)
);

NOR2xp33_ASAP7_75t_SL g4770 ( 
.A(n_4724),
.B(n_3884),
.Y(n_4770)
);

AOI22xp5_ASAP7_75t_L g4771 ( 
.A1(n_4733),
.A2(n_3891),
.B1(n_3897),
.B2(n_3892),
.Y(n_4771)
);

AOI211xp5_ASAP7_75t_L g4772 ( 
.A1(n_4720),
.A2(n_3917),
.B(n_3623),
.C(n_3803),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4725),
.Y(n_4773)
);

OAI21xp33_ASAP7_75t_L g4774 ( 
.A1(n_4733),
.A2(n_3968),
.B(n_3779),
.Y(n_4774)
);

INVxp67_ASAP7_75t_SL g4775 ( 
.A(n_4725),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4725),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_L g4777 ( 
.A(n_4725),
.B(n_657),
.Y(n_4777)
);

AND2x2_ASAP7_75t_L g4778 ( 
.A(n_4733),
.B(n_3824),
.Y(n_4778)
);

AOI22xp5_ASAP7_75t_L g4779 ( 
.A1(n_4733),
.A2(n_3985),
.B1(n_3285),
.B2(n_3506),
.Y(n_4779)
);

AOI21xp33_ASAP7_75t_L g4780 ( 
.A1(n_4720),
.A2(n_658),
.B(n_659),
.Y(n_4780)
);

NOR3xp33_ASAP7_75t_SL g4781 ( 
.A(n_4720),
.B(n_3657),
.C(n_3643),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4725),
.Y(n_4782)
);

AOI211x1_ASAP7_75t_L g4783 ( 
.A1(n_4780),
.A2(n_3782),
.B(n_3671),
.C(n_3685),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4775),
.Y(n_4784)
);

AOI22xp5_ASAP7_75t_L g4785 ( 
.A1(n_4747),
.A2(n_3505),
.B1(n_3531),
.B2(n_3509),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4756),
.Y(n_4786)
);

OAI211xp5_ASAP7_75t_SL g4787 ( 
.A1(n_4781),
.A2(n_3659),
.B(n_3174),
.C(n_3166),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4777),
.Y(n_4788)
);

XOR2x2_ASAP7_75t_L g4789 ( 
.A(n_4751),
.B(n_658),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_SL g4790 ( 
.A(n_4769),
.B(n_3762),
.Y(n_4790)
);

INVx2_ASAP7_75t_L g4791 ( 
.A(n_4766),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_SL g4792 ( 
.A(n_4773),
.B(n_3767),
.Y(n_4792)
);

OAI21xp5_ASAP7_75t_SL g4793 ( 
.A1(n_4761),
.A2(n_3691),
.B(n_3343),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4778),
.B(n_4762),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_SL g4795 ( 
.A(n_4776),
.B(n_3273),
.Y(n_4795)
);

CKINVDCx5p33_ASAP7_75t_R g4796 ( 
.A(n_4764),
.Y(n_4796)
);

INVxp67_ASAP7_75t_L g4797 ( 
.A(n_4763),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4782),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4748),
.Y(n_4799)
);

INVxp67_ASAP7_75t_L g4800 ( 
.A(n_4767),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4749),
.Y(n_4801)
);

OAI211xp5_ASAP7_75t_L g4802 ( 
.A1(n_4754),
.A2(n_3203),
.B(n_3210),
.C(n_3193),
.Y(n_4802)
);

OAI22xp5_ASAP7_75t_L g4803 ( 
.A1(n_4760),
.A2(n_3215),
.B1(n_3272),
.B2(n_3265),
.Y(n_4803)
);

AOI211x1_ASAP7_75t_L g4804 ( 
.A1(n_4752),
.A2(n_4758),
.B(n_4759),
.C(n_4757),
.Y(n_4804)
);

INVx2_ASAP7_75t_L g4805 ( 
.A(n_4753),
.Y(n_4805)
);

INVx2_ASAP7_75t_L g4806 ( 
.A(n_4779),
.Y(n_4806)
);

INVx2_ASAP7_75t_L g4807 ( 
.A(n_4765),
.Y(n_4807)
);

INVxp67_ASAP7_75t_L g4808 ( 
.A(n_4770),
.Y(n_4808)
);

HAxp5_ASAP7_75t_SL g4809 ( 
.A(n_4772),
.B(n_3824),
.CON(n_4809),
.SN(n_4809)
);

O2A1O1Ixp5_ASAP7_75t_SL g4810 ( 
.A1(n_4750),
.A2(n_4755),
.B(n_4772),
.C(n_4774),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4771),
.Y(n_4811)
);

AOI21xp33_ASAP7_75t_L g4812 ( 
.A1(n_4768),
.A2(n_660),
.B(n_661),
.Y(n_4812)
);

AOI21xp33_ASAP7_75t_L g4813 ( 
.A1(n_4775),
.A2(n_661),
.B(n_662),
.Y(n_4813)
);

INVx2_ASAP7_75t_L g4814 ( 
.A(n_4766),
.Y(n_4814)
);

OAI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_4766),
.A2(n_3573),
.B1(n_3554),
.B2(n_3655),
.Y(n_4815)
);

AND2x2_ASAP7_75t_L g4816 ( 
.A(n_4752),
.B(n_662),
.Y(n_4816)
);

NAND2xp5_ASAP7_75t_L g4817 ( 
.A(n_4775),
.B(n_664),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4816),
.B(n_665),
.Y(n_4818)
);

AOI21xp33_ASAP7_75t_L g4819 ( 
.A1(n_4784),
.A2(n_665),
.B(n_666),
.Y(n_4819)
);

OR2x2_ASAP7_75t_L g4820 ( 
.A(n_4786),
.B(n_667),
.Y(n_4820)
);

NAND3xp33_ASAP7_75t_SL g4821 ( 
.A(n_4810),
.B(n_3336),
.C(n_3317),
.Y(n_4821)
);

OR2x2_ASAP7_75t_L g4822 ( 
.A(n_4817),
.B(n_667),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4805),
.Y(n_4823)
);

XNOR2xp5_ASAP7_75t_L g4824 ( 
.A(n_4789),
.B(n_668),
.Y(n_4824)
);

NOR3xp33_ASAP7_75t_SL g4825 ( 
.A(n_4802),
.B(n_3342),
.C(n_668),
.Y(n_4825)
);

NAND5xp2_ASAP7_75t_L g4826 ( 
.A(n_4808),
.B(n_3764),
.C(n_3773),
.D(n_3776),
.E(n_672),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4791),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_L g4828 ( 
.A(n_4804),
.B(n_669),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4814),
.Y(n_4829)
);

NOR3xp33_ASAP7_75t_L g4830 ( 
.A(n_4812),
.B(n_671),
.C(n_672),
.Y(n_4830)
);

AOI22xp5_ASAP7_75t_L g4831 ( 
.A1(n_4796),
.A2(n_3765),
.B1(n_3578),
.B2(n_3615),
.Y(n_4831)
);

INVx2_ASAP7_75t_SL g4832 ( 
.A(n_4795),
.Y(n_4832)
);

NOR3xp33_ASAP7_75t_SL g4833 ( 
.A(n_4801),
.B(n_673),
.C(n_674),
.Y(n_4833)
);

NAND3x1_ASAP7_75t_L g4834 ( 
.A(n_4798),
.B(n_3482),
.C(n_4003),
.Y(n_4834)
);

AOI211xp5_ASAP7_75t_SL g4835 ( 
.A1(n_4813),
.A2(n_675),
.B(n_673),
.C(n_674),
.Y(n_4835)
);

NAND3xp33_ASAP7_75t_L g4836 ( 
.A(n_4804),
.B(n_3615),
.C(n_3288),
.Y(n_4836)
);

AND2x2_ASAP7_75t_L g4837 ( 
.A(n_4797),
.B(n_676),
.Y(n_4837)
);

OAI22xp33_ASAP7_75t_L g4838 ( 
.A1(n_4794),
.A2(n_4807),
.B1(n_4806),
.B2(n_4800),
.Y(n_4838)
);

NAND5xp2_ASAP7_75t_L g4839 ( 
.A(n_4811),
.B(n_678),
.C(n_676),
.D(n_677),
.E(n_679),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4793),
.B(n_677),
.Y(n_4840)
);

HB1xp67_ASAP7_75t_L g4841 ( 
.A(n_4799),
.Y(n_4841)
);

AND2x2_ASAP7_75t_L g4842 ( 
.A(n_4788),
.B(n_680),
.Y(n_4842)
);

NOR2xp33_ASAP7_75t_L g4843 ( 
.A(n_4790),
.B(n_681),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4792),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4783),
.Y(n_4845)
);

OAI21xp5_ASAP7_75t_L g4846 ( 
.A1(n_4787),
.A2(n_3731),
.B(n_4309),
.Y(n_4846)
);

NAND2xp33_ASAP7_75t_SL g4847 ( 
.A(n_4809),
.B(n_3273),
.Y(n_4847)
);

AOI21xp5_ASAP7_75t_L g4848 ( 
.A1(n_4815),
.A2(n_3482),
.B(n_3578),
.Y(n_4848)
);

NAND3xp33_ASAP7_75t_L g4849 ( 
.A(n_4783),
.B(n_3288),
.C(n_3273),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4785),
.B(n_681),
.Y(n_4850)
);

NAND3xp33_ASAP7_75t_SL g4851 ( 
.A(n_4803),
.B(n_682),
.C(n_683),
.Y(n_4851)
);

AOI21xp5_ASAP7_75t_L g4852 ( 
.A1(n_4817),
.A2(n_682),
.B(n_683),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4816),
.B(n_685),
.Y(n_4853)
);

NOR2x1_ASAP7_75t_L g4854 ( 
.A(n_4784),
.B(n_686),
.Y(n_4854)
);

NAND4xp25_ASAP7_75t_L g4855 ( 
.A(n_4804),
.B(n_688),
.C(n_686),
.D(n_687),
.Y(n_4855)
);

AOI22xp5_ASAP7_75t_L g4856 ( 
.A1(n_4830),
.A2(n_3350),
.B1(n_3363),
.B2(n_3288),
.Y(n_4856)
);

NAND4xp25_ASAP7_75t_L g4857 ( 
.A(n_4855),
.B(n_689),
.C(n_687),
.D(n_688),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4823),
.Y(n_4858)
);

AOI21xp5_ASAP7_75t_SL g4859 ( 
.A1(n_4828),
.A2(n_689),
.B(n_690),
.Y(n_4859)
);

OAI211xp5_ASAP7_75t_SL g4860 ( 
.A1(n_4838),
.A2(n_692),
.B(n_690),
.C(n_691),
.Y(n_4860)
);

O2A1O1Ixp33_ASAP7_75t_SL g4861 ( 
.A1(n_4827),
.A2(n_695),
.B(n_691),
.C(n_693),
.Y(n_4861)
);

AO22x2_ASAP7_75t_L g4862 ( 
.A1(n_4829),
.A2(n_4003),
.B1(n_696),
.B2(n_693),
.Y(n_4862)
);

AOI211xp5_ASAP7_75t_L g4863 ( 
.A1(n_4821),
.A2(n_697),
.B(n_695),
.C(n_696),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4820),
.Y(n_4864)
);

O2A1O1Ixp33_ASAP7_75t_L g4865 ( 
.A1(n_4840),
.A2(n_700),
.B(n_698),
.C(n_699),
.Y(n_4865)
);

NAND3xp33_ASAP7_75t_SL g4866 ( 
.A(n_4835),
.B(n_698),
.C(n_700),
.Y(n_4866)
);

OAI221xp5_ASAP7_75t_L g4867 ( 
.A1(n_4825),
.A2(n_704),
.B1(n_701),
.B2(n_702),
.C(n_706),
.Y(n_4867)
);

OAI211xp5_ASAP7_75t_L g4868 ( 
.A1(n_4851),
.A2(n_704),
.B(n_701),
.C(n_702),
.Y(n_4868)
);

OAI211xp5_ASAP7_75t_L g4869 ( 
.A1(n_4841),
.A2(n_709),
.B(n_707),
.C(n_708),
.Y(n_4869)
);

AOI22xp5_ASAP7_75t_L g4870 ( 
.A1(n_4847),
.A2(n_3363),
.B1(n_3379),
.B2(n_3350),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4824),
.B(n_708),
.Y(n_4871)
);

AOI221xp5_ASAP7_75t_L g4872 ( 
.A1(n_4832),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.C(n_713),
.Y(n_4872)
);

OAI21xp5_ASAP7_75t_L g4873 ( 
.A1(n_4836),
.A2(n_710),
.B(n_711),
.Y(n_4873)
);

AOI221xp5_ASAP7_75t_L g4874 ( 
.A1(n_4844),
.A2(n_715),
.B1(n_712),
.B2(n_714),
.C(n_716),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4837),
.B(n_714),
.Y(n_4875)
);

AOI21xp33_ASAP7_75t_L g4876 ( 
.A1(n_4854),
.A2(n_715),
.B(n_717),
.Y(n_4876)
);

OAI211xp5_ASAP7_75t_L g4877 ( 
.A1(n_4852),
.A2(n_720),
.B(n_718),
.C(n_719),
.Y(n_4877)
);

AOI22xp5_ASAP7_75t_L g4878 ( 
.A1(n_4842),
.A2(n_3363),
.B1(n_3379),
.B2(n_3350),
.Y(n_4878)
);

AOI221xp5_ASAP7_75t_L g4879 ( 
.A1(n_4819),
.A2(n_721),
.B1(n_718),
.B2(n_719),
.C(n_722),
.Y(n_4879)
);

A2O1A1Ixp33_ASAP7_75t_L g4880 ( 
.A1(n_4865),
.A2(n_4843),
.B(n_4833),
.C(n_4850),
.Y(n_4880)
);

AOI211xp5_ASAP7_75t_L g4881 ( 
.A1(n_4868),
.A2(n_4839),
.B(n_4822),
.C(n_4818),
.Y(n_4881)
);

AOI221xp5_ASAP7_75t_L g4882 ( 
.A1(n_4876),
.A2(n_4845),
.B1(n_4853),
.B2(n_4849),
.C(n_4826),
.Y(n_4882)
);

AOI21xp33_ASAP7_75t_SL g4883 ( 
.A1(n_4871),
.A2(n_4831),
.B(n_4846),
.Y(n_4883)
);

AOI221xp5_ASAP7_75t_L g4884 ( 
.A1(n_4860),
.A2(n_4848),
.B1(n_4834),
.B2(n_3412),
.C(n_3436),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_L g4885 ( 
.A(n_4858),
.B(n_4872),
.Y(n_4885)
);

AO22x2_ASAP7_75t_L g4886 ( 
.A1(n_4864),
.A2(n_724),
.B1(n_721),
.B2(n_723),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_L g4887 ( 
.A(n_4874),
.B(n_723),
.Y(n_4887)
);

XOR2xp5_ASAP7_75t_L g4888 ( 
.A(n_4857),
.B(n_4866),
.Y(n_4888)
);

OAI221xp5_ASAP7_75t_L g4889 ( 
.A1(n_4867),
.A2(n_726),
.B1(n_724),
.B2(n_725),
.C(n_727),
.Y(n_4889)
);

NAND4xp25_ASAP7_75t_L g4890 ( 
.A(n_4863),
.B(n_729),
.C(n_726),
.D(n_728),
.Y(n_4890)
);

OAI22xp5_ASAP7_75t_L g4891 ( 
.A1(n_4875),
.A2(n_3405),
.B1(n_3412),
.B2(n_3379),
.Y(n_4891)
);

AOI22xp5_ASAP7_75t_L g4892 ( 
.A1(n_4877),
.A2(n_3412),
.B1(n_3436),
.B2(n_3405),
.Y(n_4892)
);

AOI22xp5_ASAP7_75t_L g4893 ( 
.A1(n_4879),
.A2(n_3436),
.B1(n_3405),
.B2(n_3594),
.Y(n_4893)
);

INVx2_ASAP7_75t_L g4894 ( 
.A(n_4862),
.Y(n_4894)
);

AOI22xp5_ASAP7_75t_L g4895 ( 
.A1(n_4869),
.A2(n_3594),
.B1(n_3752),
.B2(n_3898),
.Y(n_4895)
);

AOI221xp5_ASAP7_75t_L g4896 ( 
.A1(n_4859),
.A2(n_3594),
.B1(n_730),
.B2(n_728),
.C(n_729),
.Y(n_4896)
);

OAI211xp5_ASAP7_75t_L g4897 ( 
.A1(n_4873),
.A2(n_733),
.B(n_731),
.C(n_732),
.Y(n_4897)
);

NOR3xp33_ASAP7_75t_SL g4898 ( 
.A(n_4861),
.B(n_734),
.C(n_735),
.Y(n_4898)
);

O2A1O1Ixp33_ASAP7_75t_L g4899 ( 
.A1(n_4862),
.A2(n_739),
.B(n_735),
.C(n_737),
.Y(n_4899)
);

OAI22xp33_ASAP7_75t_L g4900 ( 
.A1(n_4856),
.A2(n_3752),
.B1(n_3925),
.B2(n_3898),
.Y(n_4900)
);

O2A1O1Ixp33_ASAP7_75t_L g4901 ( 
.A1(n_4870),
.A2(n_742),
.B(n_739),
.C(n_740),
.Y(n_4901)
);

AND2x4_ASAP7_75t_SL g4902 ( 
.A(n_4878),
.B(n_743),
.Y(n_4902)
);

NAND2xp5_ASAP7_75t_L g4903 ( 
.A(n_4858),
.B(n_743),
.Y(n_4903)
);

OR2x2_ASAP7_75t_L g4904 ( 
.A(n_4890),
.B(n_744),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4886),
.Y(n_4905)
);

NOR2xp33_ASAP7_75t_L g4906 ( 
.A(n_4888),
.B(n_744),
.Y(n_4906)
);

NOR2x1_ASAP7_75t_L g4907 ( 
.A(n_4903),
.B(n_745),
.Y(n_4907)
);

AND2x2_ASAP7_75t_L g4908 ( 
.A(n_4898),
.B(n_4881),
.Y(n_4908)
);

OR3x2_ASAP7_75t_L g4909 ( 
.A(n_4889),
.B(n_4897),
.C(n_4896),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_SL g4910 ( 
.A(n_4882),
.B(n_745),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4886),
.Y(n_4911)
);

AO22x2_ASAP7_75t_L g4912 ( 
.A1(n_4894),
.A2(n_748),
.B1(n_746),
.B2(n_747),
.Y(n_4912)
);

BUFx12f_ASAP7_75t_L g4913 ( 
.A(n_4880),
.Y(n_4913)
);

OAI22xp5_ASAP7_75t_L g4914 ( 
.A1(n_4885),
.A2(n_3965),
.B1(n_3925),
.B2(n_750),
.Y(n_4914)
);

NAND4xp75_ASAP7_75t_L g4915 ( 
.A(n_4887),
.B(n_750),
.C(n_747),
.D(n_749),
.Y(n_4915)
);

HB1xp67_ASAP7_75t_L g4916 ( 
.A(n_4902),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4901),
.Y(n_4917)
);

AO22x2_ASAP7_75t_L g4918 ( 
.A1(n_4883),
.A2(n_752),
.B1(n_749),
.B2(n_751),
.Y(n_4918)
);

NOR2x1_ASAP7_75t_L g4919 ( 
.A(n_4899),
.B(n_751),
.Y(n_4919)
);

OR2x2_ASAP7_75t_L g4920 ( 
.A(n_4904),
.B(n_4891),
.Y(n_4920)
);

AOI221xp5_ASAP7_75t_SL g4921 ( 
.A1(n_4910),
.A2(n_4884),
.B1(n_4900),
.B2(n_4893),
.C(n_4892),
.Y(n_4921)
);

AOI221xp5_ASAP7_75t_L g4922 ( 
.A1(n_4918),
.A2(n_4895),
.B1(n_754),
.B2(n_752),
.C(n_753),
.Y(n_4922)
);

NOR3xp33_ASAP7_75t_L g4923 ( 
.A(n_4906),
.B(n_753),
.C(n_755),
.Y(n_4923)
);

OAI22xp5_ASAP7_75t_L g4924 ( 
.A1(n_4909),
.A2(n_3965),
.B1(n_758),
.B2(n_756),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4918),
.Y(n_4925)
);

NAND3xp33_ASAP7_75t_L g4926 ( 
.A(n_4919),
.B(n_756),
.C(n_757),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_L g4927 ( 
.A(n_4905),
.B(n_757),
.Y(n_4927)
);

NAND2xp5_ASAP7_75t_L g4928 ( 
.A(n_4911),
.B(n_758),
.Y(n_4928)
);

AND2x4_ASAP7_75t_L g4929 ( 
.A(n_4916),
.B(n_4908),
.Y(n_4929)
);

AOI21xp5_ASAP7_75t_L g4930 ( 
.A1(n_4912),
.A2(n_4917),
.B(n_4907),
.Y(n_4930)
);

AND2x2_ASAP7_75t_L g4931 ( 
.A(n_4912),
.B(n_759),
.Y(n_4931)
);

NAND3xp33_ASAP7_75t_L g4932 ( 
.A(n_4914),
.B(n_760),
.C(n_762),
.Y(n_4932)
);

AOI22xp5_ASAP7_75t_L g4933 ( 
.A1(n_4929),
.A2(n_4913),
.B1(n_4915),
.B2(n_763),
.Y(n_4933)
);

INVx2_ASAP7_75t_L g4934 ( 
.A(n_4920),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4931),
.Y(n_4935)
);

AND2x2_ASAP7_75t_L g4936 ( 
.A(n_4925),
.B(n_760),
.Y(n_4936)
);

OAI221xp5_ASAP7_75t_L g4937 ( 
.A1(n_4921),
.A2(n_765),
.B1(n_762),
.B2(n_764),
.C(n_766),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_L g4938 ( 
.A(n_4930),
.B(n_765),
.Y(n_4938)
);

AOI211xp5_ASAP7_75t_L g4939 ( 
.A1(n_4926),
.A2(n_768),
.B(n_766),
.C(n_767),
.Y(n_4939)
);

OAI22xp5_ASAP7_75t_SL g4940 ( 
.A1(n_4937),
.A2(n_4927),
.B1(n_4928),
.B2(n_4932),
.Y(n_4940)
);

INVx2_ASAP7_75t_L g4941 ( 
.A(n_4934),
.Y(n_4941)
);

AO22x2_ASAP7_75t_L g4942 ( 
.A1(n_4935),
.A2(n_4923),
.B1(n_4924),
.B2(n_4922),
.Y(n_4942)
);

BUFx3_ASAP7_75t_L g4943 ( 
.A(n_4936),
.Y(n_4943)
);

AOI22xp5_ASAP7_75t_L g4944 ( 
.A1(n_4938),
.A2(n_771),
.B1(n_769),
.B2(n_770),
.Y(n_4944)
);

AO22x2_ASAP7_75t_L g4945 ( 
.A1(n_4933),
.A2(n_772),
.B1(n_769),
.B2(n_771),
.Y(n_4945)
);

AO22x2_ASAP7_75t_L g4946 ( 
.A1(n_4941),
.A2(n_4939),
.B1(n_775),
.B2(n_773),
.Y(n_4946)
);

NAND2xp5_ASAP7_75t_L g4947 ( 
.A(n_4944),
.B(n_774),
.Y(n_4947)
);

AOI22xp5_ASAP7_75t_L g4948 ( 
.A1(n_4940),
.A2(n_778),
.B1(n_776),
.B2(n_777),
.Y(n_4948)
);

OAI22xp5_ASAP7_75t_SL g4949 ( 
.A1(n_4948),
.A2(n_4943),
.B1(n_4945),
.B2(n_4942),
.Y(n_4949)
);

CKINVDCx16_ASAP7_75t_R g4950 ( 
.A(n_4947),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4949),
.Y(n_4951)
);

OAI21x1_ASAP7_75t_L g4952 ( 
.A1(n_4950),
.A2(n_4946),
.B(n_776),
.Y(n_4952)
);

OAI21x1_ASAP7_75t_L g4953 ( 
.A1(n_4949),
.A2(n_778),
.B(n_780),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_L g4954 ( 
.A(n_4951),
.B(n_782),
.Y(n_4954)
);

OAI22xp5_ASAP7_75t_L g4955 ( 
.A1(n_4952),
.A2(n_784),
.B1(n_782),
.B2(n_783),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_SL g4956 ( 
.A(n_4953),
.B(n_784),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4954),
.B(n_785),
.Y(n_4957)
);

AO21x2_ASAP7_75t_L g4958 ( 
.A1(n_4956),
.A2(n_786),
.B(n_787),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4957),
.Y(n_4959)
);

NAND2xp5_ASAP7_75t_L g4960 ( 
.A(n_4958),
.B(n_4955),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4957),
.Y(n_4961)
);

OAI221xp5_ASAP7_75t_R g4962 ( 
.A1(n_4961),
.A2(n_790),
.B1(n_786),
.B2(n_787),
.C(n_791),
.Y(n_4962)
);

AOI211xp5_ASAP7_75t_L g4963 ( 
.A1(n_4962),
.A2(n_4959),
.B(n_4960),
.C(n_794),
.Y(n_4963)
);


endmodule