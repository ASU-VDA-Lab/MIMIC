module fake_jpeg_2238_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_SL g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_71),
.Y(n_75)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_61),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_64),
.B1(n_61),
.B2(n_53),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_70),
.B1(n_54),
.B2(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_57),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_73),
.B1(n_68),
.B2(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_84),
.B1(n_49),
.B2(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_48),
.B1(n_50),
.B2(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_96),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_99),
.B1(n_102),
.B2(n_8),
.Y(n_120)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_100),
.Y(n_111)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_3),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_75),
.B(n_60),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_97),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_58),
.B1(n_52),
.B2(n_4),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_3),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_82),
.B1(n_80),
.B2(n_58),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_1),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_110),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_52),
.B(n_58),
.C(n_21),
.Y(n_113)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_116),
.B1(n_16),
.B2(n_17),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_6),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_27),
.C(n_43),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_10),
.C(n_11),
.Y(n_133)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_125),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_114),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_126),
.B(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_131),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_135),
.B1(n_141),
.B2(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_136),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_11),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_13),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_140),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_15),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_141),
.Y(n_156)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_41),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_18),
.B(n_20),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_38),
.B(n_40),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_151),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_28),
.C(n_29),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_135),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_140),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_148),
.A2(n_155),
.B1(n_159),
.B2(n_154),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_36),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_157),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_42),
.B(n_45),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_133),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_164),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_153),
.C(n_158),
.Y(n_169)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_176),
.Y(n_178)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_177),
.A2(n_163),
.B1(n_161),
.B2(n_173),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_177),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_173),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_174),
.B1(n_178),
.B2(n_152),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_168),
.CI(n_152),
.CON(n_184),
.SN(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_184),
.Y(n_186)
);


endmodule