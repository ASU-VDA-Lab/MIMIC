module fake_netlist_5_1879_n_2304 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_211, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_2304);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2304;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1360;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_2248;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_314;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_16),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_124),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_138),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_59),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_52),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_191),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_187),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_167),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_15),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_115),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_122),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_55),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_186),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_160),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_118),
.Y(n_231)
);

BUFx2_ASAP7_75t_R g232 ( 
.A(n_131),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_147),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_46),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_40),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_139),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_172),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_63),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_162),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_79),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_165),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_113),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_66),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_58),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_52),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_144),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_102),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_0),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_17),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_6),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_17),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_14),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_194),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_50),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_161),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_151),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_141),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_123),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_64),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_35),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_90),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_149),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_26),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_110),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_143),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_170),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_104),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_3),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_119),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_41),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_79),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_8),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_109),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_7),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_60),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_41),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_126),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_85),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_184),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_80),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_133),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_106),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_169),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_55),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_19),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_6),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_208),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_154),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_43),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_5),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_129),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_65),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_70),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_166),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_9),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_136),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_177),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_181),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_74),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_210),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_183),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_7),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_199),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_29),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_159),
.Y(n_306)
);

INVx4_ASAP7_75t_R g307 ( 
.A(n_125),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_9),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_76),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_13),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_28),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_148),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_204),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_32),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_117),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_13),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_193),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_47),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_76),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_81),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_5),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_142),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_46),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_11),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_38),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_201),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_3),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_45),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_28),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_49),
.Y(n_330)
);

BUFx10_ASAP7_75t_L g331 ( 
.A(n_63),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_68),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_205),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_1),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_50),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_130),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_198),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_86),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_137),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_213),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_72),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_62),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_87),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_59),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_101),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_185),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_49),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_69),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_179),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_202),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_60),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_53),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_176),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_32),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_39),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_212),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_83),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_42),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_68),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_84),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_42),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_27),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_12),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_48),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_207),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_72),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_87),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_112),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_173),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_91),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_134),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_128),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_19),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_80),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_1),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_111),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_180),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_45),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_89),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_88),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_10),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_65),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_127),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_114),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_70),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_58),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_182),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_84),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_100),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_15),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_152),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_145),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_33),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_35),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_211),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_56),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_25),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_146),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_150),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_120),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_57),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_168),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_108),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_64),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_99),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_81),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_135),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_44),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_97),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_39),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_4),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_82),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_158),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_44),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_190),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_43),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_12),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_16),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_95),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_96),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_47),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_103),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_227),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_241),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_257),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_300),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_300),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_215),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_300),
.B(n_0),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_219),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_300),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_236),
.B(n_2),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_300),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_268),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_236),
.B(n_2),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_306),
.B(n_376),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_300),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_300),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_220),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_227),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_300),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_222),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_300),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_262),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_355),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_226),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_229),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_355),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_262),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_225),
.B(n_4),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_355),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_275),
.B(n_8),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_274),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_355),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_295),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_295),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_355),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_355),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_230),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_302),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_355),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_355),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_233),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_237),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_295),
.Y(n_466)
);

BUFx2_ASAP7_75t_SL g467 ( 
.A(n_225),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_L g468 ( 
.A(n_275),
.B(n_10),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_384),
.B(n_11),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_384),
.B(n_14),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_239),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_242),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_361),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_247),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_266),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_361),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_340),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_248),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_361),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_361),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_336),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_254),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_361),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_256),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_361),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_388),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_258),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_388),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_340),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_357),
.B(n_18),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_224),
.B(n_18),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_303),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_281),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_303),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_259),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_281),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_265),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_270),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_340),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_339),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_221),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_383),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_338),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_407),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_338),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_261),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_231),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_341),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_267),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_280),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_282),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_341),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_419),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_344),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_344),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_283),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_284),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_288),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_292),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_224),
.B(n_20),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_261),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_261),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_308),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_308),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_297),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_308),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_370),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_370),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_223),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_370),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_473),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_427),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_507),
.B(n_397),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_493),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_467),
.B(n_419),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_456),
.B(n_298),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_466),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_427),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_473),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_466),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_428),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_430),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_426),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_476),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_514),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_457),
.B(n_422),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_476),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_479),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_479),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_480),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_426),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_475),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_424),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_475),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_475),
.Y(n_557)
);

INVxp67_ASAP7_75t_SL g558 ( 
.A(n_530),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_466),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_431),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_480),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_517),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_483),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_431),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_425),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_433),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_495),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_477),
.B(n_397),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_437),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_437),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_500),
.B(n_397),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_508),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_483),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_485),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_438),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_439),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_485),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_438),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_441),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_514),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_441),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_443),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_434),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_443),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_522),
.B(n_406),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_445),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_454),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_445),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_461),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_510),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_442),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_448),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_446),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_467),
.B(n_436),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_448),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_481),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_451),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_451),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_522),
.B(n_406),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_453),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_447),
.Y(n_602)
);

BUFx8_ASAP7_75t_L g603 ( 
.A(n_440),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_453),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_455),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_460),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_455),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_458),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_458),
.B(n_216),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_459),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_459),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_462),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_462),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_464),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_465),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_471),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_R g617 ( 
.A(n_472),
.B(n_474),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_523),
.B(n_406),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_579),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_579),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_547),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_533),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_556),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_556),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_538),
.B(n_490),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_556),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_538),
.B(n_478),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_579),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_538),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_583),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_556),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_556),
.Y(n_632)
);

AND3x4_ASAP7_75t_L g633 ( 
.A(n_568),
.B(n_468),
.C(n_452),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_547),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_559),
.B(n_491),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_538),
.B(n_482),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_533),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g638 ( 
.A(n_537),
.B(n_350),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_583),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_542),
.B(n_484),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_533),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_583),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_533),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_581),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_556),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_573),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_542),
.B(n_490),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_556),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_540),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_569),
.B(n_490),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_542),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_542),
.B(n_523),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_559),
.B(n_487),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_585),
.Y(n_654)
);

AO21x2_ASAP7_75t_L g655 ( 
.A1(n_537),
.A2(n_429),
.B(n_470),
.Y(n_655)
);

AND2x6_ASAP7_75t_L g656 ( 
.A(n_609),
.B(n_350),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_585),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_559),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_573),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_536),
.B(n_496),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_581),
.B(n_444),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_536),
.B(n_498),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_540),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_585),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_556),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_540),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_556),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_548),
.B(n_595),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_589),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_SL g670 ( 
.A(n_617),
.B(n_470),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_540),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_540),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_555),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_557),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_555),
.Y(n_675)
);

INVx4_ASAP7_75t_SL g676 ( 
.A(n_560),
.Y(n_676)
);

NAND2x1p5_ASAP7_75t_L g677 ( 
.A(n_609),
.B(n_228),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_548),
.B(n_350),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_586),
.B(n_524),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_609),
.B(n_350),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_566),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_589),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_589),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_540),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_596),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_591),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_595),
.B(n_499),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_592),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_596),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_557),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_569),
.B(n_511),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_557),
.Y(n_692)
);

INVxp33_ASAP7_75t_L g693 ( 
.A(n_586),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_596),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_569),
.B(n_572),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_557),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_598),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_545),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_598),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_545),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_545),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_572),
.A2(n_435),
.B1(n_432),
.B2(n_450),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_535),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_557),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_572),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_557),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_535),
.B(n_444),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_598),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_608),
.B(n_512),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_534),
.B(n_531),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_608),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_608),
.Y(n_712)
);

CKINVDCx16_ASAP7_75t_R g713 ( 
.A(n_568),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_543),
.B(n_518),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_534),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_557),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_558),
.B(n_495),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_558),
.A2(n_502),
.B1(n_469),
.B2(n_449),
.Y(n_718)
);

BUFx4f_ASAP7_75t_L g719 ( 
.A(n_560),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_545),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_534),
.Y(n_721)
);

INVx4_ASAP7_75t_SL g722 ( 
.A(n_560),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_553),
.Y(n_723)
);

AND2x6_ASAP7_75t_L g724 ( 
.A(n_609),
.B(n_350),
.Y(n_724)
);

OAI221xp5_ASAP7_75t_L g725 ( 
.A1(n_611),
.A2(n_492),
.B1(n_521),
.B2(n_491),
.C(n_429),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_609),
.A2(n_440),
.B1(n_423),
.B2(n_452),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_611),
.B(n_519),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_557),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_586),
.B(n_524),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_611),
.B(n_520),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_544),
.A2(n_577),
.B1(n_615),
.B2(n_614),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_612),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_600),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_617),
.B(n_526),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_612),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_616),
.B(n_525),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_557),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_600),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_553),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_603),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_600),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_592),
.B(n_525),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_618),
.B(n_527),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_618),
.B(n_527),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_539),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_612),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_568),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_594),
.B(n_528),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_553),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_613),
.B(n_463),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_613),
.Y(n_751)
);

BUFx4f_ASAP7_75t_L g752 ( 
.A(n_560),
.Y(n_752)
);

NAND2x1p5_ASAP7_75t_L g753 ( 
.A(n_609),
.B(n_228),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_591),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_618),
.B(n_528),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_594),
.A2(n_501),
.B1(n_505),
.B2(n_503),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_613),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_576),
.B(n_463),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_553),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_576),
.B(n_322),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_602),
.B(n_529),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_562),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_539),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_532),
.B(n_529),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_539),
.Y(n_765)
);

INVx5_ASAP7_75t_L g766 ( 
.A(n_560),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_576),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_532),
.B(n_531),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_560),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_602),
.B(n_357),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_576),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_715),
.B(n_606),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_715),
.B(n_606),
.Y(n_773)
);

AND2x2_ASAP7_75t_SL g774 ( 
.A(n_740),
.B(n_216),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_668),
.B(n_576),
.Y(n_775)
);

AND2x2_ASAP7_75t_SL g776 ( 
.A(n_740),
.B(n_313),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_670),
.A2(n_603),
.B1(n_304),
.B2(n_312),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_695),
.B(n_576),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_725),
.A2(n_468),
.B1(n_263),
.B2(n_278),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_741),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_705),
.B(n_603),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_702),
.A2(n_402),
.B1(n_313),
.B2(n_263),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_741),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_687),
.B(n_580),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_705),
.B(n_603),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_742),
.B(n_562),
.Y(n_786)
);

AO22x1_ASAP7_75t_L g787 ( 
.A1(n_633),
.A2(n_603),
.B1(n_243),
.B2(n_289),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_764),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_721),
.B(n_580),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_721),
.B(n_486),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_733),
.B(n_580),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_650),
.B(n_486),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_653),
.B(n_603),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_L g794 ( 
.A1(n_693),
.A2(n_278),
.B1(n_289),
.B2(n_243),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_619),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_619),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_650),
.A2(n_593),
.B(n_580),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_620),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_733),
.B(n_580),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_738),
.B(n_301),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_738),
.B(n_580),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_620),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_748),
.B(n_566),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_652),
.B(n_593),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_691),
.A2(n_349),
.B1(n_353),
.B2(n_326),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_710),
.A2(n_365),
.B1(n_368),
.B2(n_356),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_710),
.A2(n_377),
.B1(n_389),
.B2(n_369),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_679),
.B(n_488),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_628),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_652),
.B(n_655),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_625),
.B(n_647),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_621),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_628),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_652),
.B(n_655),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_625),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_655),
.B(n_593),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_621),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_635),
.A2(n_402),
.B1(n_315),
.B2(n_317),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_762),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_629),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_625),
.B(n_593),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_764),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_769),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_679),
.A2(n_604),
.B1(n_605),
.B2(n_593),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_761),
.B(n_584),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_629),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_768),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_647),
.B(n_593),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_661),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_647),
.B(n_604),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_689),
.B(n_694),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_709),
.A2(n_554),
.B(n_564),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_769),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_736),
.B(n_395),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_697),
.B(n_604),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_630),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_658),
.B(n_770),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_644),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_699),
.B(n_604),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_658),
.B(n_398),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_630),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_708),
.B(n_604),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_639),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_639),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_635),
.A2(n_400),
.B1(n_399),
.B2(n_299),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_717),
.B(n_345),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_727),
.B(n_604),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_730),
.A2(n_554),
.B(n_564),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_642),
.B(n_605),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_769),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_679),
.A2(n_605),
.B1(n_565),
.B2(n_567),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_729),
.B(n_299),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_651),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_729),
.A2(n_605),
.B1(n_565),
.B2(n_567),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_642),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_654),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_654),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_657),
.B(n_605),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_729),
.A2(n_605),
.B1(n_565),
.B2(n_567),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_657),
.B(n_560),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_635),
.A2(n_317),
.B1(n_333),
.B2(n_315),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_755),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_664),
.B(n_560),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_664),
.B(n_560),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_660),
.B(n_584),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_661),
.Y(n_866)
);

AOI221xp5_ASAP7_75t_L g867 ( 
.A1(n_718),
.A2(n_421),
.B1(n_311),
.B2(n_354),
.C(n_378),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_755),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_743),
.A2(n_565),
.B1(n_567),
.B2(n_564),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_669),
.B(n_570),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_743),
.B(n_333),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_R g872 ( 
.A(n_762),
.B(n_588),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_662),
.B(n_588),
.Y(n_873)
);

BUFx4f_ASAP7_75t_L g874 ( 
.A(n_677),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_717),
.B(n_345),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_669),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_651),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_635),
.A2(n_337),
.B1(n_371),
.B2(n_346),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_682),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_743),
.B(n_488),
.Y(n_880)
);

OAI21xp33_ASAP7_75t_L g881 ( 
.A1(n_726),
.A2(n_408),
.B(n_363),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_682),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_683),
.B(n_570),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_744),
.B(n_489),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_683),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_707),
.B(n_363),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_685),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_685),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_707),
.B(n_345),
.Y(n_889)
);

NAND2x1p5_ASAP7_75t_L g890 ( 
.A(n_711),
.B(n_337),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_744),
.B(n_345),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_711),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_744),
.A2(n_346),
.B1(n_372),
.B2(n_371),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_646),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_646),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_768),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_714),
.B(n_590),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_634),
.B(n_408),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_712),
.B(n_570),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_627),
.B(n_350),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_703),
.B(n_590),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_712),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_768),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_732),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_634),
.B(n_489),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_732),
.B(n_570),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_735),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_633),
.A2(n_387),
.B1(n_391),
.B2(n_372),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_636),
.A2(n_391),
.B1(n_392),
.B2(n_387),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_735),
.B(n_570),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_746),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_640),
.A2(n_403),
.B1(n_405),
.B2(n_392),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_677),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_746),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_760),
.A2(n_405),
.B1(n_413),
.B2(n_403),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_751),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_751),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_757),
.B(n_570),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_757),
.B(n_570),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_767),
.B(n_570),
.Y(n_920)
);

NAND2xp33_ASAP7_75t_SL g921 ( 
.A(n_734),
.B(n_240),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_767),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_771),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_731),
.B(n_415),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_771),
.B(n_570),
.Y(n_925)
);

NOR2xp67_ASAP7_75t_L g926 ( 
.A(n_756),
.B(n_659),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_632),
.B(n_610),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_632),
.B(n_645),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_677),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_753),
.Y(n_930)
);

BUFx8_ASAP7_75t_L g931 ( 
.A(n_713),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_673),
.B(n_597),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_675),
.B(n_597),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_753),
.B(n_532),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_698),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_747),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_681),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_719),
.A2(n_554),
.B(n_564),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_632),
.B(n_610),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_624),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_659),
.B(n_214),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_698),
.Y(n_942)
);

NOR2x2_ASAP7_75t_L g943 ( 
.A(n_747),
.B(n_232),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_638),
.A2(n_582),
.B1(n_587),
.B2(n_571),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_792),
.B(n_750),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_812),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_R g947 ( 
.A(n_819),
.B(n_686),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_792),
.B(n_758),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_784),
.A2(n_753),
.B1(n_719),
.B2(n_752),
.Y(n_949)
);

INVx5_ASAP7_75t_L g950 ( 
.A(n_823),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_812),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_809),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_817),
.Y(n_953)
);

AO221x1_ASAP7_75t_L g954 ( 
.A1(n_779),
.A2(n_366),
.B1(n_250),
.B2(n_269),
.C(n_273),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_782),
.A2(n_678),
.B1(n_638),
.B2(n_656),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_SL g956 ( 
.A(n_867),
.B(n_754),
.C(n_686),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_811),
.A2(n_678),
.B1(n_674),
.B2(n_645),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_811),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_811),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_809),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_817),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_780),
.B(n_827),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_922),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_780),
.B(n_413),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_790),
.B(n_645),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_874),
.B(n_688),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_773),
.A2(n_674),
.B1(n_765),
.B2(n_716),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_826),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_852),
.A2(n_656),
.B1(n_724),
.B2(n_680),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_826),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_931),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_838),
.Y(n_972)
);

BUFx12f_ASAP7_75t_L g973 ( 
.A(n_931),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_931),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_905),
.Y(n_975)
);

INVx5_ASAP7_75t_L g976 ( 
.A(n_823),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_SL g977 ( 
.A(n_786),
.B(n_754),
.C(n_367),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_790),
.B(n_674),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_775),
.B(n_716),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_896),
.B(n_716),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_826),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_SL g982 ( 
.A(n_921),
.B(n_218),
.C(n_217),
.Y(n_982)
);

INVxp67_ASAP7_75t_SL g983 ( 
.A(n_820),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_829),
.B(n_866),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_788),
.B(n_765),
.Y(n_985)
);

NOR3xp33_ASAP7_75t_SL g986 ( 
.A(n_921),
.B(n_235),
.C(n_234),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_905),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_822),
.B(n_917),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_SL g989 ( 
.A(n_793),
.B(n_364),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_922),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_SL g991 ( 
.A(n_819),
.B(n_244),
.C(n_238),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_903),
.B(n_765),
.Y(n_992)
);

INVx5_ASAP7_75t_L g993 ( 
.A(n_823),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_937),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_773),
.A2(n_680),
.B1(n_724),
.B2(n_656),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_923),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_923),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_783),
.B(n_649),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_795),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_826),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_941),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_803),
.B(n_688),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_940),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_826),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_778),
.A2(n_250),
.B(n_269),
.C(n_223),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_877),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_808),
.B(n_700),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_856),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_874),
.B(n_688),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_913),
.B(n_623),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_795),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_808),
.B(n_700),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_880),
.B(n_701),
.Y(n_1013)
);

BUFx4f_ASAP7_75t_L g1014 ( 
.A(n_877),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_872),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_796),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_796),
.Y(n_1017)
);

OR2x6_ASAP7_75t_L g1018 ( 
.A(n_787),
.B(n_415),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_856),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_877),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_894),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_940),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_862),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_857),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_798),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_880),
.B(n_701),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_815),
.A2(n_680),
.B1(n_724),
.B2(n_656),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_877),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_877),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_798),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_884),
.B(n_720),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_884),
.B(n_649),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_SL g1033 ( 
.A(n_894),
.B(n_246),
.C(n_245),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_L g1034 ( 
.A(n_772),
.B(n_837),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_815),
.A2(n_680),
.B1(n_724),
.B2(n_656),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_913),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_R g1037 ( 
.A(n_895),
.B(n_249),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_857),
.Y(n_1038)
);

AOI22x1_ASAP7_75t_L g1039 ( 
.A1(n_876),
.A2(n_626),
.B1(n_665),
.B2(n_623),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_802),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_874),
.B(n_624),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_833),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_895),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_862),
.B(n_720),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_802),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_833),
.Y(n_1046)
);

BUFx4f_ASAP7_75t_L g1047 ( 
.A(n_774),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_868),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_820),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_852),
.A2(n_680),
.B1(n_724),
.B2(n_656),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_868),
.B(n_813),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_876),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_813),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_852),
.B(n_663),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_836),
.B(n_723),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_787),
.B(n_415),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_936),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_871),
.B(n_723),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_836),
.B(n_739),
.Y(n_1059)
);

NAND2x1p5_ASAP7_75t_L g1060 ( 
.A(n_929),
.B(n_623),
.Y(n_1060)
);

BUFx2_ASAP7_75t_R g1061 ( 
.A(n_936),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_774),
.B(n_624),
.Y(n_1062)
);

OAI221xp5_ASAP7_75t_L g1063 ( 
.A1(n_881),
.A2(n_374),
.B1(n_366),
.B2(n_360),
.C(n_352),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_841),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_929),
.B(n_626),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_R g1066 ( 
.A(n_897),
.B(n_251),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_898),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_940),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_879),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_871),
.B(n_739),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_841),
.B(n_749),
.Y(n_1071)
);

AO22x1_ASAP7_75t_L g1072 ( 
.A1(n_865),
.A2(n_873),
.B1(n_825),
.B2(n_861),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_871),
.B(n_663),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_898),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_820),
.B(n_626),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_SL g1076 ( 
.A(n_901),
.B(n_253),
.C(n_252),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_886),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_932),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_886),
.B(n_749),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_853),
.Y(n_1080)
);

BUFx12f_ASAP7_75t_L g1081 ( 
.A(n_890),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_879),
.Y(n_1082)
);

AOI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_794),
.A2(n_342),
.B1(n_335),
.B2(n_334),
.C(n_332),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_818),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_890),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_810),
.A2(n_752),
.B1(n_719),
.B2(n_667),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_933),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_887),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_887),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_943),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_853),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_892),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_892),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_R g1094 ( 
.A(n_930),
.B(n_255),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_890),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_908),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_840),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_853),
.B(n_666),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_843),
.B(n_844),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_L g1100 ( 
.A(n_781),
.B(n_665),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_SL g1101 ( 
.A(n_846),
.B(n_264),
.C(n_260),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_776),
.B(n_624),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_777),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_843),
.B(n_759),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_833),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_844),
.B(n_759),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_902),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_855),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_R g1109 ( 
.A(n_776),
.B(n_855),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_R g1110 ( 
.A(n_882),
.B(n_271),
.Y(n_1110)
);

INVx6_ASAP7_75t_L g1111 ( 
.A(n_850),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_882),
.B(n_666),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_SL g1113 ( 
.A(n_875),
.B(n_276),
.C(n_272),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_885),
.B(n_624),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_885),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_SL g1116 ( 
.A(n_889),
.B(n_286),
.C(n_277),
.Y(n_1116)
);

NAND2xp33_ASAP7_75t_SL g1117 ( 
.A(n_785),
.B(n_415),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_888),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_888),
.B(n_622),
.Y(n_1119)
);

BUFx2_ASAP7_75t_R g1120 ( 
.A(n_891),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_914),
.B(n_631),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_845),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_914),
.B(n_671),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_SL g1124 ( 
.A(n_924),
.B(n_294),
.C(n_293),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_R g1125 ( 
.A(n_814),
.B(n_296),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_847),
.B(n_631),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_902),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_789),
.B(n_631),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_831),
.B(n_631),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_943),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_904),
.Y(n_1131)
);

OR2x6_ASAP7_75t_L g1132 ( 
.A(n_926),
.B(n_415),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_904),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_907),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_907),
.B(n_671),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_911),
.B(n_672),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_911),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_824),
.B(n_631),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1039),
.A2(n_863),
.B(n_860),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_L g1140 ( 
.A(n_956),
.B(n_805),
.C(n_806),
.Y(n_1140)
);

NAND2xp33_ASAP7_75t_L g1141 ( 
.A(n_950),
.B(n_816),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_L g1142 ( 
.A(n_1072),
.B(n_807),
.C(n_834),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1128),
.A2(n_870),
.B(n_864),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1138),
.A2(n_797),
.B(n_791),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1086),
.A2(n_899),
.B(n_883),
.Y(n_1145)
);

AOI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_1002),
.A2(n_800),
.B(n_909),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1079),
.B(n_916),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1047),
.A2(n_878),
.B(n_915),
.C(n_916),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_1126),
.A2(n_910),
.B(n_906),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_973),
.B(n_821),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1041),
.A2(n_919),
.B(n_918),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_963),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1042),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1041),
.A2(n_1075),
.B(n_979),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1075),
.A2(n_925),
.B(n_920),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1114),
.A2(n_858),
.B(n_849),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_990),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1087),
.B(n_799),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1121),
.A2(n_848),
.B(n_832),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1100),
.A2(n_939),
.B(n_927),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1079),
.B(n_801),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_SL g1162 ( 
.A1(n_1046),
.A2(n_893),
.B(n_830),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1138),
.A2(n_804),
.B(n_828),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_975),
.B(n_934),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_996),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1077),
.B(n_331),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1047),
.A2(n_851),
.B1(n_859),
.B2(n_854),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1060),
.A2(n_928),
.B(n_839),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1060),
.A2(n_842),
.B(n_835),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_975),
.B(n_934),
.Y(n_1170)
);

AOI221x1_ASAP7_75t_L g1171 ( 
.A1(n_989),
.A2(n_912),
.B1(n_938),
.B2(n_942),
.C(n_935),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1065),
.A2(n_942),
.B(n_935),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1065),
.A2(n_900),
.B(n_869),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_946),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1036),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_989),
.A2(n_1122),
.B1(n_1047),
.B2(n_987),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_997),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_950),
.A2(n_850),
.B(n_752),
.Y(n_1178)
);

NAND2x1_ASAP7_75t_L g1179 ( 
.A(n_1111),
.B(n_1042),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_999),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1055),
.A2(n_944),
.B(n_637),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_950),
.A2(n_850),
.B(n_667),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_950),
.B(n_648),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1067),
.B(n_331),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_950),
.B(n_648),
.Y(n_1185)
);

AOI21xp33_ASAP7_75t_L g1186 ( 
.A1(n_1122),
.A2(n_314),
.B(n_310),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_987),
.B(n_622),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_948),
.A2(n_641),
.B(n_637),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_947),
.Y(n_1189)
);

BUFx12f_ASAP7_75t_L g1190 ( 
.A(n_973),
.Y(n_1190)
);

NOR4xp25_ASAP7_75t_L g1191 ( 
.A(n_977),
.B(n_329),
.C(n_287),
.D(n_285),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_965),
.A2(n_643),
.B(n_641),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_946),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_SL g1194 ( 
.A1(n_1046),
.A2(n_279),
.B(n_273),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_976),
.A2(n_667),
.B(n_665),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1059),
.A2(n_643),
.B(n_672),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_945),
.B(n_648),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_976),
.A2(n_706),
.B(n_696),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1071),
.A2(n_684),
.B(n_582),
.Y(n_1199)
);

CKINVDCx8_ASAP7_75t_R g1200 ( 
.A(n_1043),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1051),
.B(n_648),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1005),
.A2(n_385),
.A3(n_386),
.B(n_401),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1043),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_976),
.A2(n_706),
.B(n_696),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_988),
.B(n_648),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1104),
.A2(n_684),
.B(n_582),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1011),
.A2(n_320),
.B(n_309),
.C(n_324),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1106),
.A2(n_582),
.B(n_571),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1129),
.A2(n_546),
.B(n_541),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_976),
.A2(n_706),
.B(n_696),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1078),
.B(n_316),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_976),
.A2(n_745),
.B(n_728),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_949),
.A2(n_587),
.B(n_571),
.Y(n_1213)
);

INVxp67_ASAP7_75t_SL g1214 ( 
.A(n_1042),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1016),
.A2(n_324),
.B(n_320),
.C(n_309),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_993),
.A2(n_745),
.B(n_728),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1099),
.B(n_690),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1078),
.B(n_318),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1046),
.A2(n_285),
.B(n_279),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_958),
.B(n_728),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_1042),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1099),
.B(n_690),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1069),
.A2(n_587),
.B(n_571),
.Y(n_1223)
);

NOR3xp33_ASAP7_75t_L g1224 ( 
.A(n_1090),
.B(n_321),
.C(n_319),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1099),
.B(n_690),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1042),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1017),
.A2(n_291),
.B(n_290),
.C(n_287),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1025),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1115),
.B(n_690),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_978),
.A2(n_1012),
.B(n_1007),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1115),
.B(n_690),
.Y(n_1231)
);

AO32x2_ASAP7_75t_L g1232 ( 
.A1(n_970),
.A2(n_763),
.A3(n_745),
.B1(n_329),
.B2(n_334),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1074),
.B(n_972),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1118),
.A2(n_763),
.B1(n_737),
.B2(n_704),
.Y(n_1234)
);

OAI21xp33_ASAP7_75t_L g1235 ( 
.A1(n_1066),
.A2(n_325),
.B(n_323),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_993),
.A2(n_763),
.B(n_737),
.Y(n_1236)
);

AO32x2_ASAP7_75t_L g1237 ( 
.A1(n_970),
.A2(n_360),
.A3(n_332),
.B1(n_335),
.B2(n_416),
.Y(n_1237)
);

NOR4xp25_ASAP7_75t_L g1238 ( 
.A(n_1005),
.B(n_416),
.C(n_414),
.D(n_411),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1069),
.A2(n_599),
.B(n_587),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_993),
.A2(n_737),
.B(n_704),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1119),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1013),
.A2(n_680),
.B(n_656),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1118),
.A2(n_737),
.B1(n_704),
.B2(n_769),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1030),
.A2(n_291),
.A3(n_290),
.B(n_305),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1040),
.B(n_704),
.Y(n_1245)
);

OAI22x1_ASAP7_75t_L g1246 ( 
.A1(n_1096),
.A2(n_390),
.B1(n_328),
.B2(n_330),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1045),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1105),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1053),
.B(n_704),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1069),
.A2(n_601),
.B(n_599),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1089),
.A2(n_601),
.B(n_599),
.Y(n_1251)
);

NAND2x1_ASAP7_75t_L g1252 ( 
.A(n_1111),
.B(n_737),
.Y(n_1252)
);

AND3x2_ASAP7_75t_L g1253 ( 
.A(n_994),
.B(n_342),
.C(n_305),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1089),
.A2(n_601),
.B(n_599),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1064),
.B(n_769),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_958),
.B(n_962),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1089),
.A2(n_607),
.B(n_601),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1108),
.B(n_607),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_994),
.B(n_331),
.Y(n_1259)
);

OA22x2_ASAP7_75t_L g1260 ( 
.A1(n_1096),
.A2(n_374),
.B1(n_418),
.B2(n_352),
.Y(n_1260)
);

AOI21xp33_ASAP7_75t_L g1261 ( 
.A1(n_984),
.A2(n_343),
.B(n_327),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1001),
.B(n_331),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1093),
.A2(n_607),
.B(n_546),
.Y(n_1263)
);

AOI211x1_ASAP7_75t_L g1264 ( 
.A1(n_1063),
.A2(n_418),
.B(n_414),
.C(n_385),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1001),
.B(n_375),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1026),
.A2(n_724),
.B(n_680),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_962),
.B(n_607),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_951),
.B(n_347),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1001),
.B(n_375),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_961),
.B(n_375),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_952),
.A2(n_386),
.A3(n_411),
.B(n_401),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1021),
.B(n_494),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1083),
.A2(n_420),
.B(n_417),
.C(n_348),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1062),
.A2(n_549),
.B(n_541),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1031),
.A2(n_724),
.B(n_549),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1093),
.A2(n_549),
.B(n_541),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1093),
.A2(n_550),
.B(n_546),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_SL g1278 ( 
.A1(n_1105),
.A2(n_539),
.B(n_415),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_953),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_993),
.A2(n_1014),
.B(n_1105),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_993),
.A2(n_692),
.B(n_554),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_953),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1034),
.A2(n_1097),
.B1(n_1103),
.B2(n_962),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1044),
.B(n_550),
.Y(n_1284)
);

OA22x2_ASAP7_75t_L g1285 ( 
.A1(n_961),
.A2(n_393),
.B1(n_382),
.B2(n_381),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_967),
.A2(n_551),
.B(n_550),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1014),
.A2(n_692),
.B(n_554),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1023),
.B(n_375),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1062),
.A2(n_1102),
.B(n_985),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1014),
.A2(n_692),
.B(n_554),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1057),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_952),
.A2(n_575),
.A3(n_574),
.B(n_563),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1111),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_954),
.A2(n_266),
.B1(n_351),
.B2(n_358),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1102),
.A2(n_551),
.B(n_552),
.Y(n_1295)
);

NOR2x1_ASAP7_75t_L g1296 ( 
.A(n_958),
.B(n_551),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_966),
.B(n_98),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1107),
.A2(n_561),
.B(n_552),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1107),
.A2(n_561),
.B(n_552),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1084),
.A2(n_1036),
.B1(n_1111),
.B2(n_1085),
.Y(n_1300)
);

AOI31xp67_ASAP7_75t_L g1301 ( 
.A1(n_960),
.A2(n_722),
.A3(n_676),
.B(n_266),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1057),
.B(n_1048),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1048),
.B(n_494),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1049),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_983),
.A2(n_692),
.B(n_766),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_964),
.B(n_497),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1158),
.B(n_964),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1248),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1241),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1211),
.B(n_1109),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_SL g1311 ( 
.A1(n_1162),
.A2(n_1008),
.B(n_960),
.Y(n_1311)
);

NOR2x1_ASAP7_75t_L g1312 ( 
.A(n_1248),
.B(n_970),
.Y(n_1312)
);

OAI211xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1186),
.A2(n_1076),
.B(n_982),
.C(n_986),
.Y(n_1313)
);

NOR2xp67_ASAP7_75t_L g1314 ( 
.A(n_1142),
.B(n_959),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1241),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1211),
.A2(n_1103),
.B1(n_1015),
.B2(n_1130),
.Y(n_1316)
);

BUFx10_ASAP7_75t_L g1317 ( 
.A(n_1189),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1221),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1292),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1291),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1292),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1146),
.A2(n_1124),
.B(n_1117),
.C(n_1116),
.Y(n_1322)
);

AO21x2_ASAP7_75t_L g1323 ( 
.A1(n_1208),
.A2(n_1009),
.B(n_966),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1208),
.A2(n_1107),
.B(n_1019),
.Y(n_1324)
);

BUFx12f_ASAP7_75t_L g1325 ( 
.A(n_1190),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1196),
.A2(n_1019),
.B(n_1008),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1233),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1292),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1248),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1274),
.A2(n_1133),
.B(n_1127),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1292),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1289),
.A2(n_1070),
.B(n_1058),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1263),
.Y(n_1333)
);

AOI21xp33_ASAP7_75t_L g1334 ( 
.A1(n_1218),
.A2(n_1032),
.B(n_1054),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1258),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1152),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1144),
.A2(n_1070),
.B(n_1058),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1140),
.A2(n_1125),
.B1(n_964),
.B2(n_959),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1157),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1165),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1263),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1176),
.A2(n_1036),
.B1(n_1085),
.B2(n_1095),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1177),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1276),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1218),
.A2(n_959),
.B1(n_1032),
.B2(n_1073),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1196),
.A2(n_1038),
.B(n_1024),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1199),
.A2(n_1038),
.B(n_1024),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1163),
.A2(n_957),
.B(n_1032),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1199),
.A2(n_1082),
.B(n_1052),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1180),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1276),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1256),
.B(n_1054),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1206),
.A2(n_1082),
.B(n_1052),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1235),
.A2(n_1246),
.B1(n_1261),
.B2(n_1285),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1158),
.B(n_1036),
.Y(n_1355)
);

AO22x2_ASAP7_75t_L g1356 ( 
.A1(n_1264),
.A2(n_1300),
.B1(n_1167),
.B2(n_1171),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1283),
.A2(n_1081),
.B1(n_1009),
.B2(n_1015),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1203),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1206),
.A2(n_1298),
.B(n_1277),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1228),
.Y(n_1360)
);

AOI211xp5_ASAP7_75t_L g1361 ( 
.A1(n_1191),
.A2(n_1037),
.B(n_1110),
.C(n_1117),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1277),
.Y(n_1362)
);

INVx6_ASAP7_75t_L g1363 ( 
.A(n_1221),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1221),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1298),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1299),
.A2(n_1092),
.B(n_1088),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1247),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1299),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1223),
.A2(n_1092),
.B(n_1088),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1306),
.B(n_1131),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1223),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1147),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1164),
.B(n_1131),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1239),
.A2(n_1134),
.B(n_1137),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1187),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1239),
.A2(n_1134),
.B(n_1010),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1285),
.A2(n_1054),
.B1(n_1073),
.B2(n_1094),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1221),
.Y(n_1378)
);

CKINVDCx14_ASAP7_75t_R g1379 ( 
.A(n_1190),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_SL g1380 ( 
.A(n_1200),
.B(n_1061),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1250),
.A2(n_1254),
.B(n_1251),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1250),
.A2(n_1010),
.B(n_1003),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1251),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1193),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1145),
.A2(n_955),
.B(n_1119),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1161),
.B(n_1095),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1254),
.A2(n_1022),
.B(n_1003),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1271),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1257),
.A2(n_1022),
.B(n_1003),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1257),
.A2(n_1068),
.B(n_1022),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1213),
.A2(n_1068),
.B(n_1035),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1213),
.A2(n_1068),
.B(n_1027),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1141),
.A2(n_1020),
.B(n_1049),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1170),
.B(n_998),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1271),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1145),
.A2(n_1123),
.B(n_1112),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1159),
.A2(n_1050),
.B(n_969),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1159),
.A2(n_1160),
.B(n_1181),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1172),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1148),
.A2(n_1101),
.B(n_1113),
.C(n_995),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1270),
.A2(n_1073),
.B1(n_1081),
.B2(n_1056),
.Y(n_1401)
);

AO21x1_ASAP7_75t_L g1402 ( 
.A1(n_1141),
.A2(n_1230),
.B(n_1197),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1303),
.B(n_998),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1286),
.A2(n_1123),
.B(n_1112),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1203),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1160),
.A2(n_1181),
.B(n_1139),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1271),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1172),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1175),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1273),
.B(n_998),
.Y(n_1410)
);

OR2x6_ASAP7_75t_L g1411 ( 
.A(n_1280),
.B(n_1020),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1175),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1262),
.A2(n_1056),
.B1(n_1018),
.B2(n_980),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1139),
.A2(n_563),
.B(n_561),
.Y(n_1414)
);

INVx6_ASAP7_75t_L g1415 ( 
.A(n_1256),
.Y(n_1415)
);

AOI222xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1282),
.A2(n_516),
.B1(n_515),
.B2(n_513),
.C1(n_509),
.C2(n_506),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_1179),
.B(n_1020),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1143),
.A2(n_1123),
.B(n_1112),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1279),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1265),
.A2(n_1018),
.B1(n_1056),
.B2(n_980),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1256),
.B(n_980),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1271),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_SL g1423 ( 
.A1(n_1194),
.A2(n_578),
.B(n_575),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1291),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1209),
.Y(n_1425)
);

OR2x6_ASAP7_75t_L g1426 ( 
.A(n_1150),
.B(n_968),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1245),
.Y(n_1427)
);

CKINVDCx12_ASAP7_75t_R g1428 ( 
.A(n_1302),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1155),
.A2(n_578),
.B(n_563),
.Y(n_1429)
);

AO31x2_ASAP7_75t_L g1430 ( 
.A1(n_1207),
.A2(n_578),
.A3(n_575),
.B(n_574),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1148),
.A2(n_1136),
.B(n_1135),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1209),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1267),
.A2(n_1136),
.B(n_1135),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1174),
.B(n_981),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1260),
.B(n_992),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1260),
.A2(n_1273),
.B1(n_1224),
.B2(n_1288),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1297),
.A2(n_1033),
.B(n_991),
.C(n_992),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1155),
.A2(n_1168),
.B(n_1154),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1143),
.A2(n_1136),
.B(n_1135),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1279),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1272),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1174),
.B(n_981),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1175),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1293),
.B(n_1153),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1149),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1168),
.A2(n_574),
.B(n_497),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1249),
.Y(n_1447)
);

INVx4_ASAP7_75t_SL g1448 ( 
.A(n_1202),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1269),
.A2(n_1018),
.B1(n_1056),
.B2(n_992),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1154),
.A2(n_515),
.B(n_504),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1275),
.A2(n_1098),
.B(n_504),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_SL g1452 ( 
.A(n_1295),
.B(n_1049),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1284),
.B(n_1000),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1205),
.A2(n_1098),
.B(n_1018),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1255),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1151),
.A2(n_516),
.B(n_506),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1151),
.A2(n_509),
.B(n_513),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1220),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1149),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1156),
.A2(n_1049),
.B(n_1091),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1175),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1173),
.A2(n_1029),
.B(n_1028),
.C(n_1000),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1259),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1201),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1184),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1268),
.A2(n_1130),
.B1(n_1132),
.B2(n_1098),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1293),
.B(n_1004),
.Y(n_1467)
);

OAI21xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1214),
.A2(n_1132),
.B(n_1091),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1156),
.A2(n_394),
.B(n_359),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1200),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1217),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1169),
.A2(n_1091),
.B(n_1080),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1222),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1189),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1238),
.B(n_1004),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1225),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1153),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_SL g1478 ( 
.A1(n_1219),
.A2(n_968),
.B(n_1006),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1268),
.A2(n_1132),
.B1(n_1029),
.B2(n_1028),
.Y(n_1479)
);

AOI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1149),
.A2(n_1132),
.B(n_1091),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1166),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1295),
.A2(n_1080),
.B(n_1006),
.Y(n_1482)
);

AO21x1_ASAP7_75t_L g1483 ( 
.A1(n_1183),
.A2(n_266),
.B(n_307),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1336),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1310),
.A2(n_1150),
.B1(n_971),
.B2(n_974),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1307),
.B(n_1120),
.Y(n_1486)
);

INVx6_ASAP7_75t_L g1487 ( 
.A(n_1317),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1327),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1354),
.A2(n_1294),
.B1(n_1150),
.B2(n_974),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1404),
.A2(n_1393),
.B(n_1411),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1336),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1313),
.A2(n_1294),
.B1(n_971),
.B2(n_1296),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1357),
.A2(n_1229),
.B1(n_1231),
.B2(n_1080),
.Y(n_1493)
);

INVx5_ASAP7_75t_L g1494 ( 
.A(n_1318),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1339),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1384),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1406),
.A2(n_1173),
.B(n_1169),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1308),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1309),
.B(n_1202),
.Y(n_1499)
);

AO21x2_ASAP7_75t_L g1500 ( 
.A1(n_1311),
.A2(n_1185),
.B(n_1183),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1465),
.A2(n_1253),
.B1(n_1293),
.B2(n_1080),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1384),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1309),
.B(n_1202),
.Y(n_1503)
);

AND2x2_ASAP7_75t_SL g1504 ( 
.A(n_1385),
.B(n_968),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1339),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1315),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1441),
.B(n_1207),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1352),
.B(n_1304),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1340),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1340),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1343),
.Y(n_1511)
);

BUFx12f_ASAP7_75t_L g1512 ( 
.A(n_1325),
.Y(n_1512)
);

A2O1A1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1400),
.A2(n_1215),
.B(n_1227),
.C(n_1242),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1372),
.B(n_1215),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1463),
.A2(n_1304),
.B1(n_968),
.B2(n_1006),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1315),
.B(n_1202),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1357),
.A2(n_1006),
.B1(n_1226),
.B2(n_1153),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1308),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1343),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1363),
.Y(n_1520)
);

OAI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1436),
.A2(n_404),
.B1(n_410),
.B2(n_409),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1361),
.B(n_1226),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1446),
.A2(n_1192),
.B(n_1178),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_1327),
.Y(n_1524)
);

OAI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1436),
.A2(n_380),
.B1(n_379),
.B2(n_396),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1358),
.Y(n_1526)
);

OR2x6_ASAP7_75t_L g1527 ( 
.A(n_1411),
.B(n_1278),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1428),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1350),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1372),
.B(n_1227),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1370),
.B(n_1386),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1345),
.A2(n_1226),
.B1(n_1243),
.B2(n_1185),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1481),
.A2(n_1304),
.B1(n_1220),
.B2(n_266),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1440),
.Y(n_1534)
);

AO21x2_ASAP7_75t_L g1535 ( 
.A1(n_1311),
.A2(n_1188),
.B(n_1287),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1350),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1370),
.B(n_1244),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1386),
.B(n_1244),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1356),
.A2(n_373),
.B1(n_362),
.B2(n_412),
.C(n_1266),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1358),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_SL g1541 ( 
.A1(n_1361),
.A2(n_1290),
.B1(n_1234),
.B2(n_1240),
.C(n_1237),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1375),
.B(n_1244),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1446),
.A2(n_1182),
.B(n_1236),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1320),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1308),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1405),
.A2(n_1220),
.B1(n_1237),
.B2(n_22),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1375),
.B(n_1244),
.Y(n_1547)
);

AO21x2_ASAP7_75t_L g1548 ( 
.A1(n_1462),
.A2(n_1305),
.B(n_1210),
.Y(n_1548)
);

NOR3xp33_ASAP7_75t_L g1549 ( 
.A(n_1334),
.B(n_1322),
.C(n_1437),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_R g1550 ( 
.A1(n_1342),
.A2(n_1237),
.B(n_307),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1320),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1360),
.Y(n_1552)
);

AOI211xp5_ASAP7_75t_L g1553 ( 
.A1(n_1314),
.A2(n_1237),
.B(n_266),
.C(n_22),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1424),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1338),
.A2(n_266),
.B1(n_1252),
.B2(n_1281),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1435),
.A2(n_266),
.B1(n_1198),
.B2(n_1216),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1373),
.B(n_1232),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1435),
.A2(n_266),
.B1(n_1195),
.B2(n_1212),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1380),
.A2(n_1204),
.B1(n_1232),
.B2(n_610),
.Y(n_1559)
);

INVx8_ASAP7_75t_L g1560 ( 
.A(n_1318),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1405),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1360),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1424),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1403),
.B(n_20),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1475),
.A2(n_610),
.B1(n_539),
.B2(n_1232),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1318),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1373),
.B(n_1232),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1470),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1475),
.A2(n_1377),
.B1(n_1314),
.B2(n_1316),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1355),
.B(n_21),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1318),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1352),
.A2(n_610),
.B1(n_539),
.B2(n_692),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1367),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_SL g1574 ( 
.A(n_1404),
.B(n_1411),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1466),
.B(n_610),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1379),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1352),
.A2(n_610),
.B1(n_539),
.B2(n_1301),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1428),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1352),
.B(n_105),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1318),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1367),
.Y(n_1581)
);

NAND2x1p5_ASAP7_75t_L g1582 ( 
.A(n_1378),
.B(n_766),
.Y(n_1582)
);

NOR3xp33_ASAP7_75t_SL g1583 ( 
.A(n_1468),
.B(n_21),
.C(n_23),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1471),
.B(n_23),
.Y(n_1584)
);

CKINVDCx6p67_ASAP7_75t_R g1585 ( 
.A(n_1325),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1434),
.B(n_24),
.Y(n_1586)
);

OAI21xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1427),
.A2(n_206),
.B(n_203),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1466),
.A2(n_610),
.B1(n_25),
.B2(n_26),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1363),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1410),
.A2(n_610),
.B1(n_539),
.B2(n_766),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1471),
.B(n_107),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1473),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_SL g1593 ( 
.A1(n_1356),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1479),
.A2(n_766),
.B1(n_539),
.B2(n_33),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1473),
.B(n_200),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1476),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_SL g1597 ( 
.A1(n_1356),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1476),
.B(n_30),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1470),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1317),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1401),
.A2(n_766),
.B1(n_34),
.B2(n_36),
.Y(n_1601)
);

OAI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1474),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1356),
.A2(n_722),
.B1(n_676),
.B2(n_40),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1421),
.A2(n_722),
.B1(n_676),
.B2(n_48),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1421),
.B(n_37),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1425),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1413),
.A2(n_38),
.B1(n_51),
.B2(n_53),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1434),
.B(n_51),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1432),
.Y(n_1609)
);

OAI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1426),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1416),
.A2(n_676),
.B1(n_722),
.B2(n_62),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1464),
.B(n_54),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1388),
.Y(n_1613)
);

OAI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1420),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.C(n_69),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1415),
.A2(n_61),
.B1(n_67),
.B2(n_71),
.Y(n_1615)
);

AOI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1431),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.C(n_75),
.Y(n_1616)
);

AND2x2_ASAP7_75t_SL g1617 ( 
.A(n_1385),
.B(n_73),
.Y(n_1617)
);

OAI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1426),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1317),
.Y(n_1619)
);

OR2x6_ASAP7_75t_L g1620 ( 
.A(n_1411),
.B(n_116),
.Y(n_1620)
);

INVx3_ASAP7_75t_SL g1621 ( 
.A(n_1317),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1444),
.B(n_121),
.Y(n_1622)
);

AO21x2_ASAP7_75t_L g1623 ( 
.A1(n_1406),
.A2(n_197),
.B(n_192),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1450),
.A2(n_188),
.B(n_178),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1415),
.A2(n_77),
.B1(n_78),
.B2(n_82),
.Y(n_1625)
);

AND2x2_ASAP7_75t_SL g1626 ( 
.A(n_1385),
.B(n_83),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1464),
.B(n_85),
.Y(n_1627)
);

INVx4_ASAP7_75t_L g1628 ( 
.A(n_1363),
.Y(n_1628)
);

AND2x2_ASAP7_75t_SL g1629 ( 
.A(n_1385),
.B(n_86),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1432),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1415),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1329),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1388),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1404),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1363),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1449),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.C(n_95),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1378),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1395),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1444),
.B(n_156),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1395),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1467),
.B(n_155),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1450),
.A2(n_157),
.B(n_174),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1415),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1419),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_SL g1645 ( 
.A1(n_1454),
.A2(n_132),
.B(n_140),
.C(n_153),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1444),
.B(n_163),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1394),
.B(n_175),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1442),
.B(n_164),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1426),
.A2(n_171),
.B1(n_1419),
.B2(n_1453),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1444),
.B(n_1427),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1329),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1407),
.Y(n_1652)
);

BUFx2_ASAP7_75t_L g1653 ( 
.A(n_1443),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1407),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_SL g1655 ( 
.A(n_1332),
.B(n_1402),
.C(n_1483),
.Y(n_1655)
);

INVx6_ASAP7_75t_L g1656 ( 
.A(n_1378),
.Y(n_1656)
);

AOI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1480),
.A2(n_1330),
.B(n_1422),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1467),
.B(n_1426),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1335),
.B(n_1447),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1426),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1337),
.A2(n_1348),
.B1(n_1402),
.B2(n_1335),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1422),
.Y(n_1662)
);

OAI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1458),
.A2(n_1442),
.B1(n_1447),
.B2(n_1455),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1458),
.A2(n_1423),
.B1(n_1433),
.B2(n_1467),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1319),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1521),
.A2(n_1423),
.B1(n_1458),
.B2(n_1467),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1484),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1613),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1491),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1633),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1525),
.A2(n_1483),
.B1(n_1478),
.B2(n_1455),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1602),
.A2(n_1616),
.B1(n_1636),
.B2(n_1614),
.C(n_1588),
.Y(n_1672)
);

NAND2x1p5_ASAP7_75t_L g1673 ( 
.A(n_1617),
.B(n_1439),
.Y(n_1673)
);

NAND3xp33_ASAP7_75t_L g1674 ( 
.A(n_1549),
.B(n_1469),
.C(n_1468),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1569),
.A2(n_1478),
.B1(n_1323),
.B2(n_1448),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1489),
.A2(n_1411),
.B1(n_1417),
.B2(n_1329),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1486),
.A2(n_1417),
.B1(n_1364),
.B2(n_1312),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1538),
.B(n_1445),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1495),
.Y(n_1679)
);

AOI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1539),
.A2(n_1319),
.B1(n_1321),
.B2(n_1331),
.C(n_1328),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1593),
.A2(n_1323),
.B1(n_1448),
.B2(n_1451),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1597),
.A2(n_1323),
.B1(n_1448),
.B2(n_1451),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1487),
.Y(n_1683)
);

AO21x2_ASAP7_75t_L g1684 ( 
.A1(n_1655),
.A2(n_1438),
.B(n_1398),
.Y(n_1684)
);

CKINVDCx14_ASAP7_75t_R g1685 ( 
.A(n_1576),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1607),
.A2(n_1448),
.B1(n_1451),
.B2(n_1477),
.Y(n_1686)
);

AOI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1610),
.A2(n_1461),
.B(n_1409),
.C(n_1457),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1634),
.A2(n_1477),
.B1(n_1418),
.B2(n_1417),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1486),
.A2(n_1418),
.B1(n_1417),
.B2(n_1469),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1618),
.A2(n_1321),
.B1(n_1328),
.B2(n_1331),
.C(n_1459),
.Y(n_1690)
);

AOI222xp33_ASAP7_75t_L g1691 ( 
.A1(n_1643),
.A2(n_1452),
.B1(n_1459),
.B2(n_1445),
.C1(n_1397),
.C2(n_1461),
.Y(n_1691)
);

OAI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1615),
.A2(n_1469),
.B1(n_1417),
.B2(n_1312),
.C(n_1364),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1631),
.A2(n_1418),
.B1(n_1469),
.B2(n_1412),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1531),
.B(n_1409),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1492),
.A2(n_1412),
.B1(n_1409),
.B2(n_1439),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1528),
.A2(n_1578),
.B1(n_1626),
.B2(n_1617),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1601),
.A2(n_1365),
.B1(n_1362),
.B2(n_1368),
.C(n_1344),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1553),
.A2(n_1365),
.B1(n_1362),
.B2(n_1368),
.C(n_1344),
.Y(n_1698)
);

AOI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1594),
.A2(n_1351),
.B1(n_1341),
.B2(n_1333),
.C(n_1399),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1626),
.B(n_1396),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1546),
.A2(n_1378),
.B1(n_1452),
.B2(n_1364),
.Y(n_1701)
);

BUFx12f_ASAP7_75t_L g1702 ( 
.A(n_1512),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1490),
.A2(n_1396),
.B(n_1439),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1659),
.B(n_1409),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1524),
.B(n_1409),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_SL g1706 ( 
.A1(n_1600),
.A2(n_1412),
.B1(n_1378),
.B2(n_1396),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1501),
.A2(n_1412),
.B1(n_1480),
.B2(n_1351),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1488),
.B(n_1430),
.Y(n_1708)
);

OAI211xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1625),
.A2(n_1399),
.B(n_1408),
.C(n_1333),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1550),
.A2(n_1600),
.B1(n_1485),
.B2(n_1660),
.Y(n_1710)
);

OAI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1583),
.A2(n_1408),
.B1(n_1396),
.B2(n_1439),
.C(n_1341),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1660),
.A2(n_1507),
.B1(n_1599),
.B2(n_1611),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1629),
.A2(n_1482),
.B1(n_1397),
.B2(n_1392),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1599),
.A2(n_1330),
.B1(n_1383),
.B2(n_1371),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1629),
.A2(n_1482),
.B1(n_1392),
.B2(n_1391),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1575),
.A2(n_1482),
.B1(n_1391),
.B2(n_1383),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1575),
.A2(n_1371),
.B1(n_1460),
.B2(n_1456),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1513),
.A2(n_1645),
.B(n_1603),
.C(n_1587),
.Y(n_1718)
);

OAI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1513),
.A2(n_1430),
.B1(n_1398),
.B2(n_1457),
.C(n_1456),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1620),
.A2(n_1460),
.B1(n_1472),
.B2(n_1376),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1496),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1568),
.A2(n_1430),
.B1(n_1472),
.B2(n_1382),
.Y(n_1722)
);

NOR2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1585),
.B(n_1430),
.Y(n_1723)
);

OAI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1533),
.A2(n_1430),
.B1(n_1429),
.B2(n_1414),
.C(n_1347),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1499),
.B(n_1326),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1638),
.Y(n_1726)
);

OAI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1564),
.A2(n_1429),
.B1(n_1347),
.B2(n_1349),
.C(n_1353),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1568),
.A2(n_1534),
.B1(n_1619),
.B2(n_1515),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1505),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1502),
.A2(n_1382),
.B1(n_1376),
.B2(n_1366),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1661),
.A2(n_1349),
.B1(n_1353),
.B2(n_1346),
.C(n_1326),
.Y(n_1731)
);

AOI21xp33_ASAP7_75t_L g1732 ( 
.A1(n_1647),
.A2(n_1346),
.B(n_1374),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1620),
.A2(n_1579),
.B1(n_1522),
.B2(n_1648),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1620),
.A2(n_1366),
.B1(n_1374),
.B2(n_1369),
.Y(n_1734)
);

AOI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1570),
.A2(n_1649),
.B1(n_1559),
.B2(n_1627),
.C(n_1612),
.Y(n_1735)
);

AOI222xp33_ASAP7_75t_L g1736 ( 
.A1(n_1584),
.A2(n_1369),
.B1(n_1324),
.B2(n_1387),
.C1(n_1389),
.C2(n_1390),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1598),
.A2(n_1324),
.B1(n_1359),
.B2(n_1387),
.C(n_1389),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1487),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1650),
.B(n_1390),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1620),
.A2(n_1359),
.B1(n_1381),
.B2(n_1579),
.Y(n_1740)
);

OA21x2_ASAP7_75t_L g1741 ( 
.A1(n_1523),
.A2(n_1381),
.B(n_1541),
.Y(n_1741)
);

AOI21xp33_ASAP7_75t_L g1742 ( 
.A1(n_1514),
.A2(n_1530),
.B(n_1645),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1579),
.A2(n_1522),
.B1(n_1648),
.B2(n_1658),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1663),
.A2(n_1605),
.B1(n_1537),
.B2(n_1604),
.C(n_1493),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1658),
.A2(n_1641),
.B1(n_1508),
.B2(n_1639),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1586),
.A2(n_1608),
.B1(n_1542),
.B2(n_1547),
.C(n_1532),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1621),
.A2(n_1664),
.B1(n_1554),
.B2(n_1563),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1499),
.B(n_1503),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1650),
.B(n_1592),
.Y(n_1749)
);

OAI211xp5_ASAP7_75t_L g1750 ( 
.A1(n_1596),
.A2(n_1595),
.B(n_1591),
.C(n_1552),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1591),
.B(n_1595),
.C(n_1555),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1658),
.A2(n_1641),
.B1(n_1508),
.B2(n_1622),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1498),
.Y(n_1753)
);

AOI21xp33_ASAP7_75t_L g1754 ( 
.A1(n_1517),
.A2(n_1556),
.B(n_1558),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1653),
.B(n_1508),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1585),
.A2(n_1576),
.B1(n_1526),
.B2(n_1561),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1498),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1526),
.B(n_1540),
.Y(n_1758)
);

OAI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1621),
.A2(n_1540),
.B1(n_1561),
.B2(n_1544),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1509),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1641),
.A2(n_1639),
.B1(n_1622),
.B2(n_1646),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1665),
.B(n_1654),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1646),
.A2(n_1512),
.B1(n_1487),
.B2(n_1644),
.Y(n_1763)
);

AOI21xp33_ASAP7_75t_L g1764 ( 
.A1(n_1535),
.A2(n_1527),
.B(n_1590),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1565),
.A2(n_1581),
.B1(n_1573),
.B2(n_1562),
.C(n_1536),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1544),
.Y(n_1766)
);

AOI222xp33_ASAP7_75t_L g1767 ( 
.A1(n_1510),
.A2(n_1519),
.B1(n_1529),
.B2(n_1511),
.C1(n_1516),
.C2(n_1503),
.Y(n_1767)
);

OR2x6_ASAP7_75t_L g1768 ( 
.A(n_1527),
.B(n_1516),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1662),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1551),
.A2(n_1628),
.B1(n_1520),
.B2(n_1589),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1551),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1520),
.A2(n_1628),
.B1(n_1589),
.B2(n_1635),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1520),
.A2(n_1628),
.B1(n_1635),
.B2(n_1623),
.Y(n_1773)
);

OAI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1527),
.A2(n_1572),
.B1(n_1577),
.B2(n_1656),
.C(n_1651),
.Y(n_1774)
);

CKINVDCx20_ASAP7_75t_R g1775 ( 
.A(n_1656),
.Y(n_1775)
);

CKINVDCx11_ASAP7_75t_R g1776 ( 
.A(n_1560),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1527),
.A2(n_1656),
.B1(n_1623),
.B2(n_1637),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1640),
.Y(n_1778)
);

AOI222xp33_ASAP7_75t_L g1779 ( 
.A1(n_1557),
.A2(n_1567),
.B1(n_1504),
.B2(n_1506),
.C1(n_1574),
.C2(n_1652),
.Y(n_1779)
);

OAI211xp5_ASAP7_75t_L g1780 ( 
.A1(n_1506),
.A2(n_1657),
.B(n_1560),
.C(n_1498),
.Y(n_1780)
);

OAI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1494),
.A2(n_1571),
.B1(n_1637),
.B2(n_1580),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1518),
.A2(n_1651),
.B1(n_1632),
.B2(n_1545),
.C(n_1494),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1606),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1606),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1518),
.B(n_1651),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1504),
.A2(n_1518),
.B1(n_1632),
.B2(n_1545),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1545),
.A2(n_1632),
.B1(n_1500),
.B2(n_1535),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1566),
.B(n_1571),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1609),
.A2(n_1630),
.B1(n_1560),
.B2(n_1580),
.C(n_1637),
.Y(n_1789)
);

OAI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1494),
.A2(n_1566),
.B1(n_1637),
.B2(n_1580),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1497),
.Y(n_1791)
);

INVx4_ASAP7_75t_L g1792 ( 
.A(n_1494),
.Y(n_1792)
);

NAND4xp25_ASAP7_75t_L g1793 ( 
.A(n_1560),
.B(n_1500),
.C(n_1642),
.D(n_1624),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1494),
.A2(n_1566),
.B1(n_1580),
.B2(n_1571),
.Y(n_1794)
);

AOI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1566),
.A2(n_1571),
.B1(n_1548),
.B2(n_1500),
.C(n_1582),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1548),
.A2(n_1624),
.B1(n_1642),
.B2(n_1497),
.Y(n_1796)
);

OAI21x1_ASAP7_75t_L g1797 ( 
.A1(n_1543),
.A2(n_1523),
.B(n_1497),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1548),
.Y(n_1798)
);

OAI222xp33_ASAP7_75t_L g1799 ( 
.A1(n_1582),
.A2(n_1614),
.B1(n_1636),
.B2(n_1593),
.C1(n_1597),
.C2(n_1625),
.Y(n_1799)
);

BUFx4f_ASAP7_75t_SL g1800 ( 
.A(n_1512),
.Y(n_1800)
);

OA21x2_ASAP7_75t_L g1801 ( 
.A1(n_1523),
.A2(n_1406),
.B(n_1398),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1617),
.B(n_1626),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1521),
.A2(n_989),
.B1(n_1525),
.B2(n_1616),
.Y(n_1803)
);

NAND4xp25_ASAP7_75t_L g1804 ( 
.A(n_1616),
.B(n_867),
.C(n_1186),
.D(n_702),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1617),
.B(n_1626),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1521),
.A2(n_1186),
.B1(n_867),
.B2(n_1525),
.C(n_1072),
.Y(n_1806)
);

OAI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1614),
.A2(n_1047),
.B1(n_1078),
.B2(n_1636),
.Y(n_1807)
);

OAI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1616),
.A2(n_687),
.B1(n_1354),
.B2(n_1002),
.C(n_921),
.Y(n_1808)
);

OAI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1614),
.A2(n_1047),
.B1(n_1078),
.B2(n_1636),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_SL g1810 ( 
.A1(n_1546),
.A2(n_1002),
.B1(n_603),
.B2(n_1047),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1498),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1613),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1521),
.A2(n_989),
.B1(n_1525),
.B2(n_1616),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1617),
.B(n_1626),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1613),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1484),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1484),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1531),
.B(n_1659),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1613),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1498),
.Y(n_1820)
);

NAND2x1p5_ASAP7_75t_L g1821 ( 
.A(n_1617),
.B(n_1626),
.Y(n_1821)
);

OAI211xp5_ASAP7_75t_L g1822 ( 
.A1(n_1615),
.A2(n_867),
.B(n_1625),
.C(n_1186),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_SL g1823 ( 
.A1(n_1546),
.A2(n_1002),
.B1(n_603),
.B2(n_1047),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1490),
.A2(n_1141),
.B(n_793),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1791),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1668),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1748),
.B(n_1725),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1748),
.B(n_1725),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1678),
.B(n_1798),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1762),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1700),
.B(n_1768),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1668),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1768),
.B(n_1739),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1700),
.B(n_1768),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1791),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1670),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1670),
.Y(n_1837)
);

NOR2x1_ASAP7_75t_L g1838 ( 
.A(n_1780),
.B(n_1674),
.Y(n_1838)
);

AO31x2_ASAP7_75t_L g1839 ( 
.A1(n_1703),
.A2(n_1714),
.A3(n_1718),
.B(n_1722),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1726),
.Y(n_1840)
);

INVxp67_ASAP7_75t_SL g1841 ( 
.A(n_1708),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1726),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1768),
.B(n_1673),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1673),
.B(n_1812),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1683),
.Y(n_1845)
);

BUFx2_ASAP7_75t_L g1846 ( 
.A(n_1673),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1812),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1762),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1678),
.B(n_1818),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1815),
.B(n_1819),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1741),
.B(n_1684),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1819),
.Y(n_1852)
);

INVx4_ASAP7_75t_L g1853 ( 
.A(n_1792),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1741),
.B(n_1684),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1769),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1804),
.A2(n_1806),
.B1(n_1672),
.B2(n_1808),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1741),
.B(n_1779),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1778),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1667),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1669),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1684),
.B(n_1787),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1767),
.B(n_1746),
.Y(n_1862)
);

NAND2x1_ASAP7_75t_L g1863 ( 
.A(n_1792),
.B(n_1777),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1801),
.B(n_1749),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1679),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1729),
.B(n_1760),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1802),
.B(n_1805),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1816),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1810),
.A2(n_1823),
.B1(n_1803),
.B2(n_1813),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1802),
.B(n_1805),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1807),
.A2(n_1809),
.B1(n_1712),
.B2(n_1735),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1814),
.B(n_1821),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1817),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1783),
.B(n_1784),
.Y(n_1874)
);

AND2x4_ASAP7_75t_SL g1875 ( 
.A(n_1792),
.B(n_1721),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1814),
.B(n_1821),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_SL g1877 ( 
.A1(n_1821),
.A2(n_1822),
.B1(n_1750),
.B2(n_1710),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1715),
.B(n_1713),
.Y(n_1878)
);

BUFx3_ASAP7_75t_L g1879 ( 
.A(n_1683),
.Y(n_1879)
);

OAI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1774),
.A2(n_1698),
.B1(n_1751),
.B2(n_1692),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1797),
.Y(n_1881)
);

BUFx2_ASAP7_75t_L g1882 ( 
.A(n_1706),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1801),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1796),
.B(n_1694),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1730),
.B(n_1711),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1680),
.B(n_1704),
.Y(n_1886)
);

HB1xp67_ASAP7_75t_L g1887 ( 
.A(n_1785),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1689),
.B(n_1793),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1753),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1753),
.B(n_1757),
.Y(n_1890)
);

OAI221xp5_ASAP7_75t_SL g1891 ( 
.A1(n_1733),
.A2(n_1696),
.B1(n_1718),
.B2(n_1744),
.C(n_1687),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1716),
.B(n_1720),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1757),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1811),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1701),
.A2(n_1709),
.B1(n_1754),
.B2(n_1685),
.Y(n_1895)
);

INVxp67_ASAP7_75t_SL g1896 ( 
.A(n_1736),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1820),
.B(n_1734),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1755),
.B(n_1764),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1738),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1820),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1786),
.B(n_1820),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1795),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1727),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1705),
.B(n_1747),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1719),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1766),
.A2(n_1756),
.B1(n_1799),
.B2(n_1759),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1782),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1728),
.B(n_1677),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1707),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1731),
.B(n_1737),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1723),
.B(n_1773),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1765),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1858),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1856),
.A2(n_1743),
.B1(n_1685),
.B2(n_1676),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1856),
.A2(n_1763),
.B1(n_1752),
.B2(n_1745),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1906),
.A2(n_1775),
.B1(n_1761),
.B2(n_1702),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1906),
.A2(n_1742),
.B1(n_1681),
.B2(n_1682),
.C(n_1690),
.Y(n_1917)
);

OAI222xp33_ASAP7_75t_L g1918 ( 
.A1(n_1891),
.A2(n_1877),
.B1(n_1862),
.B2(n_1871),
.C1(n_1869),
.C2(n_1880),
.Y(n_1918)
);

OA222x2_ASAP7_75t_L g1919 ( 
.A1(n_1888),
.A2(n_1675),
.B1(n_1740),
.B2(n_1790),
.C1(n_1781),
.C2(n_1824),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1843),
.B(n_1738),
.Y(n_1920)
);

OAI321xp33_ASAP7_75t_L g1921 ( 
.A1(n_1891),
.A2(n_1880),
.A3(n_1871),
.B1(n_1869),
.B2(n_1896),
.C(n_1862),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1841),
.B(n_1693),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1827),
.B(n_1691),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1908),
.A2(n_1702),
.B1(n_1666),
.B2(n_1686),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1830),
.Y(n_1925)
);

INVx3_ASAP7_75t_L g1926 ( 
.A(n_1835),
.Y(n_1926)
);

AO21x2_ASAP7_75t_L g1927 ( 
.A1(n_1883),
.A2(n_1732),
.B(n_1724),
.Y(n_1927)
);

OAI211xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1877),
.A2(n_1770),
.B(n_1772),
.C(n_1671),
.Y(n_1928)
);

AOI221xp5_ASAP7_75t_L g1929 ( 
.A1(n_1896),
.A2(n_1771),
.B1(n_1688),
.B2(n_1695),
.C(n_1766),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1836),
.Y(n_1930)
);

OAI21x1_ASAP7_75t_L g1931 ( 
.A1(n_1883),
.A2(n_1717),
.B(n_1794),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1858),
.Y(n_1932)
);

AOI21xp33_ASAP7_75t_SL g1933 ( 
.A1(n_1908),
.A2(n_1758),
.B(n_1911),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1830),
.Y(n_1934)
);

OAI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1895),
.A2(n_1771),
.B1(n_1789),
.B2(n_1788),
.C(n_1697),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1833),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_SL g1937 ( 
.A1(n_1882),
.A2(n_1775),
.B1(n_1800),
.B2(n_1776),
.Y(n_1937)
);

INVxp67_ASAP7_75t_L g1938 ( 
.A(n_1848),
.Y(n_1938)
);

OAI33xp33_ASAP7_75t_L g1939 ( 
.A1(n_1912),
.A2(n_1699),
.A3(n_1776),
.B1(n_1902),
.B2(n_1886),
.B3(n_1907),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1827),
.B(n_1828),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_R g1941 ( 
.A(n_1882),
.B(n_1912),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1836),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1849),
.B(n_1887),
.Y(n_1943)
);

INVxp67_ASAP7_75t_SL g1944 ( 
.A(n_1900),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1825),
.Y(n_1945)
);

BUFx3_ASAP7_75t_L g1946 ( 
.A(n_1845),
.Y(n_1946)
);

BUFx2_ASAP7_75t_L g1947 ( 
.A(n_1833),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1836),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1837),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1843),
.B(n_1844),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1849),
.B(n_1887),
.Y(n_1951)
);

NOR5xp2_ASAP7_75t_SL g1952 ( 
.A(n_1838),
.B(n_1895),
.C(n_1902),
.D(n_1841),
.E(n_1839),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1848),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1844),
.Y(n_1954)
);

AOI221xp5_ASAP7_75t_L g1955 ( 
.A1(n_1910),
.A2(n_1903),
.B1(n_1907),
.B2(n_1905),
.C(n_1857),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1825),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1864),
.B(n_1829),
.Y(n_1957)
);

OAI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1911),
.A2(n_1888),
.B1(n_1905),
.B2(n_1904),
.Y(n_1958)
);

OAI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1838),
.A2(n_1888),
.B1(n_1885),
.B2(n_1863),
.C(n_1905),
.Y(n_1959)
);

NAND2xp33_ASAP7_75t_SL g1960 ( 
.A(n_1863),
.B(n_1911),
.Y(n_1960)
);

INVx2_ASAP7_75t_SL g1961 ( 
.A(n_1875),
.Y(n_1961)
);

AOI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1878),
.A2(n_1910),
.B1(n_1876),
.B2(n_1872),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1844),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1878),
.A2(n_1910),
.B1(n_1872),
.B2(n_1876),
.Y(n_1964)
);

OAI321xp33_ASAP7_75t_L g1965 ( 
.A1(n_1885),
.A2(n_1903),
.A3(n_1909),
.B1(n_1886),
.B2(n_1892),
.C(n_1878),
.Y(n_1965)
);

AOI221xp5_ASAP7_75t_L g1966 ( 
.A1(n_1903),
.A2(n_1857),
.B1(n_1909),
.B2(n_1885),
.C(n_1892),
.Y(n_1966)
);

OAI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1904),
.A2(n_1898),
.B1(n_1901),
.B2(n_1884),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1859),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1825),
.Y(n_1969)
);

OAI211xp5_ASAP7_75t_L g1970 ( 
.A1(n_1857),
.A2(n_1892),
.B(n_1901),
.C(n_1898),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1845),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1837),
.Y(n_1972)
);

OR2x2_ASAP7_75t_L g1973 ( 
.A(n_1864),
.B(n_1829),
.Y(n_1973)
);

AOI221xp5_ASAP7_75t_L g1974 ( 
.A1(n_1867),
.A2(n_1870),
.B1(n_1861),
.B2(n_1876),
.C(n_1872),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1837),
.Y(n_1975)
);

OA211x2_ASAP7_75t_L g1976 ( 
.A1(n_1874),
.A2(n_1866),
.B(n_1839),
.C(n_1853),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1859),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1826),
.Y(n_1978)
);

OAI221xp5_ASAP7_75t_L g1979 ( 
.A1(n_1898),
.A2(n_1904),
.B1(n_1884),
.B2(n_1846),
.C(n_1861),
.Y(n_1979)
);

NOR3xp33_ASAP7_75t_SL g1980 ( 
.A(n_1866),
.B(n_1874),
.C(n_1893),
.Y(n_1980)
);

OAI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1884),
.A2(n_1846),
.B1(n_1853),
.B2(n_1870),
.Y(n_1981)
);

NAND4xp25_ASAP7_75t_SL g1982 ( 
.A(n_1867),
.B(n_1870),
.C(n_1834),
.D(n_1831),
.Y(n_1982)
);

OAI211xp5_ASAP7_75t_L g1983 ( 
.A1(n_1861),
.A2(n_1846),
.B(n_1867),
.C(n_1897),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1827),
.B(n_1828),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1933),
.B(n_1833),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1930),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1925),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1943),
.B(n_1828),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1945),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1978),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1951),
.B(n_1833),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1967),
.B(n_1833),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1930),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1942),
.Y(n_1994)
);

NAND2xp33_ASAP7_75t_SL g1995 ( 
.A(n_1941),
.B(n_1831),
.Y(n_1995)
);

AND2x4_ASAP7_75t_L g1996 ( 
.A(n_1950),
.B(n_1843),
.Y(n_1996)
);

AND2x4_ASAP7_75t_L g1997 ( 
.A(n_1950),
.B(n_1834),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1945),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1940),
.B(n_1834),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1940),
.B(n_1831),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1966),
.B(n_1855),
.Y(n_2001)
);

INVx1_ASAP7_75t_SL g2002 ( 
.A(n_1971),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1923),
.B(n_1855),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1936),
.B(n_1897),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1923),
.B(n_1855),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1942),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1948),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1950),
.B(n_1879),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1936),
.B(n_1879),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1958),
.B(n_1897),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1948),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1947),
.B(n_1835),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1949),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1957),
.B(n_1864),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1949),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1970),
.B(n_1962),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1972),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1972),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1964),
.B(n_1873),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1956),
.Y(n_2020)
);

INVxp67_ASAP7_75t_L g2021 ( 
.A(n_1934),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1957),
.B(n_1973),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1973),
.B(n_1829),
.Y(n_2023)
);

NOR2x1_ASAP7_75t_L g2024 ( 
.A(n_1959),
.B(n_1845),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1916),
.A2(n_1875),
.B1(n_1868),
.B2(n_1873),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1947),
.B(n_1835),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1938),
.B(n_1868),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1953),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1954),
.B(n_1835),
.Y(n_2029)
);

NAND2xp33_ASAP7_75t_R g2030 ( 
.A(n_1952),
.B(n_1890),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1955),
.B(n_1865),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1980),
.B(n_1865),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1975),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1963),
.B(n_1835),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1984),
.B(n_1839),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1975),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1974),
.B(n_1860),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1920),
.B(n_1983),
.Y(n_2038)
);

NAND2x1_ASAP7_75t_L g2039 ( 
.A(n_1926),
.B(n_1842),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1944),
.B(n_1839),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1961),
.B(n_1920),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1913),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1920),
.B(n_1850),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1932),
.B(n_1860),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1968),
.B(n_1850),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1926),
.B(n_1850),
.Y(n_2046)
);

HB1xp67_ASAP7_75t_L g2047 ( 
.A(n_1977),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1956),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1922),
.B(n_1890),
.Y(n_2049)
);

INVx1_ASAP7_75t_SL g2050 ( 
.A(n_2002),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_2035),
.B(n_2022),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1990),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_1997),
.B(n_1961),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_2024),
.B(n_1960),
.Y(n_2054)
);

INVxp67_ASAP7_75t_SL g2055 ( 
.A(n_2032),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2001),
.B(n_1922),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2038),
.B(n_1946),
.Y(n_2057)
);

OR2x6_ASAP7_75t_L g2058 ( 
.A(n_1985),
.B(n_1931),
.Y(n_2058)
);

NAND2x1p5_ASAP7_75t_L g2059 ( 
.A(n_2039),
.B(n_2040),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_2035),
.B(n_1979),
.Y(n_2060)
);

BUFx2_ASAP7_75t_SL g2061 ( 
.A(n_2038),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_2022),
.B(n_1982),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1997),
.B(n_1946),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_2014),
.B(n_1969),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2003),
.B(n_1981),
.Y(n_2065)
);

AND2x4_ASAP7_75t_SL g2066 ( 
.A(n_2008),
.B(n_1987),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2047),
.Y(n_2067)
);

AND2x2_ASAP7_75t_SL g2068 ( 
.A(n_2016),
.B(n_2010),
.Y(n_2068)
);

NAND2x1p5_ASAP7_75t_L g2069 ( 
.A(n_2039),
.B(n_1931),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2013),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_2014),
.B(n_1969),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2005),
.B(n_1917),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1989),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_2023),
.B(n_1839),
.Y(n_2074)
);

INVxp67_ASAP7_75t_SL g2075 ( 
.A(n_2030),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2015),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_1995),
.Y(n_2077)
);

AND2x4_ASAP7_75t_L g2078 ( 
.A(n_1997),
.B(n_1926),
.Y(n_2078)
);

OAI21xp5_ASAP7_75t_SL g2079 ( 
.A1(n_2025),
.A2(n_1918),
.B(n_1914),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1996),
.B(n_1919),
.Y(n_2080)
);

NAND3xp33_ASAP7_75t_SL g2081 ( 
.A(n_1995),
.B(n_1937),
.C(n_1929),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1996),
.B(n_1839),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1986),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2023),
.B(n_1839),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_2037),
.B(n_1960),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1986),
.Y(n_2086)
);

INVxp67_ASAP7_75t_L g2087 ( 
.A(n_2031),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1991),
.B(n_2019),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_1992),
.B(n_1921),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1996),
.B(n_2004),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2021),
.B(n_1826),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2004),
.B(n_1890),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1993),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1989),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1999),
.B(n_1890),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1993),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2051),
.B(n_2040),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2073),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2073),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2061),
.B(n_1999),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2051),
.B(n_2028),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2055),
.B(n_2049),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2083),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2075),
.B(n_2090),
.Y(n_2104)
);

INVx1_ASAP7_75t_SL g2105 ( 
.A(n_2054),
.Y(n_2105)
);

INVx2_ASAP7_75t_SL g2106 ( 
.A(n_2066),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_L g2107 ( 
.A(n_2089),
.B(n_1939),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2086),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2087),
.B(n_2042),
.Y(n_2109)
);

NAND2xp33_ASAP7_75t_SL g2110 ( 
.A(n_2054),
.B(n_2008),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2090),
.B(n_2000),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2056),
.B(n_2027),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2093),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2077),
.B(n_2000),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2068),
.B(n_1994),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2060),
.B(n_2045),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2080),
.B(n_2008),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2096),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2068),
.B(n_1994),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2094),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2070),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2094),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2076),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2080),
.B(n_2041),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2059),
.Y(n_2125)
);

INVx1_ASAP7_75t_SL g2126 ( 
.A(n_2050),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2059),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2052),
.Y(n_2128)
);

INVxp67_ASAP7_75t_L g2129 ( 
.A(n_2085),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2091),
.Y(n_2130)
);

NAND3xp33_ASAP7_75t_L g2131 ( 
.A(n_2079),
.B(n_1924),
.C(n_1928),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2082),
.B(n_2041),
.Y(n_2132)
);

NAND2x1_ASAP7_75t_L g2133 ( 
.A(n_2053),
.B(n_2009),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2064),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2064),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2071),
.Y(n_2136)
);

NAND2x1_ASAP7_75t_L g2137 ( 
.A(n_2053),
.B(n_2009),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2072),
.B(n_2011),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_L g2139 ( 
.A(n_2088),
.B(n_1965),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2085),
.B(n_2043),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_2060),
.B(n_1988),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_2067),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2082),
.B(n_2078),
.Y(n_2143)
);

AOI21xp33_ASAP7_75t_SL g2144 ( 
.A1(n_2131),
.A2(n_2062),
.B(n_2058),
.Y(n_2144)
);

OAI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_2105),
.A2(n_2062),
.B1(n_2065),
.B2(n_2058),
.Y(n_2145)
);

AOI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2107),
.A2(n_2081),
.B1(n_2058),
.B2(n_2057),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2121),
.Y(n_2147)
);

OAI221xp5_ASAP7_75t_L g2148 ( 
.A1(n_2131),
.A2(n_2058),
.B1(n_2084),
.B2(n_2074),
.C(n_2069),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2139),
.B(n_2074),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2121),
.Y(n_2150)
);

AOI22xp5_ASAP7_75t_L g2151 ( 
.A1(n_2110),
.A2(n_2057),
.B1(n_1976),
.B2(n_2066),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2123),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2104),
.B(n_2063),
.Y(n_2153)
);

AOI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_2105),
.A2(n_2084),
.B(n_2044),
.Y(n_2154)
);

OAI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_2126),
.A2(n_1952),
.B1(n_1935),
.B2(n_2059),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2123),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2128),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2128),
.Y(n_2158)
);

OAI21xp33_ASAP7_75t_SL g2159 ( 
.A1(n_2115),
.A2(n_2063),
.B(n_2095),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2103),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2138),
.B(n_2071),
.Y(n_2161)
);

NAND3xp33_ASAP7_75t_L g2162 ( 
.A(n_2129),
.B(n_2119),
.C(n_2115),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2104),
.B(n_2053),
.Y(n_2163)
);

OAI221xp5_ASAP7_75t_L g2164 ( 
.A1(n_2119),
.A2(n_2069),
.B1(n_1915),
.B2(n_2018),
.C(n_2006),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2103),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2108),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_2141),
.B(n_2092),
.Y(n_2167)
);

O2A1O1Ixp33_ASAP7_75t_L g2168 ( 
.A1(n_2126),
.A2(n_2069),
.B(n_1927),
.C(n_2007),
.Y(n_2168)
);

AOI32xp33_ASAP7_75t_L g2169 ( 
.A1(n_2100),
.A2(n_2114),
.A3(n_2124),
.B1(n_2117),
.B2(n_2106),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2108),
.Y(n_2170)
);

NAND2x1p5_ASAP7_75t_L g2171 ( 
.A(n_2133),
.B(n_2009),
.Y(n_2171)
);

CKINVDCx16_ASAP7_75t_R g2172 ( 
.A(n_2106),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2124),
.B(n_2092),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2113),
.Y(n_2174)
);

AOI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_2100),
.A2(n_2078),
.B1(n_1927),
.B2(n_2041),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2138),
.B(n_2036),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2117),
.B(n_2095),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2113),
.Y(n_2178)
);

OAI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_2133),
.A2(n_2078),
.B1(n_2043),
.B2(n_2012),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2112),
.A2(n_1927),
.B1(n_2026),
.B2(n_2012),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2112),
.B(n_2033),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2142),
.B(n_2033),
.Y(n_2182)
);

NOR2xp67_ASAP7_75t_L g2183 ( 
.A(n_2151),
.B(n_2114),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2160),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2162),
.B(n_2141),
.Y(n_2185)
);

INVxp67_ASAP7_75t_L g2186 ( 
.A(n_2147),
.Y(n_2186)
);

AOI21xp33_ASAP7_75t_SL g2187 ( 
.A1(n_2155),
.A2(n_2109),
.B(n_2101),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2165),
.Y(n_2188)
);

OAI32xp33_ASAP7_75t_L g2189 ( 
.A1(n_2164),
.A2(n_2097),
.A3(n_2125),
.B1(n_2127),
.B2(n_2101),
.Y(n_2189)
);

OAI221xp5_ASAP7_75t_L g2190 ( 
.A1(n_2146),
.A2(n_2137),
.B1(n_2109),
.B2(n_2130),
.C(n_2102),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2166),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2170),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2174),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2178),
.Y(n_2194)
);

NAND3x2_ASAP7_75t_L g2195 ( 
.A(n_2153),
.B(n_2116),
.C(n_2130),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2172),
.A2(n_2140),
.B1(n_2137),
.B2(n_2116),
.Y(n_2196)
);

INVxp67_ASAP7_75t_L g2197 ( 
.A(n_2150),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2152),
.Y(n_2198)
);

OAI21xp33_ASAP7_75t_L g2199 ( 
.A1(n_2144),
.A2(n_2169),
.B(n_2149),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2163),
.B(n_2111),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2156),
.Y(n_2201)
);

OAI211xp5_ASAP7_75t_L g2202 ( 
.A1(n_2168),
.A2(n_2125),
.B(n_2127),
.C(n_2135),
.Y(n_2202)
);

INVx1_ASAP7_75t_SL g2203 ( 
.A(n_2171),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2157),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2171),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2149),
.B(n_2111),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_2177),
.B(n_2143),
.Y(n_2207)
);

OAI221xp5_ASAP7_75t_L g2208 ( 
.A1(n_2145),
.A2(n_2136),
.B1(n_2135),
.B2(n_2134),
.C(n_2127),
.Y(n_2208)
);

XOR2x2_ASAP7_75t_L g2209 ( 
.A(n_2148),
.B(n_2132),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2173),
.B(n_2143),
.Y(n_2210)
);

OAI322xp33_ASAP7_75t_L g2211 ( 
.A1(n_2180),
.A2(n_2097),
.A3(n_2136),
.B1(n_2134),
.B2(n_2118),
.C1(n_2125),
.C2(n_2099),
.Y(n_2211)
);

AOI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_2199),
.A2(n_2154),
.B(n_2182),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2210),
.B(n_2132),
.Y(n_2213)
);

AOI21xp33_ASAP7_75t_L g2214 ( 
.A1(n_2189),
.A2(n_2158),
.B(n_2159),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2184),
.Y(n_2215)
);

AOI21xp33_ASAP7_75t_L g2216 ( 
.A1(n_2185),
.A2(n_2175),
.B(n_2161),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2210),
.B(n_2207),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2187),
.B(n_2161),
.Y(n_2218)
);

INVxp67_ASAP7_75t_L g2219 ( 
.A(n_2208),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2206),
.B(n_2167),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2207),
.B(n_2181),
.Y(n_2221)
);

INVx1_ASAP7_75t_SL g2222 ( 
.A(n_2203),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2188),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2191),
.Y(n_2224)
);

NOR4xp25_ASAP7_75t_SL g2225 ( 
.A(n_2190),
.B(n_2118),
.C(n_2179),
.D(n_2182),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_L g2226 ( 
.A(n_2200),
.B(n_2181),
.Y(n_2226)
);

OAI21xp5_ASAP7_75t_SL g2227 ( 
.A1(n_2196),
.A2(n_2202),
.B(n_2205),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2192),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2193),
.Y(n_2229)
);

INVx1_ASAP7_75t_SL g2230 ( 
.A(n_2205),
.Y(n_2230)
);

INVxp33_ASAP7_75t_L g2231 ( 
.A(n_2209),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2207),
.B(n_2176),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2194),
.Y(n_2233)
);

INVx2_ASAP7_75t_SL g2234 ( 
.A(n_2198),
.Y(n_2234)
);

INVxp67_ASAP7_75t_SL g2235 ( 
.A(n_2217),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_2222),
.B(n_2209),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_2217),
.B(n_2186),
.Y(n_2237)
);

O2A1O1Ixp33_ASAP7_75t_L g2238 ( 
.A1(n_2231),
.A2(n_2211),
.B(n_2197),
.C(n_2186),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2213),
.B(n_2183),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2213),
.Y(n_2240)
);

AO22x2_ASAP7_75t_L g2241 ( 
.A1(n_2234),
.A2(n_2197),
.B1(n_2201),
.B2(n_2204),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2230),
.B(n_2176),
.Y(n_2242)
);

NAND3xp33_ASAP7_75t_L g2243 ( 
.A(n_2225),
.B(n_2195),
.C(n_2122),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2234),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_L g2245 ( 
.A(n_2232),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2219),
.B(n_2122),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2232),
.Y(n_2247)
);

INVxp67_ASAP7_75t_L g2248 ( 
.A(n_2218),
.Y(n_2248)
);

AND4x1_ASAP7_75t_L g2249 ( 
.A(n_2212),
.B(n_2026),
.C(n_2029),
.D(n_2034),
.Y(n_2249)
);

NAND3xp33_ASAP7_75t_L g2250 ( 
.A(n_2238),
.B(n_2227),
.C(n_2214),
.Y(n_2250)
);

AOI221xp5_ASAP7_75t_L g2251 ( 
.A1(n_2236),
.A2(n_2216),
.B1(n_2226),
.B2(n_2224),
.C(n_2228),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2241),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2235),
.B(n_2221),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_R g2254 ( 
.A(n_2244),
.B(n_2247),
.Y(n_2254)
);

AOI221x1_ASAP7_75t_L g2255 ( 
.A1(n_2241),
.A2(n_2233),
.B1(n_2229),
.B2(n_2228),
.C(n_2223),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2241),
.Y(n_2256)
);

NOR3xp33_ASAP7_75t_SL g2257 ( 
.A(n_2246),
.B(n_2220),
.C(n_2229),
.Y(n_2257)
);

NOR2x1_ASAP7_75t_L g2258 ( 
.A(n_2244),
.B(n_2233),
.Y(n_2258)
);

AOI221x1_ASAP7_75t_L g2259 ( 
.A1(n_2241),
.A2(n_2223),
.B1(n_2215),
.B2(n_2122),
.C(n_2120),
.Y(n_2259)
);

XNOR2xp5_ASAP7_75t_L g2260 ( 
.A(n_2239),
.B(n_2249),
.Y(n_2260)
);

AOI22xp33_ASAP7_75t_L g2261 ( 
.A1(n_2248),
.A2(n_2215),
.B1(n_2120),
.B2(n_2099),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2240),
.Y(n_2262)
);

O2A1O1Ixp33_ASAP7_75t_L g2263 ( 
.A1(n_2243),
.A2(n_2120),
.B(n_2099),
.C(n_2098),
.Y(n_2263)
);

O2A1O1Ixp33_ASAP7_75t_SL g2264 ( 
.A1(n_2245),
.A2(n_2098),
.B(n_2007),
.C(n_2036),
.Y(n_2264)
);

AOI221xp5_ASAP7_75t_L g2265 ( 
.A1(n_2247),
.A2(n_2098),
.B1(n_2018),
.B2(n_2017),
.C(n_2011),
.Y(n_2265)
);

CKINVDCx14_ASAP7_75t_R g2266 ( 
.A(n_2254),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2260),
.B(n_2237),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2262),
.B(n_2237),
.Y(n_2268)
);

XNOR2x1_ASAP7_75t_L g2269 ( 
.A(n_2250),
.B(n_2237),
.Y(n_2269)
);

OAI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2257),
.A2(n_2240),
.B1(n_2239),
.B2(n_2242),
.Y(n_2270)
);

NAND2xp33_ASAP7_75t_R g2271 ( 
.A(n_2252),
.B(n_2242),
.Y(n_2271)
);

INVx2_ASAP7_75t_SL g2272 ( 
.A(n_2258),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2255),
.A2(n_2251),
.B(n_2259),
.Y(n_2273)
);

OAI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2256),
.A2(n_2017),
.B1(n_2006),
.B2(n_2048),
.Y(n_2274)
);

BUFx2_ASAP7_75t_L g2275 ( 
.A(n_2272),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2268),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2266),
.B(n_2253),
.Y(n_2277)
);

INVxp67_ASAP7_75t_L g2278 ( 
.A(n_2271),
.Y(n_2278)
);

OAI211xp5_ASAP7_75t_SL g2279 ( 
.A1(n_2273),
.A2(n_2263),
.B(n_2261),
.C(n_2264),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2270),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2267),
.B(n_2265),
.Y(n_2281)
);

OAI211xp5_ASAP7_75t_L g2282 ( 
.A1(n_2269),
.A2(n_2265),
.B(n_1853),
.C(n_1879),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2275),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2277),
.Y(n_2284)
);

NOR3xp33_ASAP7_75t_L g2285 ( 
.A(n_2278),
.B(n_2274),
.C(n_1853),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2280),
.B(n_2048),
.Y(n_2286)
);

AOI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2279),
.A2(n_2034),
.B1(n_2029),
.B2(n_1899),
.Y(n_2287)
);

NOR3x1_ASAP7_75t_L g2288 ( 
.A(n_2281),
.B(n_1854),
.C(n_1851),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2283),
.B(n_2276),
.Y(n_2289)
);

AOI221xp5_ASAP7_75t_L g2290 ( 
.A1(n_2285),
.A2(n_2282),
.B1(n_1899),
.B2(n_2020),
.C(n_1998),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2284),
.Y(n_2291)
);

BUFx2_ASAP7_75t_L g2292 ( 
.A(n_2287),
.Y(n_2292)
);

AOI31xp33_ASAP7_75t_L g2293 ( 
.A1(n_2289),
.A2(n_2286),
.A3(n_2282),
.B(n_2288),
.Y(n_2293)
);

OA22x2_ASAP7_75t_L g2294 ( 
.A1(n_2291),
.A2(n_1875),
.B1(n_2020),
.B2(n_1998),
.Y(n_2294)
);

NOR2x1_ASAP7_75t_L g2295 ( 
.A(n_2293),
.B(n_2292),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2295),
.B(n_2290),
.Y(n_2296)
);

OR3x2_ASAP7_75t_L g2297 ( 
.A(n_2295),
.B(n_2294),
.C(n_1854),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2296),
.Y(n_2298)
);

AOI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_2297),
.A2(n_2046),
.B1(n_1899),
.B2(n_1853),
.Y(n_2299)
);

OAI222xp33_ASAP7_75t_L g2300 ( 
.A1(n_2298),
.A2(n_2046),
.B1(n_1851),
.B2(n_1854),
.C1(n_1894),
.C2(n_1889),
.Y(n_2300)
);

A2O1A1Ixp33_ASAP7_75t_L g2301 ( 
.A1(n_2299),
.A2(n_1832),
.B(n_1840),
.C(n_1852),
.Y(n_2301)
);

OAI22xp33_ASAP7_75t_L g2302 ( 
.A1(n_2301),
.A2(n_1851),
.B1(n_1881),
.B2(n_1893),
.Y(n_2302)
);

AOI221xp5_ASAP7_75t_L g2303 ( 
.A1(n_2302),
.A2(n_2300),
.B1(n_1840),
.B2(n_1852),
.C(n_1832),
.Y(n_2303)
);

AOI211xp5_ASAP7_75t_L g2304 ( 
.A1(n_2303),
.A2(n_1889),
.B(n_1894),
.C(n_1847),
.Y(n_2304)
);


endmodule