module real_jpeg_1797_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_1),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_1),
.B(n_19),
.C(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_1),
.A2(n_18),
.B1(n_29),
.B2(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_1),
.B(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_1),
.A2(n_18),
.B1(n_41),
.B2(n_61),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_1),
.B(n_27),
.C(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_1),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_1),
.B(n_48),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_1),
.B(n_23),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_19),
.B1(n_22),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_4),
.A2(n_37),
.B1(n_41),
.B2(n_61),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_4),
.A2(n_29),
.B1(n_32),
.B2(n_37),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_5),
.A2(n_29),
.B1(n_32),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_5),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_5),
.A2(n_41),
.B1(n_61),
.B2(n_69),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_5),
.A2(n_19),
.B1(n_22),
.B2(n_69),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_96),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_94),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_81),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_13),
.B(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_80),
.Y(n_13)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_38),
.B1(n_50),
.B2(n_51),
.Y(n_14)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_33),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_23),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_17),
.B(n_34),
.Y(n_104)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_19),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_19),
.A2(n_22),
.B1(n_44),
.B2(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_19),
.B(n_102),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_23),
.B(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_25),
.B(n_85),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_29),
.B(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_33),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_34),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_45),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_39),
.A2(n_40),
.B1(n_45),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_57)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_44),
.B1(n_61),
.B2(n_73),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B(n_49),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_111),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_46),
.B(n_68),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_47),
.B(n_111),
.Y(n_126)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_48),
.B(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_70),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_65),
.B(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_67),
.B(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.C(n_92),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_86),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_139),
.B(n_143),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_120),
.B(n_138),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_112),
.B1(n_113),
.B2(n_119),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_117),
.C(n_119),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_128),
.B(n_137),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_133),
.B(n_136),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_141),
.Y(n_143)
);


endmodule