module fake_jpeg_24574_n_286 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_37),
.Y(n_66)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_35),
.B1(n_27),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_35),
.B1(n_32),
.B2(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_32),
.B1(n_18),
.B2(n_21),
.Y(n_52)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_31),
.B1(n_32),
.B2(n_21),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_32),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_73),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_32),
.B1(n_18),
.B2(n_21),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_68),
.B1(n_80),
.B2(n_2),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_66),
.B(n_74),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_18),
.B1(n_37),
.B2(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_77),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_18),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_81),
.C(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_26),
.Y(n_71)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_33),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_22),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_33),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_28),
.B1(n_22),
.B2(n_20),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_23),
.B1(n_36),
.B2(n_24),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_28),
.B1(n_30),
.B2(n_34),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_34),
.B(n_30),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_23),
.C(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_87),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_39),
.B(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_19),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_29),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_49),
.B1(n_80),
.B2(n_84),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_36),
.B1(n_29),
.B2(n_4),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_115),
.B1(n_67),
.B2(n_63),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_1),
.Y(n_101)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_2),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_110),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_49),
.B1(n_53),
.B2(n_10),
.Y(n_146)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_62),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_5),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_6),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_63),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_53),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_6),
.B(n_7),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_64),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_114),
.B1(n_111),
.B2(n_105),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_118),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_125),
.Y(n_165)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_51),
.B(n_80),
.C(n_70),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_132),
.B(n_148),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_127),
.A2(n_131),
.B(n_8),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_62),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_136),
.B1(n_146),
.B2(n_120),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_80),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_85),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_9),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_54),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_99),
.B(n_61),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_61),
.B(n_76),
.C(n_78),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_69),
.B1(n_83),
.B2(n_55),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_149),
.A2(n_116),
.B1(n_120),
.B2(n_106),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_69),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_95),
.C(n_90),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_8),
.Y(n_151)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_159),
.B1(n_173),
.B2(n_177),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_163),
.A2(n_171),
.B1(n_178),
.B2(n_182),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_128),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_129),
.B(n_137),
.CI(n_130),
.CON(n_167),
.SN(n_167)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_167),
.B(n_174),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_90),
.C(n_91),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_126),
.A2(n_96),
.B1(n_117),
.B2(n_109),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_99),
.B1(n_119),
.B2(n_91),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_113),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_180),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_148),
.A2(n_112),
.B1(n_92),
.B2(n_55),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_124),
.A2(n_103),
.B(n_112),
.Y(n_178)
);

AOI22x1_ASAP7_75t_L g181 ( 
.A1(n_132),
.A2(n_103),
.B1(n_10),
.B2(n_11),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_138),
.B1(n_11),
.B2(n_12),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_121),
.A2(n_92),
.B1(n_103),
.B2(n_12),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_129),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_197),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_141),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_125),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_149),
.B(n_132),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_202),
.B(n_182),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_193),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_127),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_168),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_122),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_143),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_203),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_162),
.A2(n_152),
.B1(n_134),
.B2(n_147),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_155),
.B1(n_181),
.B2(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_176),
.B(n_153),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_206),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_9),
.B(n_11),
.C(n_13),
.D(n_14),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_173),
.C(n_153),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_138),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_200),
.B(n_199),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_221),
.B(n_225),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_167),
.C(n_178),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_171),
.Y(n_215)
);

OA21x2_ASAP7_75t_SL g221 ( 
.A1(n_201),
.A2(n_167),
.B(n_163),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_222),
.C(n_224),
.Y(n_230)
);

OA21x2_ASAP7_75t_SL g222 ( 
.A1(n_192),
.A2(n_157),
.B(n_179),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_202),
.Y(n_228)
);

OAI322xp33_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_174),
.A3(n_161),
.B1(n_164),
.B2(n_160),
.C1(n_158),
.C2(n_15),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_161),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_227),
.C(n_185),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_158),
.C(n_164),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_223),
.B(n_219),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_208),
.B1(n_220),
.B2(n_213),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_207),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_240),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_188),
.B(n_203),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_243),
.B(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_235),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_234),
.B(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_238),
.C(n_242),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_194),
.C(n_199),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_194),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_197),
.CI(n_190),
.CON(n_241),
.SN(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_186),
.C(n_190),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_242),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_236),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_231),
.A2(n_209),
.B1(n_210),
.B2(n_217),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_227),
.B1(n_210),
.B2(n_240),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_212),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_237),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_251),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_249),
.A2(n_257),
.B(n_256),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_250),
.B(n_255),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_218),
.Y(n_251)
);

AOI31xp67_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_220),
.A3(n_224),
.B(n_205),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_230),
.B(n_236),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_266),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_264),
.C(n_265),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_244),
.B(n_246),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_250),
.B1(n_246),
.B2(n_14),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_193),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_13),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_254),
.B(n_247),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_268),
.A2(n_269),
.B(n_261),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_263),
.B(n_254),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_253),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_270),
.B(n_273),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_277),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_266),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_264),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_280),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_276),
.A2(n_271),
.B(n_260),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_279),
.C(n_258),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_282),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_283),
.Y(n_286)
);


endmodule