module fake_ibex_347_n_812 (n_85, n_128, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_91, n_54, n_19, n_812);

input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_812;

wire n_151;
wire n_599;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_144;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_732;
wire n_673;
wire n_798;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_791;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_141;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_772;
wire n_810;
wire n_768;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_721;
wire n_365;
wire n_651;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_562;
wire n_564;
wire n_506;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_159;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_60),
.Y(n_146)
);

INVx4_ASAP7_75t_R g147 ( 
.A(n_99),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_102),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_1),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_57),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_48),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_19),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_50),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_56),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_37),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_3),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_61),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_38),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_63),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_46),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_4),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_41),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_47),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_14),
.B(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_40),
.Y(n_176)
);

BUFx2_ASAP7_75t_SL g177 ( 
.A(n_100),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_0),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_89),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_27),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_36),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_53),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_71),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_72),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_90),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_18),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_54),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_91),
.B(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_7),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_55),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_51),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_22),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_29),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_59),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_62),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_32),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_8),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_96),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_67),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_76),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_92),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_58),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_52),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_1),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_78),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_94),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_75),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_49),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_19),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_85),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_25),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_66),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_73),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_64),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_9),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_95),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_113),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_10),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_74),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_111),
.B(n_88),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_83),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_81),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_39),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_77),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_21),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_34),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_9),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_65),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_136),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_80),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_97),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_164),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_160),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_164),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_171),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_160),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_4),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_5),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g254 ( 
.A(n_191),
.B(n_30),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_214),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_156),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_6),
.Y(n_258)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_150),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_150),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_163),
.Y(n_262)
);

AND2x6_ASAP7_75t_L g263 ( 
.A(n_158),
.B(n_31),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_142),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_143),
.Y(n_266)
);

NOR2x1_ASAP7_75t_L g267 ( 
.A(n_144),
.B(n_33),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_178),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_190),
.B(n_11),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_190),
.B(n_11),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_158),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_183),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_168),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_195),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_205),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_168),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_195),
.B(n_12),
.Y(n_279)
);

OA21x2_ASAP7_75t_L g280 ( 
.A1(n_201),
.A2(n_69),
.B(n_140),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_206),
.B(n_13),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_149),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_209),
.B(n_13),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_206),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_207),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_207),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_202),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_145),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_218),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_151),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_152),
.Y(n_294)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_176),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_180),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_153),
.A2(n_155),
.B(n_154),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_157),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_159),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_161),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g301 ( 
.A1(n_162),
.A2(n_70),
.B(n_137),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_166),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_169),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_194),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_170),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_172),
.B(n_17),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_175),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_306),
.B(n_302),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_239),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_186),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_240),
.B(n_165),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_296),
.Y(n_317)
);

AOI21x1_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_193),
.B(n_187),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_253),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_272),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_254),
.A2(n_224),
.B1(n_237),
.B2(n_167),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_295),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_196),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_302),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_242),
.B(n_215),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_263),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_295),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_293),
.B(n_203),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_305),
.B(n_204),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_211),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_287),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

BUFx6f_ASAP7_75t_SL g339 ( 
.A(n_254),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_305),
.B(n_213),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_263),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_247),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_245),
.Y(n_344)
);

OR2x6_ASAP7_75t_L g345 ( 
.A(n_269),
.B(n_177),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_289),
.B(n_227),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_245),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_220),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_239),
.Y(n_349)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_255),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_307),
.B(n_226),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_285),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_249),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_276),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_265),
.B(n_266),
.Y(n_356)
);

INVx5_ASAP7_75t_L g357 ( 
.A(n_263),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_249),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_277),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_290),
.B(n_228),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_278),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_298),
.B(n_229),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_255),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_255),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_300),
.B(n_231),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_262),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_303),
.B(n_233),
.Y(n_367)
);

AO21x2_ASAP7_75t_L g368 ( 
.A1(n_279),
.A2(n_174),
.B(n_236),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_278),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_239),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_246),
.B(n_271),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_273),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_294),
.B(n_192),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_273),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_281),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_L g376 ( 
.A1(n_270),
.A2(n_210),
.B1(n_221),
.B2(n_217),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_294),
.B(n_141),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_252),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_275),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_257),
.B(n_146),
.Y(n_380)
);

INVx8_ASAP7_75t_L g381 ( 
.A(n_284),
.Y(n_381)
);

AND2x2_ASAP7_75t_SL g382 ( 
.A(n_280),
.B(n_147),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_299),
.B(n_148),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_317),
.B(n_258),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_297),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_382),
.A2(n_297),
.B(n_280),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_309),
.B(n_264),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_260),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_339),
.A2(n_222),
.B1(n_173),
.B2(n_219),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_378),
.A2(n_282),
.B1(n_261),
.B2(n_274),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_311),
.B(n_244),
.Y(n_391)
);

BUFx8_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_380),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_327),
.B(n_328),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_L g397 ( 
.A(n_314),
.B(n_350),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_292),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_338),
.B(n_292),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_350),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

OR2x6_ASAP7_75t_L g403 ( 
.A(n_345),
.B(n_267),
.Y(n_403)
);

OR2x6_ASAP7_75t_L g404 ( 
.A(n_345),
.B(n_280),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

OR2x6_ASAP7_75t_L g406 ( 
.A(n_345),
.B(n_301),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_363),
.Y(n_407)
);

OR2x6_ASAP7_75t_L g408 ( 
.A(n_322),
.B(n_301),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_353),
.B(n_284),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_315),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_339),
.A2(n_338),
.B1(n_314),
.B2(n_376),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_326),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_371),
.A2(n_288),
.B1(n_216),
.B2(n_212),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_343),
.Y(n_415)
);

OR2x6_ASAP7_75t_L g416 ( 
.A(n_323),
.B(n_301),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_373),
.B(n_179),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_344),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_314),
.A2(n_225),
.B1(n_182),
.B2(n_185),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_357),
.B(n_181),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_343),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_379),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_354),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_313),
.A2(n_288),
.B1(n_235),
.B2(n_223),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_316),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_359),
.B(n_188),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_324),
.B(n_199),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_357),
.B(n_200),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_319),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_324),
.Y(n_432)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_366),
.Y(n_435)
);

A2O1A1Ixp33_ASAP7_75t_L g436 ( 
.A1(n_360),
.A2(n_248),
.B(n_256),
.C(n_251),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_321),
.Y(n_438)
);

OAI221xp5_ASAP7_75t_L g439 ( 
.A1(n_365),
.A2(n_259),
.B1(n_243),
.B2(n_251),
.C(n_250),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_331),
.B(n_243),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_336),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_352),
.B(n_241),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_352),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_356),
.B(n_241),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_367),
.B(n_241),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_362),
.A2(n_256),
.B1(n_251),
.B2(n_250),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_377),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_386),
.A2(n_318),
.B(n_308),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_335),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_362),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_377),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_383),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_437),
.A2(n_340),
.B1(n_334),
.B2(n_333),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_385),
.A2(n_381),
.B(n_372),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_384),
.B(n_337),
.Y(n_455)
);

AO21x1_ASAP7_75t_L g456 ( 
.A1(n_398),
.A2(n_325),
.B(n_329),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_434),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_387),
.B(n_341),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_396),
.A2(n_397),
.B(n_428),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_411),
.B(n_35),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_392),
.Y(n_461)
);

AO21x1_ASAP7_75t_L g462 ( 
.A1(n_445),
.A2(n_355),
.B(n_375),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_400),
.B(n_20),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_391),
.B(n_20),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_393),
.B(n_21),
.Y(n_466)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_415),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_401),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_22),
.Y(n_469)
);

AO21x1_ASAP7_75t_L g470 ( 
.A1(n_442),
.A2(n_361),
.B(n_369),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_416),
.A2(n_330),
.B(n_332),
.Y(n_471)
);

O2A1O1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_413),
.A2(n_346),
.B(n_24),
.C(n_25),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_421),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_416),
.A2(n_370),
.B(n_349),
.Y(n_474)
);

OAI21xp33_ASAP7_75t_L g475 ( 
.A1(n_417),
.A2(n_256),
.B(n_250),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_416),
.A2(n_370),
.B(n_349),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_399),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_418),
.B(n_23),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_427),
.B(n_24),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_410),
.B(n_26),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_395),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_422),
.B(n_27),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_424),
.B(n_28),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_388),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_419),
.B(n_390),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_408),
.A2(n_370),
.B1(n_349),
.B2(n_310),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_29),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_401),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_402),
.Y(n_490)
);

O2A1O1Ixp33_ASAP7_75t_SL g491 ( 
.A1(n_444),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_403),
.B(n_45),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_435),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_409),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_423),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_394),
.Y(n_497)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_408),
.B(n_425),
.C(n_404),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_403),
.B(n_133),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

OA22x2_ASAP7_75t_L g501 ( 
.A1(n_403),
.A2(n_408),
.B1(n_389),
.B2(n_404),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_414),
.A2(n_82),
.B(n_84),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_455),
.B(n_440),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_474),
.A2(n_420),
.B(n_430),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_438),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_436),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_461),
.B(n_431),
.Y(n_509)
);

NAND2x1_ASAP7_75t_L g510 ( 
.A(n_468),
.B(n_446),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_473),
.B(n_439),
.Y(n_511)
);

BUFx10_ASAP7_75t_L g512 ( 
.A(n_492),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_451),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_463),
.Y(n_514)
);

AO21x1_ASAP7_75t_L g515 ( 
.A1(n_504),
.A2(n_426),
.B(n_98),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_448),
.A2(n_459),
.B(n_454),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_464),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_465),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_479),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_450),
.B(n_103),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_468),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_484),
.Y(n_523)
);

A2O1A1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_460),
.A2(n_105),
.B(n_107),
.C(n_109),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_452),
.Y(n_525)
);

AO31x2_ASAP7_75t_L g526 ( 
.A1(n_456),
.A2(n_110),
.A3(n_115),
.B(n_116),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_458),
.B(n_121),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_457),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_480),
.B(n_122),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_501),
.B(n_123),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_476),
.A2(n_124),
.B(n_127),
.Y(n_531)
);

NOR2x1_ASAP7_75t_SL g532 ( 
.A(n_502),
.B(n_503),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_466),
.B(n_457),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_488),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_478),
.B(n_496),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_469),
.B(n_494),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_481),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_482),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_453),
.B(n_497),
.Y(n_539)
);

OAI22x1_ASAP7_75t_L g540 ( 
.A1(n_498),
.A2(n_499),
.B1(n_477),
.B2(n_500),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_490),
.B(n_495),
.Y(n_541)
);

BUFx8_ASAP7_75t_L g542 ( 
.A(n_503),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_489),
.Y(n_543)
);

NAND2x1p5_ASAP7_75t_L g544 ( 
.A(n_489),
.B(n_503),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_475),
.Y(n_545)
);

OAI21x1_ASAP7_75t_SL g546 ( 
.A1(n_491),
.A2(n_499),
.B(n_504),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_449),
.B(n_433),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_449),
.B(n_433),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_492),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_455),
.B(n_432),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_455),
.B(n_432),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_448),
.A2(n_386),
.B(n_385),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_455),
.B(n_432),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_493),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_455),
.A2(n_432),
.B1(n_443),
.B2(n_441),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_449),
.B(n_433),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_455),
.B(n_432),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_455),
.B(n_432),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_SL g559 ( 
.A(n_472),
.B(n_359),
.C(n_317),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_493),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_493),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_448),
.A2(n_386),
.B(n_385),
.Y(n_562)
);

AO31x2_ASAP7_75t_L g563 ( 
.A1(n_456),
.A2(n_470),
.A3(n_462),
.B(n_386),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_461),
.Y(n_564)
);

CKINVDCx8_ASAP7_75t_R g565 ( 
.A(n_467),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_449),
.B(n_433),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_455),
.B(n_432),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_468),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_455),
.B(n_432),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_455),
.B(n_432),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_449),
.B(n_433),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_493),
.Y(n_572)
);

AOI221x1_ASAP7_75t_L g573 ( 
.A1(n_498),
.A2(n_474),
.B1(n_471),
.B2(n_476),
.C(n_386),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_448),
.A2(n_396),
.B(n_342),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_461),
.Y(n_575)
);

INVx4_ASAP7_75t_SL g576 ( 
.A(n_461),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_492),
.Y(n_577)
);

OA21x2_ASAP7_75t_L g578 ( 
.A1(n_476),
.A2(n_386),
.B(n_448),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_455),
.A2(n_432),
.B1(n_443),
.B2(n_441),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_455),
.B(n_432),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_461),
.Y(n_581)
);

AO21x2_ASAP7_75t_L g582 ( 
.A1(n_476),
.A2(n_498),
.B(n_487),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_478),
.Y(n_583)
);

AOI211x1_ASAP7_75t_L g584 ( 
.A1(n_465),
.A2(n_466),
.B(n_464),
.C(n_486),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_550),
.B(n_551),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_553),
.B(n_557),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_542),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_547),
.Y(n_588)
);

CKINVDCx11_ASAP7_75t_R g589 ( 
.A(n_576),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_558),
.B(n_567),
.Y(n_590)
);

AO21x2_ASAP7_75t_L g591 ( 
.A1(n_552),
.A2(n_562),
.B(n_546),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_530),
.B(n_548),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_556),
.B(n_566),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_569),
.B(n_570),
.Y(n_594)
);

AO31x2_ASAP7_75t_L g595 ( 
.A1(n_515),
.A2(n_545),
.A3(n_539),
.B(n_574),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_571),
.B(n_580),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_579),
.B(n_513),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_542),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_554),
.B(n_560),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_525),
.A2(n_505),
.B(n_518),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_517),
.A2(n_534),
.B(n_519),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_530),
.B(n_564),
.Y(n_602)
);

OA21x2_ASAP7_75t_L g603 ( 
.A1(n_531),
.A2(n_527),
.B(n_506),
.Y(n_603)
);

OA21x2_ASAP7_75t_L g604 ( 
.A1(n_524),
.A2(n_520),
.B(n_522),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_578),
.A2(n_510),
.B(n_544),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_561),
.B(n_572),
.Y(n_606)
);

NAND2x1p5_ASAP7_75t_L g607 ( 
.A(n_575),
.B(n_543),
.Y(n_607)
);

CKINVDCx16_ASAP7_75t_R g608 ( 
.A(n_514),
.Y(n_608)
);

BUFx2_ASAP7_75t_R g609 ( 
.A(n_581),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_565),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_583),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_535),
.B(n_523),
.Y(n_612)
);

AO21x2_ASAP7_75t_L g613 ( 
.A1(n_582),
.A2(n_529),
.B(n_508),
.Y(n_613)
);

AO31x2_ASAP7_75t_L g614 ( 
.A1(n_563),
.A2(n_532),
.A3(n_533),
.B(n_584),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_559),
.B(n_537),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_538),
.Y(n_616)
);

OR2x6_ASAP7_75t_L g617 ( 
.A(n_509),
.B(n_528),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_541),
.B(n_577),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_507),
.A2(n_536),
.B(n_511),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_563),
.Y(n_620)
);

BUFx2_ASAP7_75t_R g621 ( 
.A(n_576),
.Y(n_621)
);

NAND2x1p5_ASAP7_75t_L g622 ( 
.A(n_521),
.B(n_568),
.Y(n_622)
);

BUFx2_ASAP7_75t_R g623 ( 
.A(n_512),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_526),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_512),
.B(n_549),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_577),
.B(n_549),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_530),
.B(n_461),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_550),
.B(n_551),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_583),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_542),
.Y(n_630)
);

NAND2x1p5_ASAP7_75t_L g631 ( 
.A(n_564),
.B(n_461),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_583),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_581),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_550),
.B(n_412),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_530),
.B(n_547),
.Y(n_635)
);

NAND2x1p5_ASAP7_75t_L g636 ( 
.A(n_564),
.B(n_461),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_583),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_550),
.B(n_412),
.Y(n_638)
);

AO31x2_ASAP7_75t_L g639 ( 
.A1(n_515),
.A2(n_573),
.A3(n_516),
.B(n_540),
.Y(n_639)
);

NOR2x1_ASAP7_75t_R g640 ( 
.A(n_581),
.B(n_461),
.Y(n_640)
);

CKINVDCx6p67_ASAP7_75t_R g641 ( 
.A(n_564),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_550),
.B(n_551),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_583),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_550),
.B(n_551),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_547),
.B(n_548),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_555),
.A2(n_579),
.B1(n_501),
.B2(n_530),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_564),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_611),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_611),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_627),
.A2(n_602),
.B1(n_646),
.B2(n_592),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_617),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_602),
.B(n_627),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_617),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_629),
.B(n_632),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_632),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_637),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_643),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_643),
.B(n_616),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_620),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_594),
.B(n_585),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_586),
.A2(n_628),
.B(n_642),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_614),
.B(n_605),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_641),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_597),
.B(n_601),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_587),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_614),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_608),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_614),
.Y(n_668)
);

BUFx12f_ASAP7_75t_L g669 ( 
.A(n_589),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_590),
.B(n_644),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_622),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_634),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_612),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_624),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_608),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_588),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_596),
.B(n_646),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_592),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_635),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_591),
.Y(n_680)
);

AO21x2_ASAP7_75t_L g681 ( 
.A1(n_613),
.A2(n_600),
.B(n_619),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_599),
.Y(n_682)
);

AO21x2_ASAP7_75t_L g683 ( 
.A1(n_639),
.A2(n_595),
.B(n_615),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_593),
.B(n_645),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_618),
.B(n_606),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_639),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_647),
.Y(n_687)
);

AO21x1_ASAP7_75t_SL g688 ( 
.A1(n_626),
.A2(n_610),
.B(n_621),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_638),
.B(n_604),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_630),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_607),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_683),
.B(n_659),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_664),
.B(n_595),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_674),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_683),
.B(n_603),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_652),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_664),
.B(n_625),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_662),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_659),
.B(n_598),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_658),
.B(n_631),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_658),
.B(n_636),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_671),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_654),
.B(n_623),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_648),
.B(n_640),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_689),
.Y(n_705)
);

OAI221xp5_ASAP7_75t_L g706 ( 
.A1(n_650),
.A2(n_609),
.B1(n_633),
.B2(n_640),
.C(n_661),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_677),
.B(n_681),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_666),
.B(n_668),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_652),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_662),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_654),
.B(n_648),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_654),
.B(n_649),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_655),
.B(n_657),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_656),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_652),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_705),
.B(n_689),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_700),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_711),
.B(n_666),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_711),
.B(n_681),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_714),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_707),
.B(n_660),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_712),
.B(n_680),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_710),
.B(n_662),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_699),
.B(n_697),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_702),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_713),
.Y(n_726)
);

OR2x6_ASAP7_75t_SL g727 ( 
.A(n_704),
.B(n_690),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_713),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_692),
.B(n_680),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_692),
.B(n_686),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_694),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_719),
.B(n_692),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_719),
.B(n_698),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_731),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_729),
.B(n_698),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_726),
.B(n_697),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_727),
.A2(n_706),
.B1(n_652),
.B2(n_696),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_729),
.B(n_708),
.Y(n_738)
);

NAND3xp33_ASAP7_75t_L g739 ( 
.A(n_720),
.B(n_704),
.C(n_706),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_725),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_730),
.B(n_708),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_730),
.B(n_708),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_718),
.B(n_693),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_723),
.B(n_695),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_718),
.B(n_693),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_723),
.B(n_695),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_738),
.B(n_741),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_739),
.B(n_727),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_741),
.B(n_721),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_738),
.B(n_728),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_742),
.B(n_716),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_740),
.Y(n_752)
);

NOR2x1_ASAP7_75t_L g753 ( 
.A(n_737),
.B(n_652),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_732),
.B(n_716),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_736),
.B(n_687),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_734),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_742),
.B(n_721),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_743),
.B(n_724),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_743),
.B(n_722),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_734),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_752),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_756),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_748),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_748),
.A2(n_703),
.B(n_675),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_753),
.A2(n_746),
.B1(n_744),
.B2(n_703),
.Y(n_765)
);

OAI21xp33_ASAP7_75t_L g766 ( 
.A1(n_752),
.A2(n_735),
.B(n_733),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_749),
.A2(n_740),
.B1(n_746),
.B2(n_744),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_747),
.B(n_690),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_760),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_754),
.B(n_732),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_757),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_758),
.B(n_745),
.Y(n_772)
);

AOI211xp5_ASAP7_75t_L g773 ( 
.A1(n_764),
.A2(n_663),
.B(n_755),
.C(n_667),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_761),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_769),
.Y(n_775)
);

AOI32xp33_ASAP7_75t_L g776 ( 
.A1(n_768),
.A2(n_755),
.A3(n_754),
.B1(n_751),
.B2(n_759),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_767),
.A2(n_750),
.B(n_744),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_762),
.Y(n_778)
);

OAI21xp33_ASAP7_75t_L g779 ( 
.A1(n_776),
.A2(n_763),
.B(n_764),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_SL g780 ( 
.A(n_773),
.B(n_765),
.C(n_766),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_777),
.B(n_669),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_779),
.A2(n_774),
.B1(n_775),
.B2(n_778),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_780),
.B(n_781),
.C(n_665),
.Y(n_783)
);

OR2x6_ASAP7_75t_L g784 ( 
.A(n_783),
.B(n_669),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_782),
.B(n_772),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_785),
.B(n_770),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_784),
.B(n_771),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_787),
.A2(n_665),
.B1(n_696),
.B2(n_672),
.Y(n_788)
);

AND4x1_ASAP7_75t_L g789 ( 
.A(n_786),
.B(n_688),
.C(n_684),
.D(n_701),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_788),
.Y(n_790)
);

AOI211x1_ASAP7_75t_L g791 ( 
.A1(n_789),
.A2(n_684),
.B(n_688),
.C(n_701),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_788),
.Y(n_792)
);

XOR2xp5_ASAP7_75t_L g793 ( 
.A(n_792),
.B(n_660),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_790),
.B(n_676),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_791),
.A2(n_696),
.B1(n_709),
.B2(n_715),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_792),
.Y(n_796)
);

AND2x2_ASAP7_75t_SL g797 ( 
.A(n_790),
.B(n_670),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_796),
.A2(n_651),
.B(n_653),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_793),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_797),
.A2(n_651),
.B1(n_653),
.B2(n_696),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_SL g801 ( 
.A(n_794),
.B(n_670),
.C(n_679),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_795),
.A2(n_691),
.B(n_673),
.Y(n_802)
);

XNOR2xp5_ASAP7_75t_L g803 ( 
.A(n_793),
.B(n_685),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_798),
.A2(n_691),
.B(n_673),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_799),
.A2(n_691),
.B(n_685),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_800),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_SL g807 ( 
.A1(n_803),
.A2(n_678),
.B1(n_682),
.B2(n_709),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_806),
.A2(n_801),
.B(n_802),
.Y(n_808)
);

AOI221xp5_ASAP7_75t_L g809 ( 
.A1(n_805),
.A2(n_682),
.B1(n_678),
.B2(n_679),
.C(n_715),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_804),
.A2(n_717),
.B(n_700),
.Y(n_810)
);

OR2x6_ASAP7_75t_L g811 ( 
.A(n_808),
.B(n_807),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_SL g812 ( 
.A1(n_811),
.A2(n_810),
.B1(n_809),
.B2(n_678),
.Y(n_812)
);


endmodule