module fake_jpeg_1978_n_571 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_571);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_571;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_53),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_54),
.B(n_70),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_18),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_24),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_61),
.B(n_77),
.Y(n_120)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_99),
.Y(n_119)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_35),
.B(n_0),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_26),
.Y(n_88)
);

BUFx24_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_41),
.B(n_16),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_106),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_29),
.Y(n_90)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_58),
.Y(n_134)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_55),
.A2(n_80),
.B1(n_81),
.B2(n_101),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_109),
.A2(n_82),
.B1(n_96),
.B2(n_95),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_64),
.A2(n_52),
.B1(n_37),
.B2(n_51),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_126),
.A2(n_130),
.B1(n_40),
.B2(n_88),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_67),
.A2(n_52),
.B1(n_37),
.B2(n_51),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_75),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_133),
.B(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_134),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_41),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_65),
.B(n_42),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_141),
.B(n_143),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_72),
.B(n_42),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_76),
.B(n_48),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_154),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_102),
.A2(n_52),
.B1(n_30),
.B2(n_19),
.Y(n_153)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_153),
.A2(n_39),
.B1(n_22),
.B2(n_28),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_48),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_43),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_156),
.B(n_163),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_98),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_166),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_92),
.A2(n_40),
.B1(n_34),
.B2(n_32),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_158),
.A2(n_93),
.B1(n_40),
.B2(n_34),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_53),
.B(n_43),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_78),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_86),
.B(n_50),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_168),
.B(n_0),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_79),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_131),
.Y(n_176)
);

CKINVDCx9p33_ASAP7_75t_R g172 ( 
.A(n_116),
.Y(n_172)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

BUFx12_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_174),
.Y(n_234)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_175),
.Y(n_251)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_177),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_178),
.Y(n_260)
);

CKINVDCx9p33_ASAP7_75t_R g179 ( 
.A(n_116),
.Y(n_179)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_179),
.Y(n_258)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_181),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_182),
.A2(n_216),
.B1(n_225),
.B2(n_121),
.Y(n_284)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_139),
.A2(n_94),
.B1(n_83),
.B2(n_32),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_185),
.A2(n_186),
.B1(n_130),
.B2(n_132),
.Y(n_248)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_91),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_202),
.Y(n_240)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_192),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_110),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_193),
.B(n_205),
.Y(n_244)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_195),
.Y(n_266)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_197),
.A2(n_220),
.B1(n_228),
.B2(n_233),
.Y(n_283)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_198),
.Y(n_279)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_199),
.Y(n_280)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_120),
.B(n_25),
.CI(n_73),
.CON(n_202),
.SN(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_112),
.Y(n_203)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_122),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_107),
.B(n_50),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_148),
.B(n_97),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_208),
.B(n_212),
.Y(n_255)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_111),
.B(n_32),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_211),
.B(n_227),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_114),
.B(n_84),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_110),
.A2(n_73),
.B(n_1),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_213),
.A2(n_162),
.B(n_164),
.Y(n_271)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_129),
.Y(n_214)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_214),
.Y(n_282)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_145),
.Y(n_215)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_215),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_161),
.A2(n_62),
.B1(n_31),
.B2(n_39),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_142),
.B(n_39),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_144),
.C(n_126),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_158),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_155),
.Y(n_223)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_147),
.Y(n_224)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_132),
.A2(n_22),
.B1(n_28),
.B2(n_25),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_153),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_137),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_231),
.Y(n_270)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_232),
.Y(n_275)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_109),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_153),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_237),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_171),
.B(n_226),
.C(n_184),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_243),
.B(n_277),
.Y(n_298)
);

OA22x2_ASAP7_75t_L g320 ( 
.A1(n_248),
.A2(n_196),
.B1(n_190),
.B2(n_140),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_171),
.A2(n_127),
.B1(n_144),
.B2(n_151),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_182),
.A2(n_138),
.B1(n_151),
.B2(n_150),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_264),
.A2(n_218),
.B1(n_160),
.B2(n_136),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_173),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_267),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_210),
.A2(n_164),
.B1(n_162),
.B2(n_169),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

NOR3xp33_ASAP7_75t_L g330 ( 
.A(n_271),
.B(n_286),
.C(n_174),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_150),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_285),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_122),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_213),
.A2(n_121),
.B(n_108),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_216),
.B(n_175),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_284),
.A2(n_180),
.B1(n_232),
.B2(n_201),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_189),
.B(n_149),
.Y(n_285)
);

NOR2x1_ASAP7_75t_SL g286 ( 
.A(n_202),
.B(n_218),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_178),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_287),
.B(n_5),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_240),
.A2(n_225),
.B(n_186),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_289),
.A2(n_301),
.B(n_330),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_290),
.Y(n_346)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_253),
.Y(n_292)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_244),
.B(n_204),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_294),
.B(n_308),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_264),
.A2(n_179),
.B1(n_172),
.B2(n_192),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_270),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_335),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_235),
.A2(n_194),
.B1(n_207),
.B2(n_198),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_234),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_299),
.Y(n_357)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_303),
.A2(n_317),
.B1(n_328),
.B2(n_337),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_200),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_327),
.Y(n_340)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_257),
.Y(n_305)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_265),
.Y(n_307)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_239),
.B(n_187),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_242),
.B(n_181),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_311),
.B(n_312),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_243),
.B(n_199),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_238),
.B(n_206),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_313),
.B(n_333),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_283),
.A2(n_286),
.B1(n_248),
.B2(n_235),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_314),
.A2(n_321),
.B1(n_323),
.B2(n_258),
.Y(n_343)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_252),
.Y(n_315)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_262),
.Y(n_316)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_251),
.Y(n_318)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_318),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_322),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_283),
.A2(n_149),
.B1(n_160),
.B2(n_136),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_288),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_235),
.A2(n_125),
.B1(n_177),
.B2(n_147),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_195),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_338),
.C(n_275),
.Y(n_350)
);

OA22x2_ASAP7_75t_L g325 ( 
.A1(n_269),
.A2(n_125),
.B1(n_147),
.B2(n_108),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_325),
.B(n_329),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_255),
.B(n_3),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_237),
.A2(n_275),
.B1(n_276),
.B2(n_271),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_272),
.B(n_7),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_332),
.Y(n_353)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_262),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_268),
.B(n_7),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_254),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_256),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_261),
.Y(n_335)
);

INVx11_ASAP7_75t_L g336 ( 
.A(n_250),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_336),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_266),
.A2(n_224),
.B1(n_174),
.B2(n_10),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g338 ( 
.A(n_281),
.B(n_7),
.C(n_8),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_301),
.A2(n_275),
.B(n_263),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_342),
.A2(n_364),
.B(n_366),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_343),
.A2(n_379),
.B1(n_319),
.B2(n_335),
.Y(n_384)
);

OAI21xp33_ASAP7_75t_L g402 ( 
.A1(n_350),
.A2(n_299),
.B(n_274),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_293),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_354),
.B(n_365),
.C(n_371),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_328),
.A2(n_254),
.B(n_256),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_298),
.B(n_273),
.C(n_282),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_293),
.A2(n_259),
.B(n_247),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_317),
.A2(n_246),
.B1(n_261),
.B2(n_278),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_370),
.A2(n_381),
.B1(n_258),
.B2(n_250),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_300),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_289),
.A2(n_249),
.B(n_247),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_372),
.A2(n_377),
.B(n_260),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_304),
.B(n_259),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_375),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_300),
.B(n_246),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_306),
.B(n_245),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_376),
.B(n_260),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_326),
.A2(n_288),
.B(n_236),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_314),
.A2(n_321),
.B1(n_326),
.B2(n_303),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_331),
.B(n_249),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_279),
.C(n_241),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_319),
.A2(n_278),
.B1(n_236),
.B2(n_280),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_291),
.B(n_279),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_334),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_347),
.B(n_306),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_383),
.B(n_389),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_384),
.A2(n_397),
.B1(n_400),
.B2(n_404),
.Y(n_448)
);

AO22x1_ASAP7_75t_L g386 ( 
.A1(n_362),
.A2(n_323),
.B1(n_325),
.B2(n_315),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_386),
.B(n_398),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_345),
.B(n_296),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_382),
.Y(n_391)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_391),
.Y(n_425)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_368),
.Y(n_392)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_392),
.Y(n_428)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_368),
.Y(n_393)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_393),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_354),
.B(n_338),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_394),
.B(n_353),
.C(n_372),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_346),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_395),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_396),
.B(n_416),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_379),
.A2(n_327),
.B1(n_320),
.B2(n_307),
.Y(n_397)
);

OAI32xp33_ASAP7_75t_L g398 ( 
.A1(n_375),
.A2(n_310),
.A3(n_302),
.B1(n_305),
.B2(n_292),
.Y(n_398)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_352),
.A2(n_339),
.B1(n_360),
.B2(n_342),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_402),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g403 ( 
.A(n_341),
.B(n_364),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_410),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_365),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_350),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_320),
.B1(n_325),
.B2(n_332),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_407),
.A2(n_343),
.B1(n_362),
.B2(n_378),
.Y(n_426)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_349),
.Y(n_408)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_316),
.Y(n_409)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_355),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_349),
.Y(n_411)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_411),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_360),
.A2(n_336),
.B1(n_325),
.B2(n_318),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_412),
.A2(n_370),
.B1(n_378),
.B2(n_339),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_351),
.B(n_274),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_413),
.Y(n_441)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_363),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_414),
.B(n_415),
.Y(n_445)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_363),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_357),
.B(n_241),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_377),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_251),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_361),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_366),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_381),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_421),
.B(n_449),
.C(n_415),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_423),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_426),
.A2(n_434),
.B1(n_439),
.B2(n_386),
.Y(n_473)
);

NOR2x1_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_340),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_436),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_429),
.A2(n_417),
.B(n_419),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_430),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_388),
.A2(n_362),
.B1(n_340),
.B2(n_341),
.Y(n_434)
);

NOR2x1_ASAP7_75t_L g436 ( 
.A(n_385),
.B(n_353),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_442),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_388),
.A2(n_344),
.B1(n_373),
.B2(n_348),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_386),
.B(n_356),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_447),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_394),
.B(n_361),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_387),
.B(n_369),
.C(n_359),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_369),
.Y(n_450)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_450),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_399),
.B(n_409),
.Y(n_451)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_451),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_387),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_453),
.B(n_455),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_405),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_406),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_458),
.B(n_474),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_435),
.B(n_410),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_461),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_436),
.B(n_390),
.Y(n_462)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_462),
.Y(n_491)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_445),
.Y(n_464)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_406),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_469),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_441),
.B(n_401),
.Y(n_466)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_466),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_467),
.B(n_476),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_432),
.Y(n_468)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_468),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_420),
.B(n_391),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_477),
.C(n_452),
.Y(n_495)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_472),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_473),
.A2(n_422),
.B1(n_443),
.B2(n_440),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_420),
.B(n_403),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_439),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_429),
.A2(n_407),
.B(n_404),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_424),
.B(n_414),
.C(n_411),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_408),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_450),
.Y(n_494)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_428),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_479),
.A2(n_480),
.B1(n_424),
.B2(n_431),
.Y(n_487)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_428),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_458),
.B(n_422),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_SL g512 ( 
.A(n_482),
.B(n_495),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_463),
.A2(n_426),
.B1(n_448),
.B2(n_432),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_483),
.A2(n_476),
.B1(n_500),
.B2(n_494),
.Y(n_514)
);

INVx11_ASAP7_75t_L g484 ( 
.A(n_470),
.Y(n_484)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_484),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_434),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_494),
.Y(n_505)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_487),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_492),
.A2(n_460),
.B1(n_478),
.B2(n_462),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_429),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_498),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_474),
.B(n_455),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_440),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_469),
.C(n_454),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_457),
.A2(n_423),
.B1(n_443),
.B2(n_425),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_473),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_506),
.B(n_521),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_500),
.A2(n_456),
.B(n_467),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_508),
.A2(n_518),
.B(n_499),
.Y(n_537)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_509),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_481),
.B(n_427),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_511),
.B(n_519),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_514),
.A2(n_488),
.B1(n_493),
.B2(n_482),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_454),
.C(n_477),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_516),
.C(n_489),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_489),
.B(n_456),
.C(n_425),
.Y(n_516)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_517),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_491),
.A2(n_447),
.B(n_446),
.Y(n_518)
);

AOI322xp5_ASAP7_75t_SL g519 ( 
.A1(n_503),
.A2(n_438),
.A3(n_367),
.B1(n_395),
.B2(n_444),
.C1(n_431),
.C2(n_452),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_502),
.A2(n_446),
.B1(n_444),
.B2(n_438),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_522),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_483),
.A2(n_393),
.B1(n_392),
.B2(n_346),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_504),
.A2(n_320),
.B1(n_359),
.B2(n_290),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_518),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_524),
.B(n_526),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_496),
.C(n_486),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_530),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_490),
.C(n_498),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_510),
.Y(n_531)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_531),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_533),
.A2(n_537),
.B(n_521),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_490),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_535),
.Y(n_550)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_523),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_485),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_538),
.B(n_485),
.C(n_505),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_520),
.B(n_497),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_539),
.A2(n_513),
.B1(n_517),
.B2(n_516),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_536),
.A2(n_512),
.B(n_508),
.Y(n_541)
);

AOI31xp67_ASAP7_75t_L g555 ( 
.A1(n_541),
.A2(n_530),
.A3(n_534),
.B(n_527),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_543),
.B(n_545),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_546),
.A2(n_547),
.B(n_548),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_528),
.A2(n_505),
.B(n_523),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_537),
.A2(n_522),
.B(n_484),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_525),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_549),
.B(n_539),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_526),
.C(n_529),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_551),
.B(n_553),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_544),
.A2(n_533),
.B(n_532),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_554),
.B(n_556),
.Y(n_558)
);

OAI211xp5_ASAP7_75t_L g559 ( 
.A1(n_555),
.A2(n_545),
.B(n_546),
.C(n_548),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_550),
.B(n_538),
.Y(n_556)
);

AOI21xp33_ASAP7_75t_L g563 ( 
.A1(n_559),
.A2(n_552),
.B(n_10),
.Y(n_563)
);

AOI322xp5_ASAP7_75t_L g560 ( 
.A1(n_557),
.A2(n_542),
.A3(n_532),
.B1(n_547),
.B2(n_527),
.C1(n_13),
.C2(n_8),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_560),
.A2(n_8),
.B(n_11),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_551),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_562),
.B(n_563),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_564),
.B(n_558),
.C(n_13),
.Y(n_566)
);

NAND3xp33_ASAP7_75t_L g567 ( 
.A(n_566),
.B(n_12),
.C(n_13),
.Y(n_567)
);

NOR3xp33_ASAP7_75t_SL g568 ( 
.A(n_567),
.B(n_565),
.C(n_15),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_12),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_569),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_15),
.Y(n_571)
);


endmodule