module fake_netlist_6_2679_n_643 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_643);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_643;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_625;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_148;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_233;
wire n_617;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_327;
wire n_369;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_542;
wire n_621;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_616;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_164;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_612;
wire n_633;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_151;
wire n_412;
wire n_640;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_7),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_28),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_2),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_48),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_19),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_43),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_83),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_56),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_10),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_42),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_26),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_112),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_93),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_27),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_31),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_80),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_121),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_65),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_21),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_40),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_96),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_2),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_57),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_106),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_95),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_34),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_38),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_72),
.B(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_111),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_68),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_1),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_98),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_116),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_50),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_0),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_109),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_5),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_52),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_102),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_77),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_91),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_54),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_10),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_120),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_13),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_8),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_0),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_145),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_144),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_135),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_145),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_1),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_197),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_3),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_142),
.B(n_4),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_137),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_136),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_157),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_142),
.B(n_6),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_147),
.B(n_9),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_154),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_156),
.B(n_9),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_140),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_176),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_11),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_160),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_165),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_177),
.B(n_15),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_143),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_228),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_231),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_228),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_224),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_211),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_217),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_204),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_204),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_190),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_213),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_213),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_219),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_204),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_230),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_230),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_225),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_219),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_192),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_202),
.A2(n_200),
.B(n_194),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_219),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_233),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_238),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_247),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_238),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_222),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_R g291 ( 
.A(n_221),
.B(n_182),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_248),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_226),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_222),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_246),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_246),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_241),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_243),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_215),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_215),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_288),
.Y(n_306)
);

NOR3xp33_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_239),
.C(n_240),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_215),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_276),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_251),
.B(n_242),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_272),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_215),
.Y(n_315)
);

NOR3xp33_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_239),
.C(n_227),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_287),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_227),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_265),
.A2(n_234),
.B(n_236),
.C(n_207),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_220),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_232),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_232),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_249),
.B(n_207),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_294),
.B(n_184),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_251),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_264),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_229),
.B1(n_223),
.B2(n_203),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_270),
.B(n_220),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_268),
.B(n_148),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_278),
.B(n_149),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_255),
.B(n_250),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_274),
.B(n_281),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_283),
.B(n_220),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_254),
.B(n_243),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_243),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_256),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_296),
.Y(n_345)
);

BUFx6f_ASAP7_75t_SL g346 ( 
.A(n_287),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_284),
.B(n_220),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_273),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_257),
.B(n_244),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g350 ( 
.A(n_267),
.B(n_203),
.C(n_150),
.Y(n_350)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_253),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_280),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_282),
.B(n_244),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_262),
.B(n_244),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_295),
.B(n_245),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_245),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_258),
.B(n_245),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_259),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_279),
.B(n_152),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_279),
.B(n_153),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_L g363 ( 
.A(n_286),
.B(n_145),
.Y(n_363)
);

OR2x6_ASAP7_75t_L g364 ( 
.A(n_251),
.B(n_206),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_287),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_275),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_362),
.B(n_155),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_308),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_325),
.A2(n_180),
.B1(n_163),
.B2(n_164),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_319),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_327),
.A2(n_186),
.B1(n_166),
.B2(n_167),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_309),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_312),
.Y(n_374)
);

CKINVDCx11_ASAP7_75t_R g375 ( 
.A(n_351),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_162),
.Y(n_376)
);

CKINVDCx8_ASAP7_75t_R g377 ( 
.A(n_351),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_344),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_169),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_321),
.B(n_172),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_310),
.Y(n_381)
);

OR2x6_ASAP7_75t_L g382 ( 
.A(n_351),
.B(n_210),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_364),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_301),
.B(n_173),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_303),
.B(n_174),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_313),
.B(n_185),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_357),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_339),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_328),
.B(n_188),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_304),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_355),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_352),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_316),
.A2(n_216),
.B1(n_212),
.B2(n_199),
.Y(n_396)
);

NAND2x1p5_ASAP7_75t_L g397 ( 
.A(n_341),
.B(n_16),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_349),
.B(n_193),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_356),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_317),
.B(n_195),
.Y(n_400)
);

NAND2x1p5_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_17),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_320),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_329),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_302),
.B(n_198),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_318),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_331),
.Y(n_406)
);

NOR3xp33_ASAP7_75t_SL g407 ( 
.A(n_306),
.B(n_23),
.C(n_24),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_304),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_25),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_324),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_350),
.B(n_33),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_363),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_364),
.B(n_39),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_304),
.Y(n_416)
);

O2A1O1Ixp5_ASAP7_75t_L g417 ( 
.A1(n_354),
.A2(n_41),
.B(n_44),
.C(n_45),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_343),
.B(n_342),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_307),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_302),
.B(n_51),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_345),
.Y(n_422)
);

INVx3_ASAP7_75t_SL g423 ( 
.A(n_333),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_305),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_305),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_360),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_302),
.B(n_53),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_R g429 ( 
.A(n_335),
.B(n_55),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_305),
.Y(n_430)
);

AO21x1_ASAP7_75t_L g431 ( 
.A1(n_334),
.A2(n_58),
.B(n_60),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_330),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_376),
.B(n_302),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_389),
.B(n_302),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_315),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_392),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

O2A1O1Ixp33_ASAP7_75t_L g439 ( 
.A1(n_387),
.A2(n_322),
.B(n_311),
.C(n_347),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_420),
.A2(n_330),
.B1(n_346),
.B2(n_359),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_417),
.A2(n_340),
.B(n_332),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_367),
.B(n_61),
.Y(n_442)
);

BUFx12f_ASAP7_75t_L g443 ( 
.A(n_375),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_384),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_396),
.A2(n_346),
.B1(n_63),
.B2(n_64),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_368),
.B(n_62),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_393),
.B(n_67),
.Y(n_448)
);

O2A1O1Ixp33_ASAP7_75t_L g449 ( 
.A1(n_380),
.A2(n_69),
.B(n_71),
.C(n_73),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_75),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_404),
.A2(n_416),
.B(n_426),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_384),
.B(n_79),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_379),
.B(n_82),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_403),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_391),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_419),
.B(n_84),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_391),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_427),
.Y(n_461)
);

O2A1O1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_412),
.A2(n_85),
.B(n_86),
.C(n_89),
.Y(n_462)
);

O2A1O1Ixp33_ASAP7_75t_L g463 ( 
.A1(n_410),
.A2(n_415),
.B(n_406),
.C(n_418),
.Y(n_463)
);

BUFx12f_ASAP7_75t_L g464 ( 
.A(n_368),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_391),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_423),
.B(n_90),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_419),
.B(n_383),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_416),
.A2(n_426),
.B(n_385),
.Y(n_469)
);

BUFx12f_ASAP7_75t_L g470 ( 
.A(n_401),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_372),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_400),
.B(n_92),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_408),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_369),
.B(n_429),
.Y(n_475)
);

CKINVDCx8_ASAP7_75t_R g476 ( 
.A(n_451),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_434),
.A2(n_428),
.B(n_421),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_437),
.Y(n_478)
);

BUFx12f_ASAP7_75t_L g479 ( 
.A(n_443),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_438),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_467),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

AO21x2_ASAP7_75t_L g483 ( 
.A1(n_441),
.A2(n_386),
.B(n_407),
.Y(n_483)
);

BUFx2_ASAP7_75t_SL g484 ( 
.A(n_458),
.Y(n_484)
);

AO21x2_ASAP7_75t_L g485 ( 
.A1(n_441),
.A2(n_431),
.B(n_411),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_436),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_457),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_435),
.B(n_398),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_472),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_465),
.Y(n_490)
);

AO21x2_ASAP7_75t_L g491 ( 
.A1(n_433),
.A2(n_405),
.B(n_424),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_452),
.A2(n_397),
.B(n_425),
.Y(n_492)
);

AOI22x1_ASAP7_75t_L g493 ( 
.A1(n_471),
.A2(n_422),
.B1(n_394),
.B2(n_413),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_448),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_442),
.A2(n_430),
.B(n_395),
.Y(n_495)
);

AOI22x1_ASAP7_75t_L g496 ( 
.A1(n_474),
.A2(n_475),
.B1(n_469),
.B2(n_473),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_456),
.A2(n_395),
.B(n_414),
.Y(n_497)
);

AO21x2_ASAP7_75t_L g498 ( 
.A1(n_459),
.A2(n_371),
.B(n_409),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_432),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_474),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_450),
.A2(n_374),
.B(n_402),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_459),
.A2(n_426),
.B(n_416),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_446),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_447),
.B(n_409),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_SL g506 ( 
.A1(n_503),
.A2(n_440),
.B1(n_445),
.B2(n_466),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_503),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_478),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_480),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_499),
.A2(n_440),
.B1(n_461),
.B2(n_445),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_488),
.A2(n_447),
.B1(n_470),
.B2(n_461),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_468),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_487),
.Y(n_513)
);

BUFx4f_ASAP7_75t_SL g514 ( 
.A(n_479),
.Y(n_514)
);

BUFx8_ASAP7_75t_L g515 ( 
.A(n_479),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_486),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_435),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_489),
.Y(n_518)
);

BUFx12f_ASAP7_75t_L g519 ( 
.A(n_504),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_481),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_494),
.A2(n_504),
.B1(n_453),
.B2(n_496),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_481),
.B(n_468),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_476),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_482),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_502),
.A2(n_463),
.B1(n_465),
.B2(n_460),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_490),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_500),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_500),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_493),
.Y(n_530)
);

NAND2x1_ASAP7_75t_L g531 ( 
.A(n_505),
.B(n_460),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_493),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_527),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_508),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_507),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_518),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_506),
.A2(n_476),
.B1(n_377),
.B2(n_455),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_516),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_512),
.B(n_505),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_517),
.B(n_494),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_516),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_444),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_510),
.B(n_494),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_506),
.B(n_464),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_511),
.A2(n_501),
.B1(n_484),
.B2(n_490),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_523),
.Y(n_546)
);

AND2x4_ASAP7_75t_SL g547 ( 
.A(n_523),
.B(n_458),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_520),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_L g549 ( 
.A(n_522),
.B(n_490),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_L g550 ( 
.A(n_509),
.B(n_490),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_513),
.B(n_498),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_524),
.Y(n_552)
);

OR2x6_ASAP7_75t_L g553 ( 
.A(n_519),
.B(n_484),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_525),
.Y(n_554)
);

OR2x6_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_454),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_529),
.B(n_528),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_R g557 ( 
.A(n_514),
.B(n_490),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_527),
.B(n_498),
.Y(n_558)
);

AO31x2_ASAP7_75t_L g559 ( 
.A1(n_532),
.A2(n_495),
.A3(n_485),
.B(n_491),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_530),
.Y(n_560)
);

AO32x1_ASAP7_75t_L g561 ( 
.A1(n_526),
.A2(n_485),
.A3(n_483),
.B1(n_495),
.B2(n_498),
.Y(n_561)
);

A2O1A1Ixp33_ASAP7_75t_L g562 ( 
.A1(n_521),
.A2(n_462),
.B(n_449),
.C(n_526),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_514),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_551),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_534),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_539),
.B(n_492),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_560),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_540),
.B(n_521),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_546),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_539),
.B(n_483),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_543),
.B(n_483),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_555),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_536),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_548),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_560),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_556),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_542),
.B(n_485),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_548),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_544),
.B(n_491),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_538),
.B(n_491),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_552),
.Y(n_581)
);

AND2x4_ASAP7_75t_SL g582 ( 
.A(n_553),
.B(n_409),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_537),
.A2(n_477),
.B1(n_439),
.B2(n_515),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_554),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_541),
.B(n_492),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_533),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_564),
.B(n_558),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_584),
.Y(n_588)
);

NAND2x1p5_ASAP7_75t_L g589 ( 
.A(n_572),
.B(n_533),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_576),
.B(n_568),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_564),
.B(n_535),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_581),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_562),
.C(n_545),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_568),
.B(n_559),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_565),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_573),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_574),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_580),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_578),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_570),
.B(n_559),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_577),
.B(n_559),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_597),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_597),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_599),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_592),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_599),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_588),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_595),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_598),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_609),
.B(n_605),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_605),
.B(n_587),
.Y(n_611)
);

AOI32xp33_ASAP7_75t_L g612 ( 
.A1(n_602),
.A2(n_583),
.A3(n_591),
.B1(n_590),
.B2(n_594),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_608),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_608),
.B(n_589),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_607),
.B(n_606),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_603),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_611),
.A2(n_593),
.B1(n_579),
.B2(n_572),
.Y(n_617)
);

A2O1A1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_612),
.A2(n_569),
.B(n_572),
.C(n_582),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_616),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_615),
.B(n_604),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_613),
.Y(n_621)
);

NOR2x1_ASAP7_75t_L g622 ( 
.A(n_618),
.B(n_569),
.Y(n_622)
);

AOI322xp5_ASAP7_75t_L g623 ( 
.A1(n_617),
.A2(n_600),
.A3(n_563),
.B1(n_601),
.B2(n_587),
.C1(n_571),
.C2(n_596),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_619),
.B(n_610),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_620),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_621),
.B(n_614),
.Y(n_626)
);

AOI221xp5_ASAP7_75t_L g627 ( 
.A1(n_625),
.A2(n_571),
.B1(n_586),
.B2(n_566),
.C(n_585),
.Y(n_627)
);

NAND3xp33_ASAP7_75t_L g628 ( 
.A(n_623),
.B(n_572),
.C(n_614),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_622),
.A2(n_626),
.B(n_624),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_628),
.A2(n_582),
.B1(n_553),
.B2(n_550),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_629),
.A2(n_549),
.B(n_515),
.Y(n_631)
);

OAI221xp5_ASAP7_75t_SL g632 ( 
.A1(n_630),
.A2(n_631),
.B1(n_627),
.B2(n_555),
.C(n_567),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_632),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_633),
.B(n_575),
.Y(n_634)
);

AOI21xp33_ASAP7_75t_SL g635 ( 
.A1(n_634),
.A2(n_94),
.B(n_99),
.Y(n_635)
);

XNOR2x1_ASAP7_75t_L g636 ( 
.A(n_635),
.B(n_100),
.Y(n_636)
);

OAI31xp33_ASAP7_75t_SL g637 ( 
.A1(n_636),
.A2(n_557),
.A3(n_547),
.B(n_566),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_637),
.A2(n_567),
.B1(n_575),
.B2(n_561),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_638),
.A2(n_497),
.B(n_561),
.Y(n_639)
);

AOI21x1_ASAP7_75t_L g640 ( 
.A1(n_639),
.A2(n_101),
.B(n_103),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_640),
.A2(n_497),
.B1(n_107),
.B2(n_108),
.Y(n_641)
);

OR2x6_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_123),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_642),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_643)
);


endmodule