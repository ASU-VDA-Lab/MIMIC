module fake_jpeg_26911_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_SL g44 ( 
.A1(n_25),
.A2(n_1),
.B(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_33),
.Y(n_67)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_60),
.Y(n_105)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_54),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_26),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_35),
.B1(n_19),
.B2(n_18),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_68),
.B1(n_20),
.B2(n_32),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_35),
.B1(n_29),
.B2(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_31),
.Y(n_86)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_79),
.Y(n_91)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2x1_ASAP7_75t_R g84 ( 
.A(n_66),
.B(n_76),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_94),
.B(n_93),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_98),
.Y(n_117)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_103),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_89),
.B(n_73),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_35),
.B1(n_29),
.B2(n_24),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_63),
.A2(n_22),
.B1(n_30),
.B2(n_28),
.Y(n_98)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_69),
.A2(n_71),
.B1(n_83),
.B2(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_107),
.Y(n_113)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_31),
.B1(n_33),
.B2(n_22),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_106),
.A2(n_80),
.B1(n_81),
.B2(n_54),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_58),
.A2(n_30),
.B1(n_28),
.B2(n_20),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_73),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_58),
.A2(n_32),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_5),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_111)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_112),
.A2(n_121),
.B1(n_103),
.B2(n_110),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_107),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_115),
.Y(n_139)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_120),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_82),
.B(n_72),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_85),
.B(n_96),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_82),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_110),
.B(n_111),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_125),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_62),
.C(n_73),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_131),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

AOI22x1_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_62),
.B1(n_8),
.B2(n_9),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_12),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_144),
.B(n_148),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_129),
.B1(n_131),
.B2(n_130),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_145),
.A2(n_151),
.B1(n_121),
.B2(n_117),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_102),
.B1(n_89),
.B2(n_94),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_155),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_158),
.B(n_160),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_111),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_90),
.B1(n_122),
.B2(n_132),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_121),
.B(n_117),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_161),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_149),
.A2(n_116),
.B1(n_127),
.B2(n_124),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_174),
.B1(n_176),
.B2(n_138),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_120),
.B(n_124),
.Y(n_165)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_173),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_122),
.B1(n_97),
.B2(n_115),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_91),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_169),
.B(n_146),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_156),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_85),
.C(n_132),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_155),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_91),
.B1(n_8),
.B2(n_9),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_150),
.B(n_141),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_180),
.B(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_183),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_138),
.B(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_188),
.A2(n_189),
.B(n_191),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_171),
.B(n_164),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_145),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_190),
.A2(n_191),
.B1(n_188),
.B2(n_181),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_187),
.A2(n_162),
.B1(n_164),
.B2(n_138),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_197),
.B1(n_200),
.B2(n_186),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_173),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_194),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_182),
.B(n_158),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_167),
.B1(n_161),
.B2(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_184),
.B(n_172),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_201),
.B(n_190),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_205),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_184),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_207),
.Y(n_215)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_209),
.B1(n_192),
.B2(n_195),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_189),
.B(n_179),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_179),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_194),
.C(n_197),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_148),
.B(n_159),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_211),
.A2(n_214),
.B1(n_142),
.B2(n_140),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_212),
.B(n_213),
.Y(n_216)
);

NAND2xp33_ASAP7_75t_SL g213 ( 
.A(n_202),
.B(n_168),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_204),
.C(n_202),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_217),
.B(n_218),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_200),
.B1(n_175),
.B2(n_140),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_212),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_216),
.A2(n_210),
.B(n_215),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_222),
.B(n_218),
.Y(n_224)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_224),
.B(n_221),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_225),
.A2(n_144),
.B(n_142),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_12),
.C(n_13),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_11),
.Y(n_228)
);


endmodule