module real_jpeg_18324_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_0),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_0),
.B(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_0),
.A2(n_6),
.B1(n_211),
.B2(n_215),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_0),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_0),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_0),
.B(n_174),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_0),
.B(n_378),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_0),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_0),
.B(n_48),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_1),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_1),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_1),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_1),
.B(n_41),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_1),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_1),
.B(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_1),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_1),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_2),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_2),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_2),
.B(n_31),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_2),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_2),
.B(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_3),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_3),
.Y(n_190)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_3),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_3),
.Y(n_381)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

AND2x4_ASAP7_75t_SL g47 ( 
.A(n_5),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_5),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_5),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_6),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_6),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_6),
.B(n_190),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_6),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_7),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_7),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_7),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_7),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_7),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_7),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_7),
.B(n_437),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_8),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g313 ( 
.A(n_8),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_9),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_9),
.Y(n_175)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_9),
.Y(n_229)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_9),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_10),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_10),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_10),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_10),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_10),
.B(n_107),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_10),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_10),
.B(n_184),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_11),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_73),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_11),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_11),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_11),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_11),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_11),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_12),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_12),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_12),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_12),
.B(n_241),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_12),
.B(n_286),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_12),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_12),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_12),
.B(n_406),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_13),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_13),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_14),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_15),
.Y(n_188)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_199),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_197),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_159),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_21),
.B(n_159),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_96),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_66),
.C(n_88),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_24),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.C(n_51),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_25),
.B(n_39),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_26),
.B(n_30),
.C(n_34),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_28),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_37),
.Y(n_149)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_37),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.C(n_47),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_40),
.B(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_44),
.A2(n_47),
.B1(n_64),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_44),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_45),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_46),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_47),
.Y(n_64)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_53),
.C(n_59),
.Y(n_93)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_50),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_51),
.B(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g218 ( 
.A(n_52),
.B(n_219),
.C(n_221),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_52),
.A2(n_53),
.B1(n_221),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_59),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_59),
.A2(n_65),
.B1(n_104),
.B2(n_105),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_62),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_63),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_105),
.C(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_66),
.B(n_88),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_79),
.C(n_83),
.Y(n_66)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_67),
.B(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.C(n_76),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_68),
.B(n_76),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_70),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_71),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_72),
.B(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_79),
.Y(n_196)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_81),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_90),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_95),
.C(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_87),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_90),
.B(n_183),
.C(n_186),
.Y(n_182)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_93),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_132),
.B1(n_157),
.B2(n_158),
.Y(n_96)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

XNOR2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_113),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_109),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_121),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_121),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.C(n_128),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_128),
.Y(n_156)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_131),
.Y(n_220)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_151),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_135),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_145),
.B1(n_146),
.B2(n_150),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_155),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_160),
.B(n_162),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_164),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_181),
.C(n_194),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_165),
.B(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.C(n_179),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_166),
.B(n_169),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_176),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_170),
.A2(n_176),
.B1(n_177),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_170),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_173),
.B(n_294),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_176),
.B(n_342),
.C(n_345),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_176),
.A2(n_177),
.B1(n_342),
.B2(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_179),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_181),
.B(n_194),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_189),
.C(n_191),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_SL g244 ( 
.A(n_182),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_188),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_189),
.A2(n_191),
.B1(n_192),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_191),
.A2(n_192),
.B1(n_314),
.B2(n_315),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_192),
.B(n_307),
.C(n_314),
.Y(n_306)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AO21x2_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_301),
.B(n_474),
.Y(n_200)
);

NOR2xp67_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_296),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_254),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_203),
.B(n_254),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_247),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_204),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_224),
.C(n_243),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_206),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.C(n_218),
.Y(n_206)
);

XNOR2x2_ASAP7_75t_L g353 ( 
.A(n_207),
.B(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_209),
.A2(n_210),
.B1(n_218),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_210),
.A2(n_321),
.B(n_327),
.Y(n_320)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_214),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_218),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_219),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_224),
.A2(n_243),
.B1(n_244),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_236),
.C(n_240),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.C(n_232),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_226),
.B(n_230),
.C(n_232),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_226),
.B(n_232),
.Y(n_333)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_226),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_230),
.B(n_333),
.Y(n_332)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_235),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_236),
.A2(n_237),
.B1(n_240),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_242),
.Y(n_344)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_247)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_253),
.C(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_250),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.C(n_263),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_260),
.Y(n_362)
);

XOR2x2_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_264),
.B(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_289),
.C(n_293),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_265),
.B(n_357),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_270),
.C(n_280),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g348 ( 
.A(n_267),
.B(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_270),
.B(n_280),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_276),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_271),
.B(n_276),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_278),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.C(n_285),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_281),
.A2(n_284),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_284),
.A2(n_339),
.B1(n_414),
.B2(n_415),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_284),
.B(n_414),
.C(n_420),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_285),
.B(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_289),
.B(n_293),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_296),
.A2(n_475),
.B(n_476),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_297),
.B(n_299),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_470),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_358),
.C(n_363),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_350),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_SL g473 ( 
.A(n_304),
.B(n_350),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_334),
.C(n_348),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_305),
.B(n_468),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_319),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_306),
.B(n_320),
.C(n_332),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_307),
.B(n_459),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_311),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_308),
.B(n_311),
.Y(n_404)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_308),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_308),
.A2(n_423),
.B1(n_424),
.B2(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_313),
.Y(n_331)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_332),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_335),
.B(n_348),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_340),
.C(n_346),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_336),
.B(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_341),
.B(n_347),
.Y(n_454)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_342),
.Y(n_400)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_345),
.B(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_356),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_352),
.B(n_353),
.C(n_356),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_359),
.Y(n_472)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_360),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_465),
.B(n_469),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_450),
.B(n_464),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_408),
.B(n_449),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_395),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_367),
.B(n_395),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_382),
.C(n_389),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_369),
.B(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_373),
.C(n_377),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_377),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_382),
.A2(n_383),
.B1(n_389),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_384),
.B(n_386),
.Y(n_421)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_389),
.Y(n_446)
);

AO22x1_ASAP7_75t_SL g389 ( 
.A1(n_390),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_389)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_390),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_392),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_393),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_394),
.B(n_436),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_401),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_397),
.B(n_401),
.C(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_398),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

MAJx2_ASAP7_75t_L g461 ( 
.A(n_402),
.B(n_404),
.C(n_405),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_443),
.B(n_448),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_410),
.A2(n_425),
.B(n_442),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_422),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_422),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_420),
.B2(n_421),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_424),
.Y(n_434)
);

AOI21x1_ASAP7_75t_SL g425 ( 
.A1(n_426),
.A2(n_435),
.B(n_441),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_433),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_433),
.Y(n_441)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_447),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_444),
.B(n_447),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_462),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_462),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_453),
.B1(n_455),
.B2(n_456),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_457),
.C(n_461),
.Y(n_466)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_458),
.B1(n_460),
.B2(n_461),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_466),
.B(n_467),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_472),
.C(n_473),
.Y(n_470)
);


endmodule