module fake_jpeg_17755_n_231 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_32),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g31 ( 
.A(n_12),
.B(n_15),
.CON(n_31),
.SN(n_31)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_21),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_30),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_30),
.B(n_25),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_44),
.Y(n_50)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_26),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

XNOR2x1_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_55),
.Y(n_64)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_60),
.B1(n_62),
.B2(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_25),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_33),
.A2(n_20),
.B1(n_22),
.B2(n_14),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_20),
.B1(n_22),
.B2(n_14),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_34),
.C(n_42),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_76),
.C(n_79),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_80),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_50),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_40),
.B1(n_27),
.B2(n_32),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_48),
.B1(n_57),
.B2(n_40),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_38),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_28),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_32),
.C(n_28),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_19),
.B(n_13),
.C(n_14),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_64),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_0),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_6),
.B(n_11),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_55),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_12),
.B(n_16),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_27),
.B1(n_57),
.B2(n_48),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_54),
.B1(n_80),
.B2(n_71),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_96),
.Y(n_123)
);

AOI22x1_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_84),
.B1(n_94),
.B2(n_87),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_113),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_79),
.B1(n_65),
.B2(n_72),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_108),
.B1(n_16),
.B2(n_59),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_88),
.B(n_7),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_91),
.B1(n_70),
.B2(n_54),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_67),
.B(n_75),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_109),
.B(n_83),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_85),
.B1(n_94),
.B2(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_63),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_24),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_24),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_118),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_120),
.B(n_109),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_81),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_123),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_126),
.B1(n_100),
.B2(n_101),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_81),
.A3(n_17),
.B1(n_61),
.B2(n_24),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_61),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_133),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_16),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_106),
.B1(n_120),
.B2(n_128),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_138),
.B1(n_150),
.B2(n_59),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_106),
.B1(n_112),
.B2(n_101),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_145),
.B1(n_121),
.B2(n_117),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_104),
.Y(n_146)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_105),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_151),
.B1(n_49),
.B2(n_78),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_99),
.B1(n_113),
.B2(n_103),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_78),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_131),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_165),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_133),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_160),
.C(n_166),
.Y(n_171)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

NAND4xp25_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_141),
.C(n_152),
.D(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_162),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_119),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_121),
.C(n_129),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_11),
.B1(n_10),
.B2(n_8),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_29),
.C(n_35),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_167),
.A2(n_149),
.B1(n_147),
.B2(n_142),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_136),
.C(n_135),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_169),
.C(n_37),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_35),
.C(n_37),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_148),
.B(n_140),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_176),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_155),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_179),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_151),
.B1(n_46),
.B2(n_49),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_35),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_168),
.B(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_169),
.C(n_154),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_182),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_166),
.A2(n_46),
.B1(n_36),
.B2(n_35),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_159),
.C(n_46),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_171),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_174),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_181),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_193),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_36),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_192),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_5),
.B1(n_8),
.B2(n_7),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_5),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_175),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_176),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_0),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_203),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_172),
.B(n_178),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_202),
.B(n_186),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_191),
.A2(n_185),
.B(n_184),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_172),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_211),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_193),
.B(n_194),
.C(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_194),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_4),
.B1(n_7),
.B2(n_6),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_0),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_4),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_212),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_196),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_216),
.A3(n_218),
.B1(n_219),
.B2(n_1),
.C1(n_2),
.C2(n_3),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_1),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_222),
.B(n_223),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_206),
.C(n_23),
.Y(n_222)
);

INVxp33_ASAP7_75t_SL g223 ( 
.A(n_214),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_224),
.C(n_23),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_23),
.C(n_17),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_2),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_229),
.B(n_2),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_3),
.Y(n_231)
);


endmodule