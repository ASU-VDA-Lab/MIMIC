module fake_jpeg_29547_n_287 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_287);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_45),
.B(n_16),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_27),
.B1(n_30),
.B2(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_54),
.A2(n_57),
.B1(n_68),
.B2(n_87),
.Y(n_116)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_37),
.B1(n_34),
.B2(n_27),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_17),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_61),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_47),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_65),
.Y(n_119)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_20),
.B1(n_30),
.B2(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_75),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_35),
.B1(n_22),
.B2(n_32),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_81),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_71),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_38),
.A2(n_34),
.B1(n_23),
.B2(n_20),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_82),
.B1(n_21),
.B2(n_26),
.Y(n_108)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_35),
.Y(n_75)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_18),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_29),
.CON(n_81),
.SN(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_38),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_33),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_31),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_41),
.A2(n_34),
.B1(n_30),
.B2(n_24),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_41),
.B(n_15),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_28),
.B1(n_24),
.B2(n_29),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_97),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_28),
.B(n_29),
.C(n_17),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_103),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_26),
.B1(n_21),
.B2(n_29),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_96),
.B1(n_72),
.B2(n_56),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_26),
.B1(n_21),
.B2(n_17),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_17),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_112),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_65),
.B1(n_61),
.B2(n_73),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_111)
);

AOI32xp33_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_2),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_63),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_114),
.B(n_15),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_121),
.B(n_123),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_120),
.B(n_2),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_74),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_131),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_127),
.A2(n_113),
.B1(n_101),
.B2(n_99),
.Y(n_179)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_129),
.A2(n_133),
.B1(n_152),
.B2(n_137),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_67),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_94),
.A2(n_66),
.B1(n_77),
.B2(n_55),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_134),
.B1(n_136),
.B2(n_145),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_89),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_135),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_94),
.A2(n_111),
.B1(n_116),
.B2(n_90),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_67),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_90),
.A2(n_55),
.B1(n_63),
.B2(n_78),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_78),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_110),
.C(n_92),
.Y(n_171)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_90),
.A2(n_49),
.B1(n_65),
.B2(n_73),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_59),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_147),
.B(n_148),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_104),
.Y(n_148)
);

AO21x2_ASAP7_75t_SL g149 ( 
.A1(n_91),
.A2(n_59),
.B(n_71),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_119),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_49),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_108),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_162),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_SL g157 ( 
.A(n_141),
.B(n_112),
.C(n_95),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_157),
.B(n_164),
.Y(n_185)
);

NOR2x1p5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_124),
.Y(n_158)
);

XOR2x1_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_147),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_SL g164 ( 
.A1(n_121),
.A2(n_120),
.A3(n_92),
.B1(n_109),
.B2(n_102),
.C1(n_105),
.C2(n_110),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_115),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_R g188 ( 
.A(n_167),
.B(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_143),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_177),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_174),
.A2(n_180),
.B(n_149),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_183),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_129),
.B1(n_180),
.B2(n_174),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_117),
.B(n_106),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_196),
.Y(n_217)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_148),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_195),
.Y(n_211)
);

INVxp33_ASAP7_75t_SL g193 ( 
.A(n_181),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_194),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_178),
.B(n_124),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_205),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_207),
.B(n_183),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_122),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_202),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_122),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_197),
.B1(n_202),
.B2(n_192),
.Y(n_222)
);

HAxp5_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_173),
.CON(n_214),
.SN(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_134),
.C(n_150),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_206),
.B(n_161),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_174),
.A2(n_141),
.B(n_149),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_210),
.A2(n_212),
.B(n_218),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_179),
.B(n_159),
.Y(n_212)
);

OA21x2_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_168),
.B(n_165),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_213),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_185),
.Y(n_233)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_171),
.B(n_154),
.Y(n_218)
);

OAI322xp33_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_157),
.A3(n_182),
.B1(n_154),
.B2(n_181),
.C1(n_132),
.C2(n_136),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_110),
.C(n_99),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_205),
.A2(n_175),
.B1(n_170),
.B2(n_163),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_189),
.B1(n_163),
.B2(n_168),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_212),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_200),
.B(n_204),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_166),
.B(n_156),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_226),
.A2(n_188),
.B1(n_187),
.B2(n_194),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_235),
.B1(n_236),
.B2(n_208),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_234),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_218),
.A2(n_196),
.B1(n_184),
.B2(n_206),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_210),
.B1(n_213),
.B2(n_208),
.Y(n_253)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_195),
.C(n_166),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_221),
.C(n_216),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_233),
.B(n_239),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_217),
.B(n_191),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_220),
.A2(n_156),
.B1(n_101),
.B2(n_115),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_213),
.Y(n_255)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_241),
.Y(n_247)
);

FAx1_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_222),
.CI(n_211),
.CON(n_244),
.SN(n_244)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_250),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_220),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_245),
.B(n_248),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_253),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_237),
.B1(n_242),
.B2(n_238),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_255),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_228),
.B1(n_209),
.B2(n_237),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_232),
.C(n_238),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_263),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_240),
.B(n_213),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_254),
.B(n_235),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_216),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_247),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_267),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_257),
.A2(n_255),
.B(n_219),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_266),
.A2(n_271),
.B(n_262),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_250),
.B1(n_241),
.B2(n_225),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_270),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_236),
.Y(n_271)
);

OAI21x1_ASAP7_75t_SL g272 ( 
.A1(n_269),
.A2(n_257),
.B(n_244),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_251),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_260),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_259),
.C(n_225),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_275),
.A2(n_260),
.B(n_251),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_278),
.A2(n_279),
.B(n_276),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_274),
.Y(n_282)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

OAI321xp33_ASAP7_75t_L g284 ( 
.A1(n_282),
.A2(n_283),
.A3(n_4),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_277),
.A2(n_110),
.B(n_6),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_284),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_285),
.Y(n_287)
);


endmodule