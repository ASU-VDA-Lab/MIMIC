module fake_jpeg_2969_n_182 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_182);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_19),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_0),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_70),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_2),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_82),
.Y(n_92)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_58),
.B(n_59),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_82),
.B(n_81),
.C(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_50),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_50),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_52),
.B(n_83),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_76),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_57),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_62),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_53),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_101),
.Y(n_112)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_3),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_22),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_54),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_111),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_98),
.B(n_56),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_54),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_62),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_115),
.C(n_46),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_118),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_4),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_117),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_53),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_4),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_24),
.Y(n_126)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_98),
.B(n_56),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_131),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_56),
.B(n_6),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_5),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_134),
.B(n_138),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_9),
.C(n_10),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_5),
.B(n_6),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_11),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_118),
.B1(n_117),
.B2(n_112),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_141),
.B1(n_9),
.B2(n_11),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_7),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_8),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_139),
.B(n_140),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_28),
.B1(n_42),
.B2(n_41),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_145),
.C(n_157),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_154),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_133),
.C(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_31),
.A3(n_39),
.B1(n_38),
.B2(n_37),
.C1(n_36),
.C2(n_35),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_156),
.B(n_141),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_43),
.B(n_34),
.C(n_33),
.D(n_20),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_12),
.C(n_13),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_145),
.B(n_128),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_161),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_144),
.C(n_123),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_153),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_122),
.B1(n_144),
.B2(n_136),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_156),
.B(n_131),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_165),
.A2(n_14),
.B(n_15),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_170),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_171),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_151),
.C(n_157),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_146),
.A3(n_142),
.B1(n_16),
.B2(n_17),
.C1(n_14),
.C2(n_18),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_162),
.B(n_158),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_165),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_R g176 ( 
.A(n_168),
.B(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_174),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_175),
.C(n_171),
.Y(n_180)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_180),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_15),
.Y(n_182)
);


endmodule