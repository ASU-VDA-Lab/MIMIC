module fake_jpeg_25133_n_400 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_400);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_400;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_45),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_55),
.Y(n_84)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx8_ASAP7_75t_SL g53 ( 
.A(n_30),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_65),
.Y(n_100)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_91),
.Y(n_128)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_76),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_23),
.B1(n_26),
.B2(n_31),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_79),
.A2(n_82),
.B1(n_16),
.B2(n_25),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_23),
.B1(n_26),
.B2(n_31),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_23),
.B1(n_19),
.B2(n_31),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_83),
.A2(n_16),
.B1(n_25),
.B2(n_20),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_86),
.B(n_56),
.Y(n_129)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx2_ASAP7_75t_SL g130 ( 
.A(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_32),
.Y(n_91)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_39),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_55),
.A2(n_18),
.B1(n_26),
.B2(n_21),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_68),
.B(n_36),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_54),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_32),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_30),
.Y(n_133)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_106),
.A2(n_84),
.B(n_75),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_111),
.A2(n_122),
.B(n_148),
.Y(n_162)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_21),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_116),
.Y(n_163)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_72),
.B(n_103),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_125),
.Y(n_170)
);

OR2x2_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_21),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_144),
.B1(n_96),
.B2(n_76),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_20),
.B1(n_22),
.B2(n_29),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_129),
.Y(n_179)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_131),
.B(n_137),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_146),
.B1(n_113),
.B2(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_81),
.B(n_29),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_142),
.Y(n_186)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_29),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_104),
.A2(n_22),
.B1(n_32),
.B2(n_25),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_22),
.B1(n_16),
.B2(n_18),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_102),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_102),
.A2(n_85),
.B1(n_103),
.B2(n_72),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_151),
.B1(n_99),
.B2(n_70),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_47),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_85),
.A2(n_98),
.B1(n_99),
.B2(n_70),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_157),
.A2(n_158),
.B1(n_171),
.B2(n_172),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_121),
.A2(n_98),
.B1(n_92),
.B2(n_90),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_80),
.B(n_73),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_159),
.A2(n_140),
.B(n_77),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_161),
.A2(n_134),
.B(n_110),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_128),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_166),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_80),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_87),
.C(n_78),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_182),
.C(n_145),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_92),
.B1(n_90),
.B2(n_86),
.Y(n_172)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_118),
.A2(n_108),
.B1(n_78),
.B2(n_73),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_185),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_125),
.A2(n_36),
.B1(n_28),
.B2(n_33),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_36),
.B1(n_28),
.B2(n_33),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_41),
.C(n_50),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_132),
.A2(n_33),
.B1(n_28),
.B2(n_27),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_188),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_120),
.Y(n_190)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_187),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_191),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_187),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_192),
.Y(n_260)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_183),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_194),
.B(n_196),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_188),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_116),
.Y(n_197)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_203),
.B(n_213),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_209),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_149),
.B1(n_112),
.B2(n_115),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_211),
.B1(n_225),
.B2(n_185),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_163),
.B(n_122),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_205),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_207),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_122),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_179),
.B(n_141),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_131),
.B1(n_137),
.B2(n_139),
.Y(n_211)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_124),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_179),
.B(n_0),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_217),
.A2(n_227),
.B(n_178),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_218),
.A2(n_219),
.B(n_220),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_168),
.Y(n_220)
);

AO21x2_ASAP7_75t_SL g221 ( 
.A1(n_161),
.A2(n_140),
.B(n_123),
.Y(n_221)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_228),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_164),
.A2(n_152),
.B1(n_171),
.B2(n_170),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_157),
.B(n_77),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_153),
.B(n_152),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_231),
.A2(n_247),
.B1(n_256),
.B2(n_235),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_215),
.C(n_207),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_244),
.C(n_218),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_162),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_233),
.B(n_252),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_172),
.B1(n_162),
.B2(n_184),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_236),
.A2(n_238),
.B1(n_259),
.B2(n_135),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_223),
.B1(n_203),
.B2(n_224),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_167),
.B1(n_182),
.B2(n_184),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_243),
.A2(n_245),
.B1(n_257),
.B2(n_173),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_153),
.C(n_169),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_221),
.A2(n_169),
.B1(n_160),
.B2(n_155),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_155),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_196),
.B(n_46),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_2),
.B(n_3),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_211),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_209),
.B1(n_195),
.B2(n_213),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_195),
.A2(n_160),
.B1(n_173),
.B2(n_140),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_194),
.B(n_174),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_5),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_217),
.A2(n_0),
.B(n_1),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_263),
.A2(n_219),
.B(n_198),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_268),
.C(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_266),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_202),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_276),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_201),
.C(n_220),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_226),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_270),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_208),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_202),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_274),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_204),
.C(n_191),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_214),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_275),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_192),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

OA21x2_ASAP7_75t_L g277 ( 
.A1(n_240),
.A2(n_193),
.B(n_123),
.Y(n_277)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_287),
.B1(n_288),
.B2(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_282),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_135),
.C(n_150),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_268),
.C(n_272),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_1),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_230),
.A2(n_3),
.B(n_4),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_285),
.Y(n_311)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_230),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_240),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_245),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_288)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_238),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_236),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_291),
.A2(n_292),
.B1(n_255),
.B2(n_253),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_283),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_300),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_262),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_305),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_262),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_257),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_279),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_274),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_308),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_309),
.A2(n_293),
.B1(n_311),
.B2(n_302),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_294),
.C(n_296),
.Y(n_318)
);

BUFx24_ASAP7_75t_L g312 ( 
.A(n_277),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_313),
.Y(n_326)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_264),
.B(n_237),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_316),
.Y(n_337)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_277),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_255),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_321),
.C(n_328),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_313),
.A2(n_286),
.B1(n_231),
.B2(n_288),
.Y(n_319)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_281),
.C(n_279),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_324),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_295),
.A2(n_235),
.B1(n_267),
.B2(n_290),
.Y(n_323)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_323),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_246),
.C(n_291),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_304),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_327),
.Y(n_345)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_246),
.C(n_251),
.Y(n_328)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_329),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_303),
.A2(n_263),
.B(n_248),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_330),
.A2(n_297),
.B(n_314),
.Y(n_343)
);

OAI22x1_ASAP7_75t_L g331 ( 
.A1(n_312),
.A2(n_287),
.B1(n_248),
.B2(n_241),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_331),
.A2(n_312),
.B1(n_260),
.B2(n_234),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_334),
.B(n_299),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_251),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_305),
.Y(n_353)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_309),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_299),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_338),
.A2(n_249),
.B1(n_335),
.B2(n_298),
.Y(n_364)
);

BUFx12f_ASAP7_75t_L g339 ( 
.A(n_331),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_319),
.Y(n_356)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_258),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_341),
.B(n_349),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_353),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_321),
.B1(n_330),
.B2(n_324),
.Y(n_362)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_348),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_250),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_306),
.C(n_298),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_350),
.B(n_352),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_364),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_350),
.C(n_342),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_348),
.A2(n_337),
.B(n_293),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_359),
.A2(n_353),
.B(n_322),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_345),
.B(n_328),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_362),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_234),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_363),
.B(n_7),
.Y(n_371)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_365),
.B(n_366),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_320),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_365),
.A2(n_344),
.B1(n_346),
.B2(n_342),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_367),
.B(n_373),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_320),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_357),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_339),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_370),
.B(n_371),
.Y(n_382)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_372),
.B(n_355),
.Y(n_381)
);

XNOR2x1_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_352),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_374),
.A2(n_332),
.B1(n_8),
.B2(n_9),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_375),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_380),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_355),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_381),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_376),
.A2(n_361),
.B(n_364),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_383),
.B(n_372),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_384),
.A2(n_385),
.B1(n_377),
.B2(n_11),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_386),
.B(n_388),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_382),
.B(n_369),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_390),
.A2(n_391),
.B(n_377),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_380),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_387),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_389),
.A2(n_379),
.B(n_384),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_393),
.A2(n_374),
.B(n_378),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_395),
.A2(n_396),
.B1(n_394),
.B2(n_11),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_397),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_398),
.A2(n_10),
.B(n_12),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_399),
.B(n_12),
.Y(n_400)
);


endmodule