module real_aes_18451_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1835;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1802;
wire n_397;
wire n_1083;
wire n_1056;
wire n_1855;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_1772;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1777;
wire n_444;
wire n_1200;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_1851;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_0), .A2(n_266), .B1(n_664), .B2(n_668), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_0), .A2(n_235), .B1(n_467), .B2(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g825 ( .A(n_1), .Y(n_825) );
AND2x2_ASAP7_75t_L g446 ( .A(n_2), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g477 ( .A(n_2), .B(n_242), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_2), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g527 ( .A(n_2), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g1777 ( .A1(n_3), .A2(n_243), .B1(n_617), .B2(n_805), .Y(n_1777) );
AOI22xp33_ASAP7_75t_L g1798 ( .A1(n_3), .A2(n_177), .B1(n_412), .B2(n_681), .Y(n_1798) );
INVx1_ASAP7_75t_L g1479 ( .A(n_4), .Y(n_1479) );
OAI22xp5_ASAP7_75t_L g1491 ( .A1(n_4), .A2(n_81), .B1(n_372), .B2(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_L g655 ( .A(n_5), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_5), .A2(n_136), .B1(n_701), .B2(n_705), .C(n_710), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g1545 ( .A1(n_6), .A2(n_58), .B1(n_1528), .B2(n_1546), .Y(n_1545) );
INVx1_ASAP7_75t_L g1772 ( .A(n_7), .Y(n_1772) );
AOI22xp33_ASAP7_75t_L g1802 ( .A1(n_7), .A2(n_243), .B1(n_681), .B2(n_874), .Y(n_1802) );
INVx1_ASAP7_75t_L g755 ( .A(n_8), .Y(n_755) );
INVx1_ASAP7_75t_L g1171 ( .A(n_9), .Y(n_1171) );
INVx1_ASAP7_75t_L g1468 ( .A(n_10), .Y(n_1468) );
INVx1_ASAP7_75t_L g1044 ( .A(n_11), .Y(n_1044) );
OA222x2_ASAP7_75t_L g1057 ( .A1(n_11), .A2(n_138), .B1(n_161), .B2(n_488), .C1(n_624), .C2(n_1058), .Y(n_1057) );
INVxp67_ASAP7_75t_SL g1158 ( .A(n_12), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_12), .A2(n_115), .B1(n_660), .B2(n_850), .Y(n_1186) );
INVx1_ASAP7_75t_L g1156 ( .A(n_13), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_13), .A2(n_154), .B1(n_403), .B2(n_1188), .Y(n_1187) );
AOI22xp33_ASAP7_75t_SL g1206 ( .A1(n_14), .A2(n_193), .B1(n_412), .B2(n_661), .Y(n_1206) );
AOI221xp5_ASAP7_75t_L g1216 ( .A1(n_14), .A2(n_113), .B1(n_511), .B2(n_819), .C(n_1064), .Y(n_1216) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_15), .A2(n_330), .B1(n_372), .B2(n_377), .C(n_383), .Y(n_371) );
OAI21xp33_ASAP7_75t_SL g487 ( .A1(n_15), .A2(n_488), .B(n_491), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_16), .A2(n_71), .B1(n_551), .B2(n_997), .Y(n_996) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_16), .A2(n_305), .B1(n_934), .B2(n_1016), .C(n_1017), .Y(n_1015) );
INVx2_ASAP7_75t_L g367 ( .A(n_17), .Y(n_367) );
INVx1_ASAP7_75t_L g824 ( .A(n_18), .Y(n_824) );
OAI322xp33_ASAP7_75t_L g828 ( .A1(n_18), .A2(n_829), .A3(n_835), .B1(n_837), .B2(n_844), .C1(n_851), .C2(n_856), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_19), .A2(n_154), .B1(n_467), .B2(n_719), .Y(n_1168) );
AOI22xp5_ASAP7_75t_L g1189 ( .A1(n_19), .A2(n_304), .B1(n_1188), .B2(n_1190), .Y(n_1189) );
CKINVDCx5p33_ASAP7_75t_R g1296 ( .A(n_20), .Y(n_1296) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_21), .A2(n_164), .B1(n_1034), .B2(n_1037), .Y(n_1036) );
INVxp67_ASAP7_75t_SL g1076 ( .A(n_21), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g815 ( .A1(n_22), .A2(n_223), .B1(n_689), .B2(n_816), .C(n_818), .Y(n_815) );
INVx1_ASAP7_75t_L g842 ( .A(n_22), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_23), .A2(n_278), .B1(n_417), .B2(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g481 ( .A(n_23), .Y(n_481) );
INVx1_ASAP7_75t_L g930 ( .A(n_24), .Y(n_930) );
CKINVDCx5p33_ASAP7_75t_R g984 ( .A(n_25), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_26), .A2(n_309), .B1(n_417), .B2(n_420), .Y(n_756) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_26), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g1555 ( .A1(n_27), .A2(n_202), .B1(n_1535), .B2(n_1538), .Y(n_1555) );
INVx1_ASAP7_75t_L g1246 ( .A(n_28), .Y(n_1246) );
AOI221xp5_ASAP7_75t_L g1261 ( .A1(n_28), .A2(n_133), .B1(n_551), .B2(n_1262), .C(n_1264), .Y(n_1261) );
INVx1_ASAP7_75t_L g595 ( .A(n_29), .Y(n_595) );
AOI221x1_ASAP7_75t_SL g601 ( .A1(n_29), .A2(n_183), .B1(n_467), .B2(n_602), .C(n_606), .Y(n_601) );
OA22x2_ASAP7_75t_L g1361 ( .A1(n_30), .A2(n_1362), .B1(n_1460), .B2(n_1461), .Y(n_1361) );
INVxp67_ASAP7_75t_L g1461 ( .A(n_30), .Y(n_1461) );
AOI22xp5_ASAP7_75t_L g1544 ( .A1(n_30), .A2(n_174), .B1(n_1535), .B2(n_1538), .Y(n_1544) );
HB1xp67_ASAP7_75t_L g1515 ( .A(n_31), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1529 ( .A(n_31), .B(n_1513), .Y(n_1529) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_32), .A2(n_214), .B1(n_1041), .B2(n_1108), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_32), .A2(n_291), .B1(n_939), .B2(n_1139), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_33), .A2(n_290), .B1(n_617), .B2(n_821), .Y(n_820) );
INVxp67_ASAP7_75t_L g833 ( .A(n_33), .Y(n_833) );
INVx1_ASAP7_75t_L g586 ( .A(n_34), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_34), .A2(n_165), .B1(n_512), .B2(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g1401 ( .A(n_35), .Y(n_1401) );
INVx1_ASAP7_75t_L g790 ( .A(n_36), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g1580 ( .A1(n_36), .A2(n_268), .B1(n_1535), .B2(n_1538), .Y(n_1580) );
OAI211xp5_ASAP7_75t_SL g926 ( .A1(n_37), .A2(n_927), .B(n_929), .C(n_932), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_37), .A2(n_265), .B1(n_645), .B2(n_859), .Y(n_975) );
INVx1_ASAP7_75t_L g744 ( .A(n_38), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_39), .A2(n_288), .B1(n_617), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_39), .A2(n_223), .B1(n_660), .B2(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g1253 ( .A(n_40), .Y(n_1253) );
OAI22xp33_ASAP7_75t_L g1259 ( .A1(n_40), .A2(n_53), .B1(n_372), .B2(n_377), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_41), .A2(n_235), .B1(n_664), .B2(n_668), .Y(n_1204) );
AOI221xp5_ASAP7_75t_L g1213 ( .A1(n_41), .A2(n_266), .B1(n_533), .B2(n_535), .C(n_715), .Y(n_1213) );
AOI22xp5_ASAP7_75t_L g1551 ( .A1(n_42), .A2(n_112), .B1(n_1535), .B2(n_1538), .Y(n_1551) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_43), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_44), .A2(n_263), .B1(n_1033), .B2(n_1034), .Y(n_1032) );
INVxp67_ASAP7_75t_SL g1066 ( .A(n_44), .Y(n_1066) );
INVxp67_ASAP7_75t_SL g1161 ( .A(n_45), .Y(n_1161) );
AOI22xp33_ASAP7_75t_SL g1191 ( .A1(n_45), .A2(n_92), .B1(n_660), .B2(n_850), .Y(n_1191) );
INVx1_ASAP7_75t_L g885 ( .A(n_46), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g1549 ( .A1(n_47), .A2(n_158), .B1(n_1528), .B2(n_1550), .Y(n_1549) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_48), .A2(n_396), .B1(n_1284), .B2(n_1287), .Y(n_1283) );
INVx1_ASAP7_75t_L g1301 ( .A(n_48), .Y(n_1301) );
CKINVDCx5p33_ASAP7_75t_R g1198 ( .A(n_49), .Y(n_1198) );
INVx1_ASAP7_75t_L g882 ( .A(n_50), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_50), .A2(n_256), .B1(n_535), .B2(n_911), .C(n_912), .Y(n_910) );
OAI221xp5_ASAP7_75t_L g940 ( .A1(n_51), .A2(n_114), .B1(n_706), .B2(n_941), .C(n_942), .Y(n_940) );
OAI22xp33_ASAP7_75t_L g968 ( .A1(n_51), .A2(n_114), .B1(n_969), .B2(n_971), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1832 ( .A1(n_52), .A2(n_176), .B1(n_467), .B2(n_720), .Y(n_1832) );
INVx1_ASAP7_75t_L g1857 ( .A(n_52), .Y(n_1857) );
OAI221xp5_ASAP7_75t_L g1249 ( .A1(n_53), .A2(n_299), .B1(n_491), .B2(n_620), .C(n_622), .Y(n_1249) );
INVx1_ASAP7_75t_L g730 ( .A(n_54), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g947 ( .A1(n_55), .A2(n_246), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_55), .A2(n_333), .B1(n_660), .B2(n_681), .Y(n_959) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_56), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g1769 ( .A(n_57), .Y(n_1769) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_59), .A2(n_660), .B(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_59), .Y(n_768) );
INVx1_ASAP7_75t_L g1208 ( .A(n_60), .Y(n_1208) );
CKINVDCx5p33_ASAP7_75t_R g1241 ( .A(n_61), .Y(n_1241) );
INVx1_ASAP7_75t_L g1290 ( .A(n_62), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_62), .A2(n_65), .B1(n_686), .B2(n_720), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1834 ( .A1(n_63), .A2(n_204), .B1(n_719), .B2(n_1131), .Y(n_1834) );
INVx1_ASAP7_75t_L g1852 ( .A(n_63), .Y(n_1852) );
AOI22xp33_ASAP7_75t_L g1659 ( .A1(n_64), .A2(n_228), .B1(n_1528), .B2(n_1546), .Y(n_1659) );
AOI221xp5_ASAP7_75t_L g1278 ( .A1(n_65), .A2(n_325), .B1(n_751), .B2(n_1188), .C(n_1279), .Y(n_1278) );
OAI222xp33_ASAP7_75t_L g1317 ( .A1(n_66), .A2(n_82), .B1(n_1318), .B2(n_1319), .C1(n_1325), .C2(n_1331), .Y(n_1317) );
INVx1_ASAP7_75t_L g1345 ( .A(n_66), .Y(n_1345) );
INVxp67_ASAP7_75t_SL g1251 ( .A(n_67), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_67), .A2(n_396), .B1(n_1267), .B2(n_1268), .Y(n_1266) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_68), .A2(n_244), .B1(n_372), .B2(n_377), .C(n_383), .Y(n_731) );
OAI221xp5_ASAP7_75t_L g781 ( .A1(n_68), .A2(n_309), .B1(n_491), .B2(n_620), .C(n_622), .Y(n_781) );
OAI222xp33_ASAP7_75t_L g1756 ( .A1(n_69), .A2(n_166), .B1(n_538), .B2(n_1441), .C1(n_1757), .C2(n_1759), .Y(n_1756) );
OAI222xp33_ASAP7_75t_L g1781 ( .A1(n_69), .A2(n_166), .B1(n_210), .B2(n_1782), .C1(n_1783), .C2(n_1785), .Y(n_1781) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_70), .A2(n_275), .B1(n_389), .B2(n_396), .Y(n_886) );
INVxp67_ASAP7_75t_SL g891 ( .A(n_70), .Y(n_891) );
AOI22xp33_ASAP7_75t_SL g1013 ( .A1(n_71), .A2(n_137), .B1(n_805), .B2(n_938), .Y(n_1013) );
AOI21xp33_ASAP7_75t_L g423 ( .A1(n_72), .A2(n_424), .B(n_427), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_72), .A2(n_105), .B1(n_532), .B2(n_534), .C(n_536), .Y(n_531) );
INVx1_ASAP7_75t_L g1087 ( .A(n_73), .Y(n_1087) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_74), .Y(n_860) );
INVx1_ASAP7_75t_L g811 ( .A(n_75), .Y(n_811) );
OAI211xp5_ASAP7_75t_L g861 ( .A1(n_75), .A2(n_862), .B(n_863), .C(n_866), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g1096 ( .A(n_76), .Y(n_1096) );
INVx1_ASAP7_75t_L g1255 ( .A(n_77), .Y(n_1255) );
OAI222xp33_ASAP7_75t_L g1258 ( .A1(n_77), .A2(n_284), .B1(n_299), .B2(n_393), .C1(n_580), .C2(n_843), .Y(n_1258) );
AOI21xp33_ASAP7_75t_L g945 ( .A1(n_78), .A2(n_497), .B(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g955 ( .A(n_78), .Y(n_955) );
XOR2x2_ASAP7_75t_L g353 ( .A(n_79), .B(n_354), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g1564 ( .A1(n_80), .A2(n_159), .B1(n_1528), .B2(n_1535), .Y(n_1564) );
INVx1_ASAP7_75t_L g1473 ( .A(n_81), .Y(n_1473) );
INVx1_ASAP7_75t_L g1347 ( .A(n_82), .Y(n_1347) );
OAI22xp33_ASAP7_75t_L g1392 ( .A1(n_83), .A2(n_172), .B1(n_1393), .B2(n_1395), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g1443 ( .A1(n_83), .A2(n_172), .B1(n_1444), .B2(n_1448), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g1563 ( .A1(n_84), .A2(n_294), .B1(n_1538), .B2(n_1546), .Y(n_1563) );
OAI221xp5_ASAP7_75t_L g1816 ( .A1(n_85), .A2(n_119), .B1(n_1067), .B2(n_1817), .C(n_1818), .Y(n_1816) );
INVx1_ASAP7_75t_L g1839 ( .A(n_85), .Y(n_1839) );
AOI22xp5_ASAP7_75t_L g1527 ( .A1(n_86), .A2(n_146), .B1(n_1528), .B2(n_1532), .Y(n_1527) );
XNOR2xp5_ASAP7_75t_L g1810 ( .A(n_87), .B(n_1811), .Y(n_1810) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_88), .A2(n_338), .B1(n_660), .B2(n_661), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_88), .A2(n_187), .B1(n_602), .B2(n_689), .C(n_690), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g1178 ( .A(n_89), .Y(n_1178) );
XOR2xp5_ASAP7_75t_L g1194 ( .A(n_90), .B(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1415 ( .A(n_91), .Y(n_1415) );
AOI221xp5_ASAP7_75t_L g1167 ( .A1(n_92), .A2(n_115), .B1(n_497), .B2(n_901), .C(n_936), .Y(n_1167) );
INVx1_ASAP7_75t_L g1820 ( .A(n_93), .Y(n_1820) );
OAI221xp5_ASAP7_75t_SL g1844 ( .A1(n_93), .A2(n_116), .B1(n_375), .B2(n_565), .C(n_876), .Y(n_1844) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_94), .A2(n_198), .B1(n_389), .B2(n_396), .Y(n_388) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_94), .Y(n_519) );
INVx1_ASAP7_75t_L g1221 ( .A(n_95), .Y(n_1221) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_96), .A2(n_111), .B1(n_736), .B2(n_1040), .C(n_1041), .Y(n_1039) );
AOI22xp33_ASAP7_75t_SL g1077 ( .A1(n_96), .A2(n_263), .B1(n_720), .B2(n_939), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1660 ( .A1(n_97), .A2(n_316), .B1(n_1535), .B2(n_1538), .Y(n_1660) );
AOI222xp33_ASAP7_75t_L g428 ( .A1(n_98), .A2(n_142), .B1(n_322), .B2(n_398), .C1(n_429), .C2(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g539 ( .A(n_98), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g1242 ( .A(n_99), .Y(n_1242) );
INVx1_ASAP7_75t_L g878 ( .A(n_100), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_100), .A2(n_181), .B1(n_901), .B2(n_903), .C(n_905), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g1297 ( .A1(n_101), .A2(n_139), .B1(n_372), .B2(n_377), .Y(n_1297) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_101), .A2(n_282), .B1(n_620), .B2(n_622), .Y(n_1311) );
INVxp67_ASAP7_75t_SL g1326 ( .A(n_102), .Y(n_1326) );
AOI22xp33_ASAP7_75t_SL g1352 ( .A1(n_102), .A2(n_270), .B1(n_660), .B2(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1416 ( .A(n_103), .Y(n_1416) );
CKINVDCx5p33_ASAP7_75t_R g1247 ( .A(n_104), .Y(n_1247) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_105), .A2(n_213), .B1(n_401), .B2(n_404), .C(n_408), .Y(n_400) );
INVx1_ASAP7_75t_L g1513 ( .A(n_106), .Y(n_1513) );
INVx1_ASAP7_75t_L g1286 ( .A(n_107), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_107), .A2(n_325), .B1(n_467), .B2(n_720), .Y(n_1306) );
INVx1_ASAP7_75t_L g1252 ( .A(n_108), .Y(n_1252) );
INVx1_ASAP7_75t_L g370 ( .A(n_109), .Y(n_370) );
OAI21xp33_ASAP7_75t_L g461 ( .A1(n_109), .A2(n_462), .B(n_471), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g1833 ( .A1(n_110), .A2(n_144), .B1(n_602), .B2(n_689), .C(n_936), .Y(n_1833) );
INVx1_ASAP7_75t_L g1848 ( .A(n_110), .Y(n_1848) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_111), .A2(n_149), .B1(n_689), .B2(n_1064), .C(n_1065), .Y(n_1063) );
XOR2xp5_ASAP7_75t_L g1749 ( .A(n_112), .B(n_1750), .Y(n_1749) );
AOI22xp5_ASAP7_75t_L g1808 ( .A1(n_112), .A2(n_1809), .B1(n_1860), .B2(n_1864), .Y(n_1808) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_113), .A2(n_240), .B1(n_1202), .B2(n_1203), .Y(n_1201) );
INVx1_ASAP7_75t_L g1827 ( .A(n_116), .Y(n_1827) );
INVx1_ASAP7_75t_L g555 ( .A(n_117), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_117), .A2(n_238), .B1(n_620), .B2(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g1338 ( .A(n_118), .Y(n_1338) );
INVx1_ASAP7_75t_L g1837 ( .A(n_119), .Y(n_1837) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_120), .A2(n_227), .B1(n_938), .B2(n_939), .Y(n_937) );
INVx1_ASAP7_75t_L g958 ( .A(n_120), .Y(n_958) );
XOR2x2_ASAP7_75t_L g634 ( .A(n_121), .B(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g1083 ( .A1(n_122), .A2(n_1084), .B1(n_1085), .B2(n_1146), .Y(n_1083) );
INVx1_ASAP7_75t_L g1146 ( .A(n_122), .Y(n_1146) );
INVx1_ASAP7_75t_L g1824 ( .A(n_123), .Y(n_1824) );
OAI21xp33_ASAP7_75t_L g1842 ( .A1(n_123), .A2(n_639), .B(n_1843), .Y(n_1842) );
CKINVDCx5p33_ASAP7_75t_R g985 ( .A(n_124), .Y(n_985) );
AOI22xp33_ASAP7_75t_SL g1579 ( .A1(n_125), .A2(n_190), .B1(n_1528), .B2(n_1546), .Y(n_1579) );
CKINVDCx5p33_ASAP7_75t_R g1281 ( .A(n_126), .Y(n_1281) );
AOI22xp33_ASAP7_75t_SL g1477 ( .A1(n_127), .A2(n_247), .B1(n_719), .B2(n_939), .Y(n_1477) );
AOI221xp5_ASAP7_75t_L g1497 ( .A1(n_127), .A2(n_321), .B1(n_660), .B2(n_736), .C(n_1040), .Y(n_1497) );
INVx1_ASAP7_75t_L g808 ( .A(n_128), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_129), .Y(n_643) );
OAI211xp5_ASAP7_75t_SL g1164 ( .A1(n_130), .A2(n_1165), .B(n_1166), .C(n_1169), .Y(n_1164) );
INVx1_ASAP7_75t_L g1184 ( .A(n_130), .Y(n_1184) );
AOI22xp33_ASAP7_75t_SL g992 ( .A1(n_131), .A2(n_295), .B1(n_993), .B2(n_995), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_131), .A2(n_280), .B1(n_805), .B2(n_938), .Y(n_1018) );
OAI222xp33_ASAP7_75t_L g1153 ( .A1(n_132), .A2(n_258), .B1(n_706), .B2(n_941), .C1(n_1154), .C2(n_1157), .Y(n_1153) );
INVx1_ASAP7_75t_L g1181 ( .A(n_132), .Y(n_1181) );
INVx1_ASAP7_75t_L g1232 ( .A(n_133), .Y(n_1232) );
INVx1_ASAP7_75t_L g1323 ( .A(n_134), .Y(n_1323) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_134), .A2(n_192), .B1(n_664), .B2(n_999), .Y(n_1354) );
XNOR2x1_ASAP7_75t_L g1149 ( .A(n_135), .B(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g652 ( .A(n_136), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_137), .A2(n_305), .B1(n_431), .B2(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1054 ( .A(n_138), .Y(n_1054) );
INVx1_ASAP7_75t_L g1302 ( .A(n_139), .Y(n_1302) );
AOI221xp5_ASAP7_75t_SL g1831 ( .A1(n_140), .A2(n_302), .B1(n_602), .B2(n_689), .C(n_715), .Y(n_1831) );
INVx1_ASAP7_75t_L g1854 ( .A(n_140), .Y(n_1854) );
CKINVDCx5p33_ASAP7_75t_R g1829 ( .A(n_141), .Y(n_1829) );
INVx1_ASAP7_75t_L g504 ( .A(n_142), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_143), .A2(n_197), .B1(n_511), .B2(n_799), .C(n_802), .Y(n_798) );
INVxp67_ASAP7_75t_L g830 ( .A(n_143), .Y(n_830) );
INVx1_ASAP7_75t_L g1858 ( .A(n_144), .Y(n_1858) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_145), .A2(n_298), .B1(n_664), .B2(n_666), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_145), .A2(n_253), .B1(n_692), .B2(n_693), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g933 ( .A1(n_147), .A2(n_333), .B1(n_934), .B2(n_935), .C(n_936), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_147), .A2(n_246), .B1(n_660), .B2(n_965), .Y(n_964) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_148), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g1035 ( .A1(n_149), .A2(n_171), .B1(n_748), .B2(n_850), .C(n_997), .Y(n_1035) );
AOI221xp5_ASAP7_75t_L g879 ( .A1(n_150), .A2(n_181), .B1(n_551), .B2(n_880), .C(n_881), .Y(n_879) );
INVx1_ASAP7_75t_L g916 ( .A(n_150), .Y(n_916) );
INVxp67_ASAP7_75t_SL g1091 ( .A(n_151), .Y(n_1091) );
OAI221xp5_ASAP7_75t_L g1109 ( .A1(n_151), .A2(n_383), .B1(n_389), .B2(n_1110), .C(n_1115), .Y(n_1109) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_152), .A2(n_748), .B(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1128 ( .A(n_152), .Y(n_1128) );
INVx1_ASAP7_75t_L g1114 ( .A(n_153), .Y(n_1114) );
AOI22xp33_ASAP7_75t_SL g1130 ( .A1(n_153), .A2(n_214), .B1(n_692), .B2(n_1131), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_155), .A2(n_335), .B1(n_398), .B2(n_751), .Y(n_750) );
INVxp67_ASAP7_75t_SL g778 ( .A(n_155), .Y(n_778) );
INVx1_ASAP7_75t_L g1197 ( .A(n_156), .Y(n_1197) );
INVx1_ASAP7_75t_L g1292 ( .A(n_157), .Y(n_1292) );
INVx1_ASAP7_75t_L g734 ( .A(n_160), .Y(n_734) );
OAI221xp5_ASAP7_75t_L g1049 ( .A1(n_161), .A2(n_163), .B1(n_587), .B2(n_1050), .C(n_1051), .Y(n_1049) );
INVx1_ASAP7_75t_L g1170 ( .A(n_162), .Y(n_1170) );
INVxp67_ASAP7_75t_SL g1060 ( .A(n_163), .Y(n_1060) );
INVxp33_ASAP7_75t_SL g1068 ( .A(n_164), .Y(n_1068) );
INVx1_ASAP7_75t_L g578 ( .A(n_165), .Y(n_578) );
INVx2_ASAP7_75t_L g1531 ( .A(n_167), .Y(n_1531) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_167), .B(n_292), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_167), .B(n_1537), .Y(n_1539) );
INVxp67_ASAP7_75t_SL g1330 ( .A(n_168), .Y(n_1330) );
AOI22xp33_ASAP7_75t_SL g1357 ( .A1(n_168), .A2(n_307), .B1(n_562), .B2(n_995), .Y(n_1357) );
XNOR2xp5_ASAP7_75t_L g923 ( .A(n_169), .B(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g1209 ( .A(n_170), .Y(n_1209) );
INVx1_ASAP7_75t_L g1074 ( .A(n_171), .Y(n_1074) );
AOI22xp5_ASAP7_75t_L g1557 ( .A1(n_173), .A2(n_234), .B1(n_1528), .B2(n_1538), .Y(n_1557) );
OAI21xp33_ASAP7_75t_L g1470 ( .A1(n_175), .A2(n_624), .B(n_1471), .Y(n_1470) );
OAI221xp5_ASAP7_75t_L g1500 ( .A1(n_175), .A2(n_274), .B1(n_961), .B2(n_1501), .C(n_1502), .Y(n_1500) );
INVx1_ASAP7_75t_L g1847 ( .A(n_176), .Y(n_1847) );
INVx1_ASAP7_75t_L g1773 ( .A(n_177), .Y(n_1773) );
INVx1_ASAP7_75t_L g742 ( .A(n_178), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g1558 ( .A1(n_179), .A2(n_184), .B1(n_1532), .B2(n_1535), .Y(n_1558) );
OAI221xp5_ASAP7_75t_L g887 ( .A1(n_180), .A2(n_267), .B1(n_372), .B2(n_377), .C(n_383), .Y(n_887) );
INVx1_ASAP7_75t_L g921 ( .A(n_180), .Y(n_921) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_182), .Y(n_570) );
INVx1_ASAP7_75t_L g581 ( .A(n_183), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g989 ( .A(n_185), .Y(n_989) );
INVx1_ASAP7_75t_L g1053 ( .A(n_186), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_186), .A2(n_225), .B1(n_474), .B2(n_483), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_187), .A2(n_199), .B1(n_660), .B2(n_661), .Y(n_659) );
OAI211xp5_ASAP7_75t_L g1752 ( .A1(n_188), .A2(n_1753), .B(n_1754), .C(n_1763), .Y(n_1752) );
INVx1_ASAP7_75t_L g1790 ( .A(n_188), .Y(n_1790) );
CKINVDCx5p33_ASAP7_75t_R g1117 ( .A(n_189), .Y(n_1117) );
AOI22xp33_ASAP7_75t_SL g1476 ( .A1(n_191), .A2(n_310), .B1(n_604), .B2(n_911), .Y(n_1476) );
AOI221xp5_ASAP7_75t_L g1496 ( .A1(n_191), .A2(n_221), .B1(n_664), .B2(n_748), .C(n_1040), .Y(n_1496) );
AOI22xp33_ASAP7_75t_L g1335 ( .A1(n_192), .A2(n_339), .B1(n_617), .B2(n_804), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_193), .A2(n_240), .B1(n_719), .B2(n_939), .Y(n_1214) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_194), .A2(n_280), .B1(n_978), .B2(n_995), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_194), .A2(n_295), .B1(n_534), .B2(n_819), .C(n_1009), .Y(n_1008) );
INVx2_ASAP7_75t_L g369 ( .A(n_195), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_195), .B(n_367), .Y(n_392) );
INVx1_ASAP7_75t_L g434 ( .A(n_195), .Y(n_434) );
INVx1_ASAP7_75t_L g974 ( .A(n_196), .Y(n_974) );
INVxp67_ASAP7_75t_L g847 ( .A(n_197), .Y(n_847) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_198), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_199), .A2(n_338), .B1(n_693), .B2(n_719), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g1534 ( .A1(n_200), .A2(n_327), .B1(n_1535), .B2(n_1538), .Y(n_1534) );
XOR2xp5_ASAP7_75t_L g543 ( .A(n_201), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g1226 ( .A(n_202), .Y(n_1226) );
OAI22xp33_ASAP7_75t_L g556 ( .A1(n_203), .A2(n_301), .B1(n_557), .B2(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g629 ( .A(n_203), .Y(n_629) );
INVx1_ASAP7_75t_L g1855 ( .A(n_204), .Y(n_1855) );
INVx1_ASAP7_75t_L g1407 ( .A(n_205), .Y(n_1407) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_206), .Y(n_1005) );
INVx1_ASAP7_75t_L g1762 ( .A(n_207), .Y(n_1762) );
OAI22xp5_ASAP7_75t_L g1787 ( .A1(n_207), .A2(n_241), .B1(n_1394), .B2(n_1397), .Y(n_1787) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_208), .A2(n_320), .B1(n_719), .B2(n_1483), .Y(n_1482) );
AOI22xp33_ASAP7_75t_L g1495 ( .A1(n_208), .A2(n_247), .B1(n_660), .B2(n_1188), .Y(n_1495) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_209), .A2(n_297), .B1(n_645), .B2(n_647), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g683 ( .A1(n_209), .A2(n_684), .B(n_687), .C(n_695), .Y(n_683) );
INVx1_ASAP7_75t_L g1755 ( .A(n_210), .Y(n_1755) );
INVx1_ASAP7_75t_L g1322 ( .A(n_211), .Y(n_1322) );
AOI22xp33_ASAP7_75t_SL g1355 ( .A1(n_211), .A2(n_339), .B1(n_999), .B2(n_1356), .Y(n_1355) );
BUFx3_ASAP7_75t_L g361 ( .A(n_212), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_213), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g410 ( .A(n_215), .Y(n_410) );
OAI21xp5_ASAP7_75t_SL g1022 ( .A1(n_216), .A2(n_794), .B(n_1023), .Y(n_1022) );
OAI221xp5_ASAP7_75t_L g1293 ( .A1(n_217), .A2(n_282), .B1(n_1103), .B2(n_1294), .C(n_1295), .Y(n_1293) );
OAI211xp5_ASAP7_75t_L g1299 ( .A1(n_217), .A2(n_893), .B(n_1300), .C(n_1303), .Y(n_1299) );
INVx1_ASAP7_75t_L g1472 ( .A(n_218), .Y(n_1472) );
OAI21xp5_ASAP7_75t_SL g1339 ( .A1(n_219), .A2(n_794), .B(n_1340), .Y(n_1339) );
CKINVDCx5p33_ASAP7_75t_R g1280 ( .A(n_220), .Y(n_1280) );
AOI22xp33_ASAP7_75t_L g1485 ( .A1(n_221), .A2(n_321), .B1(n_1016), .B2(n_1486), .Y(n_1485) );
OAI21xp5_ASAP7_75t_L g1172 ( .A1(n_222), .A2(n_645), .B(n_1173), .Y(n_1172) );
OAI22xp33_ASAP7_75t_L g672 ( .A1(n_224), .A2(n_331), .B1(n_673), .B2(n_677), .Y(n_672) );
INVx1_ASAP7_75t_L g696 ( .A(n_224), .Y(n_696) );
INVx1_ASAP7_75t_L g1043 ( .A(n_225), .Y(n_1043) );
OAI211xp5_ASAP7_75t_SL g1377 ( .A1(n_226), .A2(n_1378), .B(n_1380), .C(n_1382), .Y(n_1377) );
INVx1_ASAP7_75t_L g1439 ( .A(n_226), .Y(n_1439) );
INVx1_ASAP7_75t_L g963 ( .A(n_227), .Y(n_963) );
INVx1_ASAP7_75t_L g1768 ( .A(n_229), .Y(n_1768) );
NAND2xp5_ASAP7_75t_L g1799 ( .A(n_229), .B(n_1034), .Y(n_1799) );
INVx1_ASAP7_75t_L g754 ( .A(n_230), .Y(n_754) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_231), .Y(n_1090) );
INVx1_ASAP7_75t_L g1391 ( .A(n_232), .Y(n_1391) );
OAI211xp5_ASAP7_75t_SL g1430 ( .A1(n_232), .A2(n_1431), .B(n_1432), .C(n_1435), .Y(n_1430) );
CKINVDCx5p33_ASAP7_75t_R g1237 ( .A(n_233), .Y(n_1237) );
INVx1_ASAP7_75t_L g1337 ( .A(n_236), .Y(n_1337) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_237), .A2(n_253), .B1(n_664), .B2(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g711 ( .A(n_237), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g564 ( .A1(n_238), .A2(n_257), .B1(n_375), .B2(n_565), .C(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g931 ( .A(n_239), .Y(n_931) );
INVx1_ASAP7_75t_L g1765 ( .A(n_241), .Y(n_1765) );
INVx1_ASAP7_75t_L g447 ( .A(n_242), .Y(n_447) );
BUFx3_ASAP7_75t_L g518 ( .A(n_242), .Y(n_518) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_244), .Y(n_785) );
OAI211xp5_ASAP7_75t_L g1332 ( .A1(n_245), .A2(n_1165), .B(n_1333), .C(n_1336), .Y(n_1332) );
INVx1_ASAP7_75t_L g1349 ( .A(n_245), .Y(n_1349) );
NOR2xp33_ASAP7_75t_L g1142 ( .A(n_248), .B(n_1143), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_249), .Y(n_591) );
INVxp67_ASAP7_75t_SL g1464 ( .A(n_250), .Y(n_1464) );
CKINVDCx5p33_ASAP7_75t_R g1819 ( .A(n_251), .Y(n_1819) );
INVx1_ASAP7_75t_L g1098 ( .A(n_252), .Y(n_1098) );
CKINVDCx5p33_ASAP7_75t_R g1288 ( .A(n_254), .Y(n_1288) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_255), .A2(n_319), .B1(n_551), .B2(n_874), .C(n_875), .Y(n_873) );
INVx1_ASAP7_75t_L g906 ( .A(n_255), .Y(n_906) );
INVx1_ASAP7_75t_L g877 ( .A(n_256), .Y(n_877) );
OA222x2_ASAP7_75t_L g623 ( .A1(n_257), .A2(n_271), .B1(n_323), .B2(n_462), .C1(n_488), .C2(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g1182 ( .A(n_258), .Y(n_1182) );
XOR2xp5_ASAP7_75t_L g868 ( .A(n_259), .B(n_869), .Y(n_868) );
OAI21xp5_ASAP7_75t_L g1222 ( .A1(n_260), .A2(n_794), .B(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g413 ( .A(n_261), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g1113 ( .A(n_262), .Y(n_1113) );
XOR2x2_ASAP7_75t_L g1314 ( .A(n_264), .B(n_1315), .Y(n_1314) );
INVxp67_ASAP7_75t_SL g896 ( .A(n_267), .Y(n_896) );
INVx1_ASAP7_75t_L g364 ( .A(n_269), .Y(n_364) );
INVx1_ASAP7_75t_L g382 ( .A(n_269), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g1334 ( .A1(n_270), .A2(n_307), .B1(n_511), .B2(n_602), .C(n_936), .Y(n_1334) );
INVx1_ASAP7_75t_L g561 ( .A(n_271), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g1235 ( .A(n_272), .Y(n_1235) );
INVx1_ASAP7_75t_L g1480 ( .A(n_273), .Y(n_1480) );
INVxp67_ASAP7_75t_SL g1505 ( .A(n_274), .Y(n_1505) );
INVx1_ASAP7_75t_L g899 ( .A(n_275), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_276), .A2(n_312), .B1(n_417), .B2(n_420), .Y(n_872) );
INVx1_ASAP7_75t_L g897 ( .A(n_276), .Y(n_897) );
INVx1_ASAP7_75t_L g1409 ( .A(n_277), .Y(n_1409) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_278), .Y(n_455) );
AOI21xp33_ASAP7_75t_L g747 ( .A1(n_279), .A2(n_559), .B(n_748), .Y(n_747) );
INVxp67_ASAP7_75t_L g771 ( .A(n_279), .Y(n_771) );
INVx1_ASAP7_75t_L g1410 ( .A(n_281), .Y(n_1410) );
INVx1_ASAP7_75t_L g1052 ( .A(n_283), .Y(n_1052) );
NOR2xp33_ASAP7_75t_L g1055 ( .A(n_283), .B(n_760), .Y(n_1055) );
INVx1_ASAP7_75t_L g1271 ( .A(n_284), .Y(n_1271) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_285), .Y(n_1006) );
INVx1_ASAP7_75t_L g1404 ( .A(n_286), .Y(n_1404) );
AOI22xp5_ASAP7_75t_SL g1554 ( .A1(n_287), .A2(n_337), .B1(n_1528), .B2(n_1532), .Y(n_1554) );
INVxp33_ASAP7_75t_L g838 ( .A(n_288), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_289), .Y(n_943) );
INVx1_ASAP7_75t_L g848 ( .A(n_290), .Y(n_848) );
INVx1_ASAP7_75t_L g1118 ( .A(n_291), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_292), .B(n_1531), .Y(n_1530) );
INVx1_ASAP7_75t_L g1537 ( .A(n_292), .Y(n_1537) );
CKINVDCx5p33_ASAP7_75t_R g1342 ( .A(n_293), .Y(n_1342) );
OAI22xp33_ASAP7_75t_L g1370 ( .A1(n_296), .A2(n_343), .B1(n_1371), .B2(n_1374), .Y(n_1370) );
OAI22xp33_ASAP7_75t_L g1451 ( .A1(n_296), .A2(n_343), .B1(n_1452), .B2(n_1454), .Y(n_1451) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_298), .A2(n_602), .B(n_715), .Y(n_714) );
XOR2x2_ASAP7_75t_L g726 ( .A(n_300), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g628 ( .A(n_301), .Y(n_628) );
INVx1_ASAP7_75t_L g1850 ( .A(n_302), .Y(n_1850) );
CKINVDCx5p33_ASAP7_75t_R g1775 ( .A(n_303), .Y(n_1775) );
INVx1_ASAP7_75t_L g1155 ( .A(n_304), .Y(n_1155) );
INVx1_ASAP7_75t_L g1220 ( .A(n_306), .Y(n_1220) );
INVx1_ASAP7_75t_L g1099 ( .A(n_308), .Y(n_1099) );
OAI221xp5_ASAP7_75t_L g1132 ( .A1(n_308), .A2(n_488), .B1(n_610), .B2(n_1133), .C(n_1141), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_310), .A2(n_320), .B1(n_1188), .B2(n_1190), .Y(n_1498) );
INVx1_ASAP7_75t_L g814 ( .A(n_311), .Y(n_814) );
INVxp67_ASAP7_75t_SL g919 ( .A(n_312), .Y(n_919) );
INVx1_ASAP7_75t_L g1387 ( .A(n_313), .Y(n_1387) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_314), .Y(n_450) );
INVx1_ASAP7_75t_L g739 ( .A(n_315), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g988 ( .A(n_317), .Y(n_988) );
CKINVDCx5p33_ASAP7_75t_R g1285 ( .A(n_318), .Y(n_1285) );
INVx1_ASAP7_75t_L g913 ( .A(n_319), .Y(n_913) );
AOI21xp33_ASAP7_75t_L g510 ( .A1(n_322), .A2(n_511), .B(n_514), .Y(n_510) );
INVx1_ASAP7_75t_L g552 ( .A(n_323), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g1233 ( .A(n_324), .Y(n_1233) );
INVx1_ASAP7_75t_L g1081 ( .A(n_326), .Y(n_1081) );
XOR2xp5_ASAP7_75t_L g981 ( .A(n_327), .B(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g437 ( .A(n_328), .Y(n_437) );
INVx1_ASAP7_75t_L g444 ( .A(n_328), .Y(n_444) );
INVx1_ASAP7_75t_L g466 ( .A(n_328), .Y(n_466) );
INVx1_ASAP7_75t_L g883 ( .A(n_329), .Y(n_883) );
INVx1_ASAP7_75t_L g472 ( .A(n_330), .Y(n_472) );
INVx1_ASAP7_75t_L g698 ( .A(n_331), .Y(n_698) );
INVx1_ASAP7_75t_L g1274 ( .A(n_332), .Y(n_1274) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_334), .Y(n_1101) );
INVxp67_ASAP7_75t_SL g766 ( .A(n_335), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_336), .Y(n_795) );
AOI21xp33_ASAP7_75t_L g1776 ( .A1(n_340), .A2(n_497), .B(n_946), .Y(n_1776) );
INVx1_ASAP7_75t_L g1796 ( .A(n_340), .Y(n_1796) );
INVx1_ASAP7_75t_L g1406 ( .A(n_341), .Y(n_1406) );
CKINVDCx5p33_ASAP7_75t_R g1760 ( .A(n_342), .Y(n_1760) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_1508), .B(n_1520), .Y(n_344) );
XNOR2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_1359), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_1314), .B2(n_1358), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI22x1_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B1(n_979), .B2(n_1312), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
XOR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_788), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_631), .B1(n_632), .B2(n_787), .Y(n_351) );
INVx1_ASAP7_75t_L g787 ( .A(n_352), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_541), .B1(n_542), .B2(n_630), .Y(n_352) );
INVx2_ASAP7_75t_L g630 ( .A(n_353), .Y(n_630) );
NOR2x1_ASAP7_75t_L g354 ( .A(n_355), .B(n_453), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_399), .B(n_435), .C(n_438), .Y(n_355) );
AOI211xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_370), .B(n_371), .C(n_388), .Y(n_356) );
AOI211xp5_ASAP7_75t_L g729 ( .A1(n_357), .A2(n_730), .B(n_731), .C(n_732), .Y(n_729) );
AOI211xp5_ASAP7_75t_SL g884 ( .A1(n_357), .A2(n_885), .B(n_886), .C(n_887), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_357), .A2(n_1047), .B1(n_1049), .B2(n_1054), .Y(n_1046) );
AOI221xp5_ASAP7_75t_L g1257 ( .A1(n_357), .A2(n_548), .B1(n_1252), .B2(n_1258), .C(n_1259), .Y(n_1257) );
AOI221xp5_ASAP7_75t_L g1291 ( .A1(n_357), .A2(n_548), .B1(n_1292), .B2(n_1293), .C(n_1297), .Y(n_1291) );
INVx2_ASAP7_75t_L g1504 ( .A(n_357), .Y(n_1504) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g647 ( .A(n_358), .B(n_648), .Y(n_647) );
OR2x6_ASAP7_75t_L g859 ( .A(n_358), .B(n_648), .Y(n_859) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_359), .B(n_365), .Y(n_358) );
BUFx3_ASAP7_75t_L g412 ( .A(n_359), .Y(n_412) );
AND2x2_ASAP7_75t_L g418 ( .A(n_359), .B(n_419), .Y(n_418) );
INVx8_ASAP7_75t_L g563 ( .A(n_359), .Y(n_563) );
BUFx3_ASAP7_75t_L g751 ( .A(n_359), .Y(n_751) );
HB1xp67_ASAP7_75t_L g1202 ( .A(n_359), .Y(n_1202) );
AND2x4_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
AND2x4_ASAP7_75t_L g394 ( .A(n_360), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_361), .Y(n_376) );
AND2x4_ASAP7_75t_L g422 ( .A(n_361), .B(n_381), .Y(n_422) );
OR2x2_ASAP7_75t_L g430 ( .A(n_361), .B(n_363), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_361), .B(n_382), .Y(n_576) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g395 ( .A(n_364), .Y(n_395) );
AND2x6_ASAP7_75t_L g373 ( .A(n_365), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g378 ( .A(n_365), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g387 ( .A(n_365), .Y(n_387) );
AND2x4_ASAP7_75t_L g654 ( .A(n_365), .B(n_522), .Y(n_654) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g433 ( .A(n_366), .B(n_434), .Y(n_433) );
NAND3x1_ASAP7_75t_L g854 ( .A(n_366), .B(n_434), .C(n_855), .Y(n_854) );
OR2x4_ASAP7_75t_L g1373 ( .A(n_366), .B(n_430), .Y(n_1373) );
INVx1_ASAP7_75t_L g1376 ( .A(n_366), .Y(n_1376) );
AND2x4_ASAP7_75t_L g1381 ( .A(n_366), .B(n_422), .Y(n_1381) );
OR2x6_ASAP7_75t_L g1397 ( .A(n_366), .B(n_575), .Y(n_1397) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g415 ( .A(n_367), .Y(n_415) );
NAND2xp33_ASAP7_75t_SL g749 ( .A(n_367), .B(n_369), .Y(n_749) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g414 ( .A(n_369), .B(n_415), .Y(n_414) );
AND3x4_ASAP7_75t_L g662 ( .A(n_369), .B(n_415), .C(n_436), .Y(n_662) );
HB1xp67_ASAP7_75t_L g1366 ( .A(n_369), .Y(n_1366) );
INVx4_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g1042 ( .A1(n_373), .A2(n_378), .B1(n_1043), .B2(n_1044), .C(n_1045), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_373), .A2(n_378), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
AND2x2_ASAP7_75t_L g653 ( .A(n_374), .B(n_654), .Y(n_653) );
NAND2x1_ASAP7_75t_L g865 ( .A(n_374), .B(n_654), .Y(n_865) );
AND2x4_ASAP7_75t_SL g970 ( .A(n_374), .B(n_654), .Y(n_970) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_374), .B(n_654), .Y(n_1346) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_376), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g398 ( .A(n_376), .B(n_380), .Y(n_398) );
BUFx2_ASAP7_75t_L g1386 ( .A(n_376), .Y(n_1386) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g1493 ( .A(n_378), .Y(n_1493) );
INVx1_ASAP7_75t_L g565 ( .A(n_379), .Y(n_565) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g386 ( .A(n_382), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g1045 ( .A(n_383), .Y(n_1045) );
OR2x6_ASAP7_75t_L g383 ( .A(n_384), .B(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g426 ( .A(n_384), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g1284 ( .A1(n_384), .A2(n_432), .B1(n_841), .B2(n_1285), .C(n_1286), .Y(n_1284) );
INVx1_ASAP7_75t_L g1379 ( .A(n_384), .Y(n_1379) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_385), .Y(n_407) );
BUFx3_ASAP7_75t_L g876 ( .A(n_385), .Y(n_876) );
BUFx2_ASAP7_75t_L g1390 ( .A(n_386), .Y(n_1390) );
INVx1_ASAP7_75t_L g567 ( .A(n_387), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_389), .Y(n_753) );
OR2x6_ASAP7_75t_SL g389 ( .A(n_390), .B(n_393), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g397 ( .A(n_391), .B(n_398), .Y(n_397) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_391), .Y(n_549) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g419 ( .A(n_392), .Y(n_419) );
OR2x2_ASAP7_75t_L g642 ( .A(n_392), .B(n_530), .Y(n_642) );
INVx1_ASAP7_75t_L g832 ( .A(n_393), .Y(n_832) );
INVx3_ASAP7_75t_L g1175 ( .A(n_393), .Y(n_1175) );
BUFx2_ASAP7_75t_L g1801 ( .A(n_393), .Y(n_1801) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_394), .Y(n_403) );
BUFx8_ASAP7_75t_L g431 ( .A(n_394), .Y(n_431) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_394), .Y(n_559) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_397), .A2(n_753), .B1(n_754), .B2(n_755), .C(n_756), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_397), .B(n_598), .Y(n_1145) );
INVx5_ASAP7_75t_L g409 ( .A(n_398), .Y(n_409) );
BUFx3_ASAP7_75t_L g551 ( .A(n_398), .Y(n_551) );
BUFx3_ASAP7_75t_L g999 ( .A(n_398), .Y(n_999) );
BUFx2_ASAP7_75t_L g1034 ( .A(n_398), .Y(n_1034) );
BUFx12f_ASAP7_75t_L g1188 ( .A(n_398), .Y(n_1188) );
NOR3xp33_ASAP7_75t_SL g399 ( .A(n_400), .B(n_416), .C(n_423), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_403), .Y(n_594) );
BUFx6f_ASAP7_75t_L g846 ( .A(n_403), .Y(n_846) );
INVx2_ASAP7_75t_L g1282 ( .A(n_403), .Y(n_1282) );
AND2x4_ASAP7_75t_L g1375 ( .A(n_403), .B(n_1376), .Y(n_1375) );
INVx2_ASAP7_75t_L g1501 ( .A(n_403), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1791 ( .A(n_403), .B(n_1376), .Y(n_1791) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g579 ( .A(n_406), .Y(n_579) );
INVx1_ASAP7_75t_L g592 ( .A(n_406), .Y(n_592) );
INVx2_ASAP7_75t_L g1782 ( .A(n_406), .Y(n_1782) );
INVx4_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_407), .Y(n_566) );
OR2x2_ASAP7_75t_L g646 ( .A(n_407), .B(n_642), .Y(n_646) );
INVx3_ASAP7_75t_L g746 ( .A(n_407), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g1279 ( .A1(n_407), .A2(n_414), .B1(n_1280), .B2(n_1281), .C(n_1282), .Y(n_1279) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_411), .B2(n_413), .C(n_414), .Y(n_408) );
INVx2_ASAP7_75t_L g666 ( .A(n_409), .Y(n_666) );
INVx2_ASAP7_75t_R g668 ( .A(n_409), .Y(n_668) );
INVx1_ASAP7_75t_L g1108 ( .A(n_409), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_410), .A2(n_537), .B1(n_539), .B2(n_540), .Y(n_536) );
INVx2_ASAP7_75t_L g1033 ( .A(n_411), .Y(n_1033) );
INVx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g994 ( .A(n_412), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_412), .B(n_1296), .Y(n_1295) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_413), .A2(n_500), .B1(n_504), .B2(n_505), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_414), .A2(n_591), .B1(n_592), .B2(n_593), .C(n_595), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g875 ( .A1(n_414), .A2(n_558), .B1(n_876), .B2(n_877), .C(n_878), .Y(n_875) );
OAI221xp5_ASAP7_75t_L g1264 ( .A1(n_414), .A2(n_876), .B1(n_1237), .B2(n_1241), .C(n_1265), .Y(n_1264) );
INVx3_ASAP7_75t_L g1385 ( .A(n_415), .Y(n_1385) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g421 ( .A(n_419), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g554 ( .A(n_422), .Y(n_554) );
BUFx2_ASAP7_75t_L g661 ( .A(n_422), .Y(n_661) );
BUFx2_ASAP7_75t_L g681 ( .A(n_422), .Y(n_681) );
BUFx2_ASAP7_75t_L g850 ( .A(n_422), .Y(n_850) );
BUFx2_ASAP7_75t_L g995 ( .A(n_422), .Y(n_995) );
BUFx3_ASAP7_75t_L g1040 ( .A(n_422), .Y(n_1040) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .Y(n_427) );
INVx3_ASAP7_75t_L g585 ( .A(n_429), .Y(n_585) );
INVx2_ASAP7_75t_SL g674 ( .A(n_429), .Y(n_674) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g557 ( .A(n_430), .Y(n_557) );
BUFx3_ASAP7_75t_L g580 ( .A(n_430), .Y(n_580) );
BUFx4f_ASAP7_75t_L g841 ( .A(n_430), .Y(n_841) );
OR2x4_ASAP7_75t_L g1394 ( .A(n_430), .B(n_1376), .Y(n_1394) );
AND2x4_ASAP7_75t_L g678 ( .A(n_431), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g738 ( .A(n_431), .Y(n_738) );
INVx3_ASAP7_75t_L g954 ( .A(n_431), .Y(n_954) );
INVx3_ASAP7_75t_L g1106 ( .A(n_431), .Y(n_1106) );
INVx2_ASAP7_75t_SL g1116 ( .A(n_431), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1356 ( .A(n_431), .Y(n_1356) );
OAI221xp5_ASAP7_75t_L g577 ( .A1(n_432), .A2(n_578), .B1(n_579), .B2(n_580), .C(n_581), .Y(n_577) );
INVx3_ASAP7_75t_L g736 ( .A(n_432), .Y(n_736) );
OAI221xp5_ASAP7_75t_L g881 ( .A1(n_432), .A2(n_841), .B1(n_876), .B2(n_882), .C(n_883), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g1110 ( .A1(n_432), .A2(n_839), .B1(n_1111), .B2(n_1113), .C(n_1114), .Y(n_1110) );
OAI221xp5_ASAP7_75t_L g1267 ( .A1(n_432), .A2(n_557), .B1(n_876), .B2(n_1233), .C(n_1242), .Y(n_1267) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x6_ASAP7_75t_L g670 ( .A(n_433), .B(n_516), .Y(n_670) );
OR2x2_ASAP7_75t_L g1859 ( .A(n_433), .B(n_516), .Y(n_1859) );
O2A1O1Ixp5_ASAP7_75t_L g1316 ( .A1(n_435), .A2(n_1317), .B(n_1332), .C(n_1339), .Y(n_1316) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g724 ( .A(n_436), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g1488 ( .A1(n_436), .A2(n_892), .B1(n_1489), .B2(n_1505), .Y(n_1488) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_437), .B(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g516 ( .A(n_437), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_440), .A2(n_456), .B1(n_628), .B2(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_440), .B(n_754), .Y(n_786) );
INVx1_ASAP7_75t_L g893 ( .A(n_440), .Y(n_893) );
HB1xp67_ASAP7_75t_L g1061 ( .A(n_440), .Y(n_1061) );
AOI222xp33_ASAP7_75t_L g1086 ( .A1(n_440), .A2(n_456), .B1(n_1087), .B2(n_1088), .C1(n_1090), .C2(n_1091), .Y(n_1086) );
NAND2xp33_ASAP7_75t_SL g1270 ( .A(n_440), .B(n_1271), .Y(n_1270) );
AND2x4_ASAP7_75t_L g440 ( .A(n_441), .B(n_445), .Y(n_440) );
AND2x4_ASAP7_75t_L g456 ( .A(n_441), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g483 ( .A(n_442), .B(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g622 ( .A(n_442), .B(n_484), .Y(n_622) );
INVxp67_ASAP7_75t_L g648 ( .A(n_442), .Y(n_648) );
INVx1_ASAP7_75t_L g1459 ( .A(n_442), .Y(n_1459) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g530 ( .A(n_443), .Y(n_530) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
AND2x2_ASAP7_75t_L g457 ( .A(n_446), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_446), .B(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g685 ( .A(n_446), .B(n_686), .Y(n_685) );
AND2x4_ASAP7_75t_L g699 ( .A(n_446), .B(n_448), .Y(n_699) );
AND2x4_ASAP7_75t_SL g704 ( .A(n_446), .B(n_512), .Y(n_704) );
AND2x2_ASAP7_75t_L g928 ( .A(n_446), .B(n_467), .Y(n_928) );
BUFx2_ASAP7_75t_L g1821 ( .A(n_446), .Y(n_1821) );
HB1xp67_ASAP7_75t_L g1447 ( .A(n_447), .Y(n_1447) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_448), .Y(n_497) );
INVx2_ASAP7_75t_L g801 ( .A(n_448), .Y(n_801) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx3_ASAP7_75t_L g535 ( .A(n_449), .Y(n_535) );
INVx2_ASAP7_75t_L g605 ( .A(n_449), .Y(n_605) );
AND2x4_ASAP7_75t_L g1455 ( .A(n_449), .B(n_1447), .Y(n_1455) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx2_ASAP7_75t_L g459 ( .A(n_450), .Y(n_459) );
INVx2_ASAP7_75t_L g470 ( .A(n_450), .Y(n_470) );
INVx1_ASAP7_75t_L g486 ( .A(n_450), .Y(n_486) );
NAND2x1_ASAP7_75t_L g490 ( .A(n_450), .B(n_452), .Y(n_490) );
OR2x2_ASAP7_75t_L g503 ( .A(n_450), .B(n_452), .Y(n_503) );
AND2x2_ASAP7_75t_L g513 ( .A(n_450), .B(n_452), .Y(n_513) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g460 ( .A(n_452), .Y(n_460) );
AND2x2_ASAP7_75t_L g469 ( .A(n_452), .B(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g480 ( .A(n_452), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_452), .B(n_470), .Y(n_509) );
OR2x2_ASAP7_75t_L g614 ( .A(n_452), .B(n_459), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_494), .Y(n_453) );
AOI211xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B(n_461), .C(n_487), .Y(n_454) );
INVx3_ASAP7_75t_L g760 ( .A(n_456), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_456), .B(n_919), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_456), .B(n_1255), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_456), .B(n_1296), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_456), .B(n_1468), .Y(n_1467) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_457), .Y(n_697) );
INVx1_ASAP7_75t_L g810 ( .A(n_457), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_458), .B(n_477), .Y(n_524) );
INVx3_ASAP7_75t_L g618 ( .A(n_458), .Y(n_618) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_458), .Y(n_720) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI222xp33_ASAP7_75t_L g782 ( .A1(n_463), .A2(n_520), .B1(n_730), .B2(n_755), .C1(n_783), .C2(n_785), .Y(n_782) );
AOI222xp33_ASAP7_75t_L g895 ( .A1(n_463), .A2(n_473), .B1(n_482), .B2(n_885), .C1(n_896), .C2(n_897), .Y(n_895) );
INVxp67_ASAP7_75t_L g1058 ( .A(n_463), .Y(n_1058) );
INVx1_ASAP7_75t_L g1089 ( .A(n_463), .Y(n_1089) );
AOI222xp33_ASAP7_75t_L g1250 ( .A1(n_463), .A2(n_520), .B1(n_783), .B2(n_1251), .C1(n_1252), .C2(n_1253), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1471 ( .A1(n_463), .A2(n_783), .B1(n_1472), .B2(n_1473), .Y(n_1471) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_467), .Y(n_463) );
AOI332xp33_ASAP7_75t_L g1300 ( .A1(n_464), .A2(n_467), .A3(n_521), .B1(n_523), .B2(n_783), .B3(n_1292), .C1(n_1301), .C2(n_1302), .Y(n_1300) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g488 ( .A(n_465), .B(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g784 ( .A(n_465), .B(n_489), .Y(n_784) );
INVx1_ASAP7_75t_L g522 ( .A(n_466), .Y(n_522) );
INVx1_ASAP7_75t_L g855 ( .A(n_466), .Y(n_855) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g949 ( .A(n_468), .Y(n_949) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_469), .Y(n_686) );
BUFx3_ASAP7_75t_L g805 ( .A(n_469), .Y(n_805) );
BUFx3_ASAP7_75t_L g939 ( .A(n_469), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_481), .B2(n_482), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_473), .A2(n_482), .B1(n_1096), .B2(n_1098), .Y(n_1141) );
AOI22xp33_ASAP7_75t_SL g1478 ( .A1(n_473), .A2(n_482), .B1(n_1479), .B2(n_1480), .Y(n_1478) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_SL g621 ( .A(n_474), .Y(n_621) );
NAND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_478), .Y(n_474) );
INVx1_ASAP7_75t_L g493 ( .A(n_475), .Y(n_493) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_477), .B(n_485), .Y(n_484) );
AND2x6_ASAP7_75t_L g694 ( .A(n_477), .B(n_512), .Y(n_694) );
INVx1_ASAP7_75t_L g709 ( .A(n_477), .Y(n_709) );
AND2x2_ASAP7_75t_L g806 ( .A(n_477), .B(n_807), .Y(n_806) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g708 ( .A(n_480), .Y(n_708) );
BUFx2_ASAP7_75t_L g807 ( .A(n_480), .Y(n_807) );
AND2x4_ASAP7_75t_L g1437 ( .A(n_480), .B(n_1438), .Y(n_1437) );
AND2x2_ASAP7_75t_L g1758 ( .A(n_480), .B(n_1434), .Y(n_1758) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
AND2x4_ASAP7_75t_L g645 ( .A(n_483), .B(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g794 ( .A(n_483), .B(n_646), .Y(n_794) );
INVx1_ASAP7_75t_L g1828 ( .A(n_484), .Y(n_1828) );
AND2x4_ASAP7_75t_L g1442 ( .A(n_485), .B(n_518), .Y(n_1442) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx3_ASAP7_75t_L g608 ( .A(n_489), .Y(n_608) );
INVx2_ASAP7_75t_SL g1321 ( .A(n_489), .Y(n_1321) );
BUFx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_490), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_491), .A2(n_610), .B(n_611), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g922 ( .A(n_491), .Y(n_922) );
OAI21xp5_ASAP7_75t_L g1069 ( .A1(n_491), .A2(n_1070), .B(n_1078), .Y(n_1069) );
OAI21xp5_ASAP7_75t_SL g1120 ( .A1(n_491), .A2(n_1121), .B(n_1125), .Y(n_1120) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx4_ASAP7_75t_L g713 ( .A(n_492), .Y(n_713) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_492), .Y(n_774) );
BUFx4f_ASAP7_75t_L g944 ( .A(n_492), .Y(n_944) );
BUFx4f_ASAP7_75t_L g1129 ( .A(n_492), .Y(n_1129) );
BUFx4f_ASAP7_75t_L g1137 ( .A(n_492), .Y(n_1137) );
AOI322xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .A3(n_510), .B1(n_519), .B2(n_520), .C1(n_525), .C2(n_531), .Y(n_494) );
BUFx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g1231 ( .A1(n_500), .A2(n_917), .B1(n_1232), .B2(n_1233), .Y(n_1231) );
OAI22xp5_ASAP7_75t_L g1767 ( .A1(n_500), .A2(n_505), .B1(n_1768), .B2(n_1769), .Y(n_1767) );
BUFx4f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g915 ( .A(n_501), .Y(n_915) );
INVxp67_ASAP7_75t_L g1245 ( .A(n_501), .Y(n_1245) );
OR2x6_ASAP7_75t_L g1446 ( .A(n_501), .B(n_1447), .Y(n_1446) );
OR2x6_ASAP7_75t_L g1452 ( .A(n_501), .B(n_1453), .Y(n_1452) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g538 ( .A(n_502), .Y(n_538) );
BUFx4f_ASAP7_75t_L g908 ( .A(n_502), .Y(n_908) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g1400 ( .A1(n_505), .A2(n_1401), .B1(n_1402), .B2(n_1404), .Y(n_1400) );
INVx5_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx6_ASAP7_75t_L g615 ( .A(n_506), .Y(n_615) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g540 ( .A(n_507), .Y(n_540) );
INVx4_ASAP7_75t_L g909 ( .A(n_507), .Y(n_909) );
INVx2_ASAP7_75t_SL g917 ( .A(n_507), .Y(n_917) );
INVx1_ASAP7_75t_L g1163 ( .A(n_507), .Y(n_1163) );
INVx2_ASAP7_75t_L g1329 ( .A(n_507), .Y(n_1329) );
INVx8_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g769 ( .A(n_508), .Y(n_769) );
OR2x2_ASAP7_75t_L g1450 ( .A(n_508), .B(n_1438), .Y(n_1450) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g1818 ( .A1(n_511), .A2(n_805), .B1(n_1819), .B2(n_1820), .Y(n_1818) );
A2O1A1Ixp33_ASAP7_75t_L g1823 ( .A1(n_511), .A2(n_1139), .B(n_1824), .C(n_1825), .Y(n_1823) );
BUFx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_512), .Y(n_533) );
BUFx3_ASAP7_75t_L g689 ( .A(n_512), .Y(n_689) );
INVx1_ASAP7_75t_L g902 ( .A(n_512), .Y(n_902) );
BUFx3_ASAP7_75t_L g911 ( .A(n_512), .Y(n_911) );
BUFx3_ASAP7_75t_L g934 ( .A(n_512), .Y(n_934) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_512), .B(n_1434), .Y(n_1433) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g1012 ( .A(n_513), .Y(n_1012) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_515), .Y(n_600) );
INVx2_ASAP7_75t_L g764 ( .A(n_515), .Y(n_764) );
AOI222xp33_ASAP7_75t_L g898 ( .A1(n_515), .A2(n_520), .B1(n_525), .B2(n_899), .C1(n_900), .C2(n_910), .Y(n_898) );
INVx2_ASAP7_75t_L g1079 ( .A(n_515), .Y(n_1079) );
INVx4_ASAP7_75t_L g1124 ( .A(n_515), .Y(n_1124) );
AOI31xp33_ASAP7_75t_L g1475 ( .A1(n_515), .A2(n_922), .A3(n_1476), .B(n_1477), .Y(n_1475) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g598 ( .A(n_516), .Y(n_598) );
AND2x4_ASAP7_75t_L g526 ( .A(n_518), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g717 ( .A(n_518), .Y(n_717) );
BUFx2_ASAP7_75t_L g1438 ( .A(n_518), .Y(n_1438) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g626 ( .A(n_522), .B(n_524), .Y(n_626) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_525), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g1062 ( .A1(n_525), .A2(n_1063), .B(n_1069), .C(n_1080), .Y(n_1062) );
NAND3xp33_ASAP7_75t_L g1481 ( .A(n_525), .B(n_1482), .C(n_1485), .Y(n_1481) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_528), .Y(n_525) );
INVx1_ASAP7_75t_SL g690 ( .A(n_526), .Y(n_690) );
AND2x2_ASAP7_75t_SL g780 ( .A(n_526), .B(n_530), .Y(n_780) );
INVx4_ASAP7_75t_L g819 ( .A(n_526), .Y(n_819) );
INVx4_ASAP7_75t_L g936 ( .A(n_526), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_526), .B(n_528), .Y(n_1307) );
OAI221xp5_ASAP7_75t_L g1770 ( .A1(n_526), .A2(n_1239), .B1(n_1771), .B2(n_1772), .C(n_1773), .Y(n_1770) );
AND2x4_ASAP7_75t_L g716 ( .A(n_527), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g1458 ( .A(n_527), .Y(n_1458) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g836 ( .A(n_530), .B(n_749), .Y(n_836) );
HB1xp67_ASAP7_75t_L g1368 ( .A(n_530), .Y(n_1368) );
BUFx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g904 ( .A(n_535), .Y(n_904) );
BUFx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g607 ( .A(n_538), .Y(n_607) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_538), .Y(n_767) );
INVx2_ASAP7_75t_SL g777 ( .A(n_538), .Y(n_777) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND4xp75_ASAP7_75t_L g544 ( .A(n_545), .B(n_599), .C(n_623), .D(n_627), .Y(n_544) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_568), .B(n_596), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_550), .B(n_560), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g1499 ( .A1(n_548), .A2(n_1472), .B1(n_1500), .B2(n_1503), .Y(n_1499) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g1048 ( .A(n_549), .Y(n_1048) );
AOI221xp5_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_552), .B1(n_553), .B2(n_555), .C(n_556), .Y(n_550) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g965 ( .A(n_554), .Y(n_965) );
INVx2_ASAP7_75t_L g1203 ( .A(n_554), .Y(n_1203) );
INVx1_ASAP7_75t_L g1422 ( .A(n_557), .Y(n_1422) );
INVx2_ASAP7_75t_L g997 ( .A(n_558), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g1424 ( .A1(n_558), .A2(n_1406), .B1(n_1415), .B2(n_1425), .Y(n_1424) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_559), .Y(n_572) );
INVx5_ASAP7_75t_L g665 ( .A(n_559), .Y(n_665) );
INVx2_ASAP7_75t_SL g1038 ( .A(n_559), .Y(n_1038) );
INVx3_ASAP7_75t_L g1050 ( .A(n_559), .Y(n_1050) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B(n_564), .C(n_567), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g1502 ( .A1(n_562), .A2(n_681), .B1(n_1468), .B2(n_1480), .Y(n_1502) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx8_ASAP7_75t_L g660 ( .A(n_563), .Y(n_660) );
INVx2_ASAP7_75t_L g874 ( .A(n_563), .Y(n_874) );
INVx2_ASAP7_75t_L g978 ( .A(n_563), .Y(n_978) );
INVx2_ASAP7_75t_L g657 ( .A(n_565), .Y(n_657) );
HB1xp67_ASAP7_75t_L g1423 ( .A(n_566), .Y(n_1423) );
OAI22xp33_ASAP7_75t_L g1846 ( .A1(n_566), .A2(n_841), .B1(n_1847), .B2(n_1848), .Y(n_1846) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_577), .B1(n_582), .B2(n_590), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B1(n_573), .B2(n_574), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_570), .A2(n_583), .B1(n_607), .B2(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_573), .A2(n_591), .B1(n_612), .B2(n_615), .C(n_616), .Y(n_611) );
OAI221xp5_ASAP7_75t_L g844 ( .A1(n_574), .A2(n_845), .B1(n_847), .B2(n_848), .C(n_849), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g1426 ( .A1(n_574), .A2(n_1265), .B1(n_1407), .B2(n_1416), .Y(n_1426) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g589 ( .A(n_575), .Y(n_589) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g641 ( .A(n_576), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B1(n_586), .B2(n_587), .Y(n_582) );
BUFx4f_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
OAI21xp33_ASAP7_75t_L g957 ( .A1(n_587), .A2(n_958), .B(n_959), .Y(n_957) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g1851 ( .A(n_589), .Y(n_1851) );
OAI21xp33_ASAP7_75t_L g733 ( .A1(n_592), .A2(n_734), .B(n_735), .Y(n_733) );
OAI221xp5_ASAP7_75t_L g960 ( .A1(n_593), .A2(n_943), .B1(n_961), .B2(n_963), .C(n_964), .Y(n_960) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_SL g1797 ( .A(n_594), .Y(n_1797) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx2_ASAP7_75t_L g889 ( .A(n_598), .Y(n_889) );
AOI21xp5_ASAP7_75t_SL g1814 ( .A1(n_598), .A2(n_1815), .B(n_1830), .Y(n_1814) );
AOI211x1_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B(n_609), .C(n_619), .Y(n_599) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g1016 ( .A(n_603), .Y(n_1016) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g817 ( .A(n_604), .Y(n_817) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g1064 ( .A(n_605), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_608), .A2(n_612), .B1(n_739), .B2(n_771), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g1238 ( .A1(n_608), .A2(n_1239), .B1(n_1241), .B2(n_1242), .Y(n_1238) );
BUFx2_ASAP7_75t_L g1431 ( .A(n_608), .Y(n_1431) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx2_ASAP7_75t_L g773 ( .A(n_614), .Y(n_773) );
BUFx3_ASAP7_75t_L g1073 ( .A(n_614), .Y(n_1073) );
INVx2_ASAP7_75t_L g1127 ( .A(n_614), .Y(n_1127) );
BUFx2_ASAP7_75t_L g1136 ( .A(n_614), .Y(n_1136) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_615), .A2(n_1066), .B1(n_1067), .B2(n_1068), .Y(n_1065) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g692 ( .A(n_618), .Y(n_692) );
INVx2_ASAP7_75t_SL g938 ( .A(n_618), .Y(n_938) );
INVx1_ASAP7_75t_L g948 ( .A(n_618), .Y(n_948) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g638 ( .A(n_626), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_626), .B(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_725), .B2(n_726), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND3xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_649), .C(n_682), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_643), .B(n_644), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_637), .A2(n_825), .B1(n_858), .B2(n_860), .C(n_861), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g973 ( .A1(n_637), .A2(n_974), .B(n_975), .Y(n_973) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_637), .A2(n_858), .B1(n_984), .B2(n_985), .C(n_986), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_637), .B(n_1178), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_637), .A2(n_858), .B1(n_1197), .B2(n_1198), .C(n_1199), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_637), .B(n_1342), .Y(n_1341) );
INVx8_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g741 ( .A(n_640), .Y(n_741) );
BUFx3_ASAP7_75t_L g834 ( .A(n_640), .Y(n_834) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx6f_ASAP7_75t_L g962 ( .A(n_641), .Y(n_962) );
INVx1_ASAP7_75t_L g676 ( .A(n_642), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_642), .Y(n_679) );
INVx2_ASAP7_75t_L g1840 ( .A(n_646), .Y(n_1840) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_647), .B(n_1089), .Y(n_1088) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_672), .C(n_680), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_658), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_655), .B2(n_656), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_653), .A2(n_656), .B1(n_1208), .B2(n_1209), .Y(n_1207) );
AND2x4_ASAP7_75t_L g656 ( .A(n_654), .B(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g680 ( .A(n_654), .B(n_681), .Y(n_680) );
AND2x4_ASAP7_75t_SL g972 ( .A(n_654), .B(n_657), .Y(n_972) );
A2O1A1Ixp33_ASAP7_75t_L g1843 ( .A1(n_654), .A2(n_660), .B(n_1819), .C(n_1844), .Y(n_1843) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_656), .A2(n_808), .B1(n_814), .B2(n_864), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_656), .A2(n_864), .B1(n_988), .B2(n_989), .Y(n_987) );
AOI22xp5_ASAP7_75t_L g1344 ( .A1(n_656), .A2(n_1345), .B1(n_1346), .B2(n_1347), .Y(n_1344) );
AOI33xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .A3(n_663), .B1(n_667), .B2(n_669), .B3(n_671), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_660), .A2(n_850), .B1(n_1090), .B2(n_1096), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_661), .A2(n_874), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
BUFx3_ASAP7_75t_L g991 ( .A(n_662), .Y(n_991) );
AOI33xp33_ASAP7_75t_L g1185 ( .A1(n_662), .A2(n_1186), .A3(n_1187), .B1(n_1189), .B2(n_1191), .B3(n_1192), .Y(n_1185) );
AOI33xp33_ASAP7_75t_L g1200 ( .A1(n_662), .A2(n_669), .A3(n_1201), .B1(n_1204), .B2(n_1205), .B3(n_1206), .Y(n_1200) );
INVx8_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g1849 ( .A1(n_665), .A2(n_1850), .B1(n_1851), .B2(n_1852), .Y(n_1849) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
OR2x6_ASAP7_75t_L g862 ( .A(n_674), .B(n_675), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g1428 ( .A1(n_674), .A2(n_843), .B1(n_1404), .B2(n_1410), .Y(n_1428) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_676), .B(n_1175), .Y(n_1174) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g856 ( .A(n_678), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_678), .A2(n_930), .B1(n_931), .B2(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_678), .A2(n_1005), .B1(n_1006), .B2(n_1024), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_678), .A2(n_1024), .B1(n_1337), .B2(n_1338), .Y(n_1340) );
AND2x4_ASAP7_75t_L g977 ( .A(n_679), .B(n_978), .Y(n_977) );
AND2x4_ASAP7_75t_L g1024 ( .A(n_679), .B(n_978), .Y(n_1024) );
INVx3_ASAP7_75t_L g866 ( .A(n_680), .Y(n_866) );
NOR3xp33_ASAP7_75t_L g951 ( .A(n_680), .B(n_952), .C(n_968), .Y(n_951) );
INVx3_ASAP7_75t_L g1193 ( .A(n_680), .Y(n_1193) );
BUFx2_ASAP7_75t_L g1353 ( .A(n_681), .Y(n_1353) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_700), .B(n_721), .Y(n_682) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_685), .A2(n_823), .B1(n_824), .B2(n_825), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_685), .A2(n_694), .B1(n_984), .B2(n_1008), .C(n_1013), .Y(n_1007) );
INVx3_ASAP7_75t_L g1165 ( .A(n_685), .Y(n_1165) );
AOI221xp5_ASAP7_75t_L g1215 ( .A1(n_685), .A2(n_694), .B1(n_1197), .B2(n_1216), .C(n_1217), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_686), .Y(n_693) );
BUFx2_ASAP7_75t_L g1131 ( .A(n_686), .Y(n_1131) );
INVx1_ASAP7_75t_L g1484 ( .A(n_686), .Y(n_1484) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_691), .B(n_694), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g812 ( .A1(n_694), .A2(n_813), .B1(n_814), .B2(n_815), .C(n_820), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_694), .A2(n_933), .B(n_937), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g1166 ( .A1(n_694), .A2(n_1167), .B(n_1168), .Y(n_1166) );
AOI21xp5_ASAP7_75t_L g1333 ( .A1(n_694), .A2(n_1334), .B(n_1335), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_697), .A2(n_699), .B1(n_930), .B2(n_931), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_697), .A2(n_823), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_697), .A2(n_699), .B1(n_1170), .B2(n_1171), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_697), .A2(n_699), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_697), .A2(n_823), .B1(n_1337), .B2(n_1338), .Y(n_1336) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_699), .Y(n_823) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g941 ( .A(n_702), .Y(n_941) );
INVx2_ASAP7_75t_L g1318 ( .A(n_702), .Y(n_1318) );
INVx4_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
BUFx3_ASAP7_75t_L g813 ( .A(n_704), .Y(n_813) );
BUFx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g1331 ( .A(n_707), .Y(n_1331) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g1825 ( .A(n_709), .Y(n_1825) );
OAI211xp5_ASAP7_75t_SL g710 ( .A1(n_711), .A2(n_712), .B(n_714), .C(n_718), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_712), .A2(n_1235), .B1(n_1236), .B2(n_1237), .Y(n_1234) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g1075 ( .A(n_713), .Y(n_1075) );
INVx1_ASAP7_75t_L g1771 ( .A(n_713), .Y(n_1771) );
INVx3_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g802 ( .A(n_716), .Y(n_802) );
INVx2_ASAP7_75t_L g946 ( .A(n_716), .Y(n_946) );
INVx1_ASAP7_75t_L g1017 ( .A(n_716), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g1154 ( .A1(n_716), .A2(n_944), .B1(n_1071), .B2(n_1155), .C(n_1156), .Y(n_1154) );
INVx1_ASAP7_75t_L g1434 ( .A(n_717), .Y(n_1434) );
INVxp67_ASAP7_75t_L g1453 ( .A(n_717), .Y(n_1453) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g1140 ( .A(n_720), .Y(n_1140) );
AOI21xp5_ASAP7_75t_L g1210 ( .A1(n_721), .A2(n_1211), .B(n_1222), .Y(n_1210) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI21xp33_ASAP7_75t_L g1092 ( .A1(n_722), .A2(n_1093), .B(n_1109), .Y(n_1092) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_SL g728 ( .A1(n_723), .A2(n_729), .B(n_752), .C(n_757), .Y(n_728) );
INVx1_ASAP7_75t_L g827 ( .A(n_723), .Y(n_827) );
BUFx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_724), .Y(n_950) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_761), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_737), .B(n_743), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_734), .A2(n_744), .B1(n_773), .B2(n_774), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B1(n_740), .B2(n_742), .Y(n_737) );
INVx1_ASAP7_75t_L g880 ( .A(n_738), .Y(n_880) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_742), .A2(n_769), .B1(n_776), .B2(n_778), .Y(n_775) );
OAI211xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_747), .C(n_750), .Y(n_743) );
INVx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g843 ( .A(n_746), .Y(n_843) );
INVx2_ASAP7_75t_L g1103 ( .A(n_746), .Y(n_1103) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_751), .Y(n_1041) );
INVx1_ASAP7_75t_L g1263 ( .A(n_751), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_782), .C(n_786), .Y(n_761) );
NOR2xp33_ASAP7_75t_SL g762 ( .A(n_763), .B(n_781), .Y(n_762) );
OAI33xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .A3(n_770), .B1(n_772), .B2(n_775), .B3(n_779), .Y(n_763) );
OAI33xp33_ASAP7_75t_L g1230 ( .A1(n_764), .A2(n_1231), .A3(n_1234), .B1(n_1238), .B2(n_1243), .B3(n_1248), .Y(n_1230) );
OAI22xp5_ASAP7_75t_SL g1304 ( .A1(n_764), .A2(n_1305), .B1(n_1307), .B2(n_1308), .Y(n_1304) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B1(n_768), .B2(n_769), .Y(n_765) );
OAI221xp5_ASAP7_75t_L g1308 ( .A1(n_774), .A2(n_1280), .B1(n_1285), .B2(n_1309), .C(n_1310), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1405 ( .A1(n_774), .A2(n_1134), .B1(n_1406), .B2(n_1407), .Y(n_1405) );
OAI22xp5_ASAP7_75t_L g1325 ( .A1(n_776), .A2(n_1326), .B1(n_1327), .B2(n_1330), .Y(n_1325) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g1248 ( .A(n_780), .Y(n_1248) );
AOI21xp5_ASAP7_75t_L g920 ( .A1(n_783), .A2(n_921), .B(n_922), .Y(n_920) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
XOR2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_867), .Y(n_788) );
XNOR2x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_857), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .B1(n_796), .B2(n_826), .C(n_828), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_812), .C(n_822), .Y(n_796) );
AOI222xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_803), .B1(n_806), .B2(n_808), .C1(n_809), .C2(n_811), .Y(n_797) );
BUFx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g935 ( .A(n_801), .Y(n_935) );
INVx1_ASAP7_75t_L g1324 ( .A(n_802), .Y(n_1324) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_805), .Y(n_821) );
INVx1_ASAP7_75t_L g1020 ( .A(n_806), .Y(n_1020) );
AOI222xp33_ASAP7_75t_L g1212 ( .A1(n_806), .A2(n_813), .B1(n_1208), .B2(n_1209), .C1(n_1213), .C2(n_1214), .Y(n_1212) );
AOI22xp33_ASAP7_75t_SL g1826 ( .A1(n_806), .A2(n_1827), .B1(n_1828), .B2(n_1829), .Y(n_1826) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AOI222xp33_ASAP7_75t_L g1014 ( .A1(n_813), .A2(n_988), .B1(n_989), .B2(n_1015), .C1(n_1018), .C2(n_1019), .Y(n_1014) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
HB1xp67_ASAP7_75t_SL g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_831), .B1(n_833), .B2(n_834), .Y(n_829) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_835), .Y(n_956) );
BUFx8_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
BUFx4f_ASAP7_75t_L g1419 ( .A(n_836), .Y(n_1419) );
BUFx2_ASAP7_75t_L g1794 ( .A(n_836), .Y(n_1794) );
OAI22xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_839), .B1(n_842), .B2(n_843), .Y(n_837) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g1856 ( .A1(n_841), .A2(n_876), .B1(n_1857), .B2(n_1858), .Y(n_1856) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
BUFx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_853), .Y(n_1000) );
BUFx2_ASAP7_75t_L g1192 ( .A(n_853), .Y(n_1192) );
INVx3_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx3_ASAP7_75t_L g967 ( .A(n_854), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_858), .B(n_1184), .Y(n_1183) );
INVx3_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx5_ASAP7_75t_L g1350 ( .A(n_859), .Y(n_1350) );
AOI22xp5_ASAP7_75t_L g1180 ( .A1(n_864), .A2(n_972), .B1(n_1181), .B2(n_1182), .Y(n_1180) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
NAND3xp33_ASAP7_75t_SL g986 ( .A(n_866), .B(n_987), .C(n_990), .Y(n_986) );
XNOR2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_923), .Y(n_867) );
OR2x2_ASAP7_75t_L g869 ( .A(n_870), .B(n_894), .Y(n_869) );
A2O1A1Ixp33_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_884), .B(n_888), .C(n_890), .Y(n_870) );
NOR3xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .C(n_879), .Y(n_871) );
INVx2_ASAP7_75t_L g1112 ( .A(n_876), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_883), .A2(n_906), .B1(n_907), .B2(n_909), .Y(n_905) );
A2O1A1Ixp33_ASAP7_75t_L g1256 ( .A1(n_888), .A2(n_1257), .B(n_1260), .C(n_1270), .Y(n_1256) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g1021 ( .A(n_889), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g1029 ( .A1(n_889), .A2(n_1030), .B(n_1055), .Y(n_1029) );
OAI21xp5_ASAP7_75t_L g1750 ( .A1(n_889), .A2(n_1751), .B(n_1778), .Y(n_1750) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
NAND4xp25_ASAP7_75t_L g894 ( .A(n_895), .B(n_898), .C(n_918), .D(n_920), .Y(n_894) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx4_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx3_ASAP7_75t_L g1067 ( .A(n_908), .Y(n_1067) );
BUFx6f_ASAP7_75t_L g1160 ( .A(n_908), .Y(n_1160) );
O2A1O1Ixp33_ASAP7_75t_L g1754 ( .A1(n_911), .A2(n_1438), .B(n_1755), .C(n_1756), .Y(n_1754) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_914), .B1(n_916), .B2(n_917), .Y(n_912) );
INVx1_ASAP7_75t_L g1403 ( .A(n_914), .Y(n_1403) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_917), .A2(n_1244), .B1(n_1246), .B2(n_1247), .Y(n_1243) );
NOR3xp33_ASAP7_75t_L g1303 ( .A(n_922), .B(n_1304), .C(n_1311), .Y(n_1303) );
AND4x1_ASAP7_75t_L g924 ( .A(n_925), .B(n_951), .C(n_973), .D(n_976), .Y(n_924) );
OAI21xp33_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_940), .B(n_950), .Y(n_925) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
OAI211xp5_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_944), .B(n_945), .C(n_947), .Y(n_942) );
OAI211xp5_ASAP7_75t_SL g1774 ( .A1(n_944), .A2(n_1775), .B(n_1776), .C(n_1777), .Y(n_1774) );
A2O1A1Ixp33_ASAP7_75t_L g1276 ( .A1(n_950), .A2(n_1277), .B(n_1291), .C(n_1298), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_957), .B1(n_960), .B2(n_966), .Y(n_952) );
OAI21xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B(n_956), .Y(n_953) );
INVx1_ASAP7_75t_L g1190 ( .A(n_954), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_961), .A2(n_1116), .B1(n_1117), .B2(n_1118), .Y(n_1115) );
OAI221xp5_ASAP7_75t_L g1800 ( .A1(n_961), .A2(n_1769), .B1(n_1775), .B2(n_1801), .C(n_1802), .Y(n_1800) );
CKINVDCx8_ASAP7_75t_R g961 ( .A(n_962), .Y(n_961) );
INVx3_ASAP7_75t_L g1269 ( .A(n_962), .Y(n_1269) );
INVx3_ASAP7_75t_L g1289 ( .A(n_962), .Y(n_1289) );
INVx3_ASAP7_75t_L g1425 ( .A(n_962), .Y(n_1425) );
OAI22xp5_ASAP7_75t_L g1793 ( .A1(n_966), .A2(n_1794), .B1(n_1795), .B2(n_1800), .Y(n_1793) );
CKINVDCx5p33_ASAP7_75t_R g966 ( .A(n_967), .Y(n_966) );
INVx2_ASAP7_75t_L g1427 ( .A(n_967), .Y(n_1427) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_977), .A2(n_1170), .B1(n_1171), .B2(n_1174), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_977), .A2(n_1174), .B1(n_1220), .B2(n_1221), .Y(n_1223) );
XNOR2xp5_ASAP7_75t_L g979 ( .A(n_980), .B(n_1025), .Y(n_979) );
XNOR2x1_ASAP7_75t_L g1313 ( .A(n_980), .B(n_1025), .Y(n_1313) );
BUFx3_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_983), .B(n_1002), .Y(n_982) );
AOI33xp33_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_992), .A3(n_996), .B1(n_998), .B2(n_1000), .B3(n_1001), .Y(n_990) );
AOI33xp33_ASAP7_75t_L g1351 ( .A1(n_991), .A2(n_1000), .A3(n_1352), .B1(n_1354), .B2(n_1355), .B3(n_1357), .Y(n_1351) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
AOI21xp5_ASAP7_75t_SL g1002 ( .A1(n_1003), .A2(n_1021), .B(n_1022), .Y(n_1002) );
NAND3xp33_ASAP7_75t_SL g1003 ( .A(n_1004), .B(n_1007), .C(n_1014), .Y(n_1003) );
INVx2_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1487 ( .A(n_1012), .Y(n_1487) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
O2A1O1Ixp33_ASAP7_75t_SL g1152 ( .A1(n_1021), .A2(n_1153), .B(n_1164), .C(n_1172), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1836 ( .A(n_1024), .B(n_1837), .Y(n_1836) );
XNOR2x1_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1147), .Y(n_1025) );
XNOR2x2_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1083), .Y(n_1026) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1081), .B(n_1082), .Y(n_1027) );
AND3x1_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1056), .C(n_1062), .Y(n_1028) );
AOI31xp33_ASAP7_75t_L g1082 ( .A1(n_1029), .A2(n_1056), .A3(n_1062), .B(n_1081), .Y(n_1082) );
NAND3xp33_ASAP7_75t_SL g1030 ( .A(n_1031), .B(n_1042), .C(n_1046), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1031 ( .A1(n_1032), .A2(n_1035), .B1(n_1036), .B2(n_1039), .Y(n_1031) );
INVx2_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
NOR3xp33_ASAP7_75t_L g1260 ( .A(n_1045), .B(n_1261), .C(n_1266), .Y(n_1260) );
NOR3xp33_ASAP7_75t_L g1277 ( .A(n_1045), .B(n_1278), .C(n_1283), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1490 ( .A(n_1045), .B(n_1491), .Y(n_1490) );
INVxp67_ASAP7_75t_L g1094 ( .A(n_1047), .Y(n_1094) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g1287 ( .A1(n_1050), .A2(n_1288), .B1(n_1289), .B2(n_1290), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1059), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1061), .Y(n_1059) );
OAI221xp5_ASAP7_75t_L g1070 ( .A1(n_1071), .A2(n_1074), .B1(n_1075), .B2(n_1076), .C(n_1077), .Y(n_1070) );
INVx3_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
OAI221xp5_ASAP7_75t_L g1305 ( .A1(n_1073), .A2(n_1129), .B1(n_1281), .B2(n_1288), .C(n_1306), .Y(n_1305) );
OAI33xp33_ASAP7_75t_L g1399 ( .A1(n_1078), .A2(n_1400), .A3(n_1405), .B1(n_1408), .B2(n_1411), .B3(n_1413), .Y(n_1399) );
BUFx6f_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NAND3xp33_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1092), .C(n_1119), .Y(n_1085) );
OAI211xp5_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1095), .B(n_1097), .C(n_1100), .Y(n_1093) );
OAI211xp5_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1102), .B(n_1104), .C(n_1107), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g1133 ( .A1(n_1101), .A2(n_1113), .B1(n_1134), .B2(n_1137), .C(n_1138), .Y(n_1133) );
HB1xp67_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
OAI22xp5_ASAP7_75t_L g1268 ( .A1(n_1106), .A2(n_1235), .B1(n_1247), .B2(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
OAI221xp5_ASAP7_75t_L g1125 ( .A1(n_1117), .A2(n_1126), .B1(n_1128), .B2(n_1129), .C(n_1130), .Y(n_1125) );
NOR3xp33_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1132), .C(n_1142), .Y(n_1119) );
INVxp67_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx2_ASAP7_75t_SL g1123 ( .A(n_1124), .Y(n_1123) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
BUFx2_ASAP7_75t_L g1240 ( .A(n_1127), .Y(n_1240) );
INVx2_ASAP7_75t_L g1309 ( .A(n_1127), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_1134), .A2(n_1320), .B1(n_1409), .B2(n_1410), .Y(n_1408) );
INVx2_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
INVx4_ASAP7_75t_L g1236 ( .A(n_1135), .Y(n_1236) );
INVx2_ASAP7_75t_L g1817 ( .A(n_1135), .Y(n_1817) );
INVx4_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1140), .Y(n_1218) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
XNOR2xp5_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1224), .Y(n_1147) );
XNOR2xp5_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1194), .Y(n_1148) );
NOR2x1p5_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1176), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1159), .B1(n_1161), .B2(n_1162), .Y(n_1157) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx2_ASAP7_75t_SL g1414 ( .A(n_1160), .Y(n_1414) );
OAI22xp5_ASAP7_75t_L g1413 ( .A1(n_1162), .A2(n_1414), .B1(n_1415), .B2(n_1416), .Y(n_1413) );
BUFx3_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1838 ( .A1(n_1174), .A2(n_1829), .B1(n_1839), .B2(n_1840), .Y(n_1838) );
INVx2_ASAP7_75t_L g1265 ( .A(n_1175), .Y(n_1265) );
INVx2_ASAP7_75t_L g1294 ( .A(n_1175), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1179), .Y(n_1176) );
AND4x1_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1183), .C(n_1185), .D(n_1193), .Y(n_1179) );
NAND3xp33_ASAP7_75t_L g1199 ( .A(n_1193), .B(n_1200), .C(n_1207), .Y(n_1199) );
AND4x1_ASAP7_75t_SL g1343 ( .A(n_1193), .B(n_1344), .C(n_1348), .D(n_1351), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1210), .Y(n_1195) );
NAND3xp33_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1215), .C(n_1219), .Y(n_1211) );
XNOR2x1_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1272), .Y(n_1224) );
XNOR2x1_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1227), .Y(n_1225) );
NOR2x1_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1256), .Y(n_1227) );
NAND3xp33_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1250), .C(n_1254), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1249), .Y(n_1229) );
INVx4_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
OAI22xp5_ASAP7_75t_L g1853 ( .A1(n_1265), .A2(n_1851), .B1(n_1854), .B2(n_1855), .Y(n_1853) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
XNOR2x1_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1275), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1299), .Y(n_1275) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1307), .Y(n_1412) );
OAI221xp5_ASAP7_75t_L g1319 ( .A1(n_1309), .A2(n_1320), .B1(n_1322), .B2(n_1323), .C(n_1324), .Y(n_1319) );
INVx2_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1314), .Y(n_1358) );
NAND3x1_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1341), .C(n_1343), .Y(n_1315) );
INVx5_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
BUFx2_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
BUFx6f_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1349), .B(n_1350), .Y(n_1348) );
AOI22xp5_ASAP7_75t_L g1359 ( .A1(n_1360), .A2(n_1361), .B1(n_1462), .B2(n_1507), .Y(n_1359) );
INVx2_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1362), .Y(n_1460) );
OAI211xp5_ASAP7_75t_L g1362 ( .A1(n_1363), .A2(n_1369), .B(n_1398), .C(n_1429), .Y(n_1362) );
CKINVDCx14_ASAP7_75t_R g1363 ( .A(n_1364), .Y(n_1363) );
AND2x4_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1367), .Y(n_1364) );
AND2x2_ASAP7_75t_SL g1792 ( .A(n_1365), .B(n_1367), .Y(n_1792) );
INVx1_ASAP7_75t_SL g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
NOR3xp33_ASAP7_75t_SL g1369 ( .A(n_1370), .B(n_1377), .C(n_1392), .Y(n_1369) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx2_ASAP7_75t_SL g1372 ( .A(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1373), .Y(n_1789) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
CKINVDCx8_ASAP7_75t_R g1380 ( .A(n_1381), .Y(n_1380) );
NOR3xp33_ASAP7_75t_L g1780 ( .A(n_1381), .B(n_1781), .C(n_1787), .Y(n_1780) );
AOI22xp33_ASAP7_75t_L g1382 ( .A1(n_1383), .A2(n_1387), .B1(n_1388), .B2(n_1391), .Y(n_1382) );
BUFx3_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1385), .B(n_1386), .Y(n_1384) );
AND2x4_ASAP7_75t_L g1389 ( .A(n_1385), .B(n_1390), .Y(n_1389) );
AND2x4_ASAP7_75t_L g1784 ( .A(n_1385), .B(n_1386), .Y(n_1784) );
AND2x2_ASAP7_75t_L g1786 ( .A(n_1385), .B(n_1390), .Y(n_1786) );
AOI22xp33_ASAP7_75t_L g1435 ( .A1(n_1387), .A2(n_1436), .B1(n_1439), .B2(n_1440), .Y(n_1435) );
BUFx6f_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
BUFx2_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
INVx2_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
NOR2xp33_ASAP7_75t_L g1398 ( .A(n_1399), .B(n_1417), .Y(n_1398) );
OAI22xp33_ASAP7_75t_L g1420 ( .A1(n_1401), .A2(n_1409), .B1(n_1421), .B2(n_1423), .Y(n_1420) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
INVx2_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
OAI33xp33_ASAP7_75t_L g1417 ( .A1(n_1418), .A2(n_1420), .A3(n_1424), .B1(n_1426), .B2(n_1427), .B3(n_1428), .Y(n_1417) );
BUFx3_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
OAI33xp33_ASAP7_75t_L g1845 ( .A1(n_1419), .A2(n_1846), .A3(n_1849), .B1(n_1853), .B2(n_1856), .B3(n_1859), .Y(n_1845) );
INVx2_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
OAI31xp33_ASAP7_75t_L g1429 ( .A1(n_1430), .A2(n_1443), .A3(n_1451), .B(n_1456), .Y(n_1429) );
INVx3_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
BUFx3_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1438), .Y(n_1761) );
INVx2_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
INVx2_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
HB1xp67_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
BUFx2_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1450), .Y(n_1764) );
INVx3_ASAP7_75t_L g1519 ( .A(n_1452), .Y(n_1519) );
AOI22xp5_ASAP7_75t_L g1759 ( .A1(n_1453), .A2(n_1760), .B1(n_1761), .B2(n_1762), .Y(n_1759) );
CKINVDCx16_ASAP7_75t_R g1454 ( .A(n_1455), .Y(n_1454) );
INVx3_ASAP7_75t_SL g1753 ( .A(n_1455), .Y(n_1753) );
BUFx3_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
AND2x4_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1459), .Y(n_1457) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1458), .Y(n_1518) );
AOI21xp5_ASAP7_75t_SL g1751 ( .A1(n_1458), .A2(n_1752), .B(n_1766), .Y(n_1751) );
NOR2xp33_ASAP7_75t_L g1807 ( .A(n_1458), .B(n_1510), .Y(n_1807) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1462), .Y(n_1507) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
OAI21x1_ASAP7_75t_SL g1463 ( .A1(n_1464), .A2(n_1465), .B(n_1506), .Y(n_1463) );
NAND4xp25_ASAP7_75t_L g1506 ( .A(n_1464), .B(n_1467), .C(n_1469), .D(n_1488), .Y(n_1506) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
NAND3xp33_ASAP7_75t_L g1466 ( .A(n_1467), .B(n_1469), .C(n_1488), .Y(n_1466) );
NOR2xp33_ASAP7_75t_L g1469 ( .A(n_1470), .B(n_1474), .Y(n_1469) );
NAND3xp33_ASAP7_75t_SL g1474 ( .A(n_1475), .B(n_1478), .C(n_1481), .Y(n_1474) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
NAND3xp33_ASAP7_75t_L g1489 ( .A(n_1490), .B(n_1494), .C(n_1499), .Y(n_1489) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_1495), .A2(n_1496), .B1(n_1497), .B2(n_1498), .Y(n_1494) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
INVx2_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
OR2x2_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1516), .Y(n_1509) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
NOR2xp33_ASAP7_75t_L g1511 ( .A(n_1512), .B(n_1514), .Y(n_1511) );
NOR2xp33_ASAP7_75t_L g1863 ( .A(n_1512), .B(n_1515), .Y(n_1863) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1512), .Y(n_1867) );
HB1xp67_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
NOR2xp33_ASAP7_75t_L g1870 ( .A(n_1515), .B(n_1867), .Y(n_1870) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1519), .Y(n_1517) );
AND2x4_ASAP7_75t_SL g1806 ( .A(n_1519), .B(n_1807), .Y(n_1806) );
OAI221xp5_ASAP7_75t_L g1520 ( .A1(n_1521), .A2(n_1746), .B1(n_1748), .B2(n_1803), .C(n_1808), .Y(n_1520) );
NOR5xp2_ASAP7_75t_L g1521 ( .A(n_1522), .B(n_1661), .C(n_1723), .D(n_1729), .E(n_1740), .Y(n_1521) );
AOI31xp33_ASAP7_75t_L g1522 ( .A1(n_1523), .A2(n_1605), .A3(n_1635), .B(n_1655), .Y(n_1522) );
AOI211xp5_ASAP7_75t_SL g1523 ( .A1(n_1524), .A2(n_1540), .B(n_1559), .C(n_1573), .Y(n_1523) );
A2O1A1Ixp33_ASAP7_75t_L g1662 ( .A1(n_1524), .A2(n_1663), .B(n_1665), .C(n_1677), .Y(n_1662) );
CKINVDCx6p67_ASAP7_75t_R g1524 ( .A(n_1525), .Y(n_1524) );
CKINVDCx6p67_ASAP7_75t_R g1525 ( .A(n_1526), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1526), .B(n_1601), .Y(n_1603) );
INVx2_ASAP7_75t_L g1613 ( .A(n_1526), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_1526), .B(n_1673), .Y(n_1672) );
OAI22xp5_ASAP7_75t_L g1683 ( .A1(n_1526), .A2(n_1684), .B1(n_1686), .B2(n_1688), .Y(n_1683) );
AND2x4_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1534), .Y(n_1526) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1527), .B(n_1534), .Y(n_1565) );
AND2x6_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1530), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1529), .B(n_1533), .Y(n_1532) );
AND2x4_ASAP7_75t_L g1535 ( .A(n_1529), .B(n_1536), .Y(n_1535) );
AND2x6_ASAP7_75t_L g1538 ( .A(n_1529), .B(n_1539), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1529), .B(n_1533), .Y(n_1546) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1529), .B(n_1533), .Y(n_1550) );
NAND2xp5_ASAP7_75t_L g1747 ( .A(n_1529), .B(n_1536), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1531), .B(n_1537), .Y(n_1536) );
HB1xp67_ASAP7_75t_L g1868 ( .A(n_1536), .Y(n_1868) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1547), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1542), .B(n_1588), .Y(n_1587) );
NAND2xp5_ASAP7_75t_SL g1609 ( .A(n_1542), .B(n_1610), .Y(n_1609) );
OR2x2_ASAP7_75t_L g1688 ( .A(n_1542), .B(n_1689), .Y(n_1688) );
INVx2_ASAP7_75t_L g1692 ( .A(n_1542), .Y(n_1692) );
INVx2_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
INVx3_ASAP7_75t_L g1567 ( .A(n_1543), .Y(n_1567) );
NOR2xp33_ASAP7_75t_L g1585 ( .A(n_1543), .B(n_1548), .Y(n_1585) );
NAND2xp5_ASAP7_75t_L g1617 ( .A(n_1543), .B(n_1618), .Y(n_1617) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1543), .B(n_1548), .Y(n_1640) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1543), .B(n_1582), .Y(n_1644) );
NAND2xp5_ASAP7_75t_L g1674 ( .A(n_1543), .B(n_1631), .Y(n_1674) );
NOR2xp33_ASAP7_75t_L g1682 ( .A(n_1543), .B(n_1593), .Y(n_1682) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1545), .Y(n_1543) );
NAND2xp5_ASAP7_75t_L g1727 ( .A(n_1547), .B(n_1577), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1552), .Y(n_1547) );
CKINVDCx5p33_ASAP7_75t_R g1608 ( .A(n_1548), .Y(n_1608) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1548), .B(n_1620), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1548), .B(n_1571), .Y(n_1697) );
OR2x2_ASAP7_75t_L g1709 ( .A(n_1548), .B(n_1584), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1712 ( .A(n_1548), .B(n_1645), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1551), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1549), .B(n_1551), .Y(n_1569) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1552), .Y(n_1593) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1552), .B(n_1640), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1670 ( .A(n_1552), .B(n_1608), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1556), .Y(n_1552) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1553), .Y(n_1572) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1553), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1555), .Y(n_1553) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1556), .Y(n_1571) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1556), .Y(n_1584) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1556), .B(n_1572), .Y(n_1597) );
OR2x2_ASAP7_75t_L g1611 ( .A(n_1556), .B(n_1572), .Y(n_1611) );
NAND2xp5_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1558), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1566), .Y(n_1559) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
OR2x2_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1565), .Y(n_1561) );
INVx3_ASAP7_75t_L g1582 ( .A(n_1562), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1562), .B(n_1599), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1562), .B(n_1613), .Y(n_1612) );
OR2x2_ASAP7_75t_L g1615 ( .A(n_1562), .B(n_1600), .Y(n_1615) );
NOR2xp33_ASAP7_75t_L g1623 ( .A(n_1562), .B(n_1576), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1637 ( .A(n_1562), .B(n_1565), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1651 ( .A(n_1562), .B(n_1576), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1562), .B(n_1627), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1562), .B(n_1631), .Y(n_1687) );
AND2x2_ASAP7_75t_L g1695 ( .A(n_1562), .B(n_1677), .Y(n_1695) );
INVx3_ASAP7_75t_L g1739 ( .A(n_1562), .Y(n_1739) );
AND2x4_ASAP7_75t_SL g1562 ( .A(n_1563), .B(n_1564), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1565), .B(n_1582), .Y(n_1581) );
OR2x2_ASAP7_75t_L g1589 ( .A(n_1565), .B(n_1578), .Y(n_1589) );
OR2x2_ASAP7_75t_L g1600 ( .A(n_1565), .B(n_1601), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1565), .B(n_1578), .Y(n_1627) );
NOR2xp33_ASAP7_75t_L g1710 ( .A(n_1565), .B(n_1658), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1568), .Y(n_1566) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1567), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1664 ( .A(n_1567), .B(n_1597), .Y(n_1664) );
NOR2xp33_ASAP7_75t_L g1667 ( .A(n_1567), .B(n_1611), .Y(n_1667) );
O2A1O1Ixp33_ASAP7_75t_L g1669 ( .A1(n_1567), .A2(n_1627), .B(n_1670), .C(n_1671), .Y(n_1669) );
NAND2xp5_ASAP7_75t_L g1699 ( .A(n_1567), .B(n_1601), .Y(n_1699) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1567), .B(n_1703), .Y(n_1702) );
NOR2xp33_ASAP7_75t_L g1708 ( .A(n_1567), .B(n_1709), .Y(n_1708) );
NOR2xp33_ASAP7_75t_L g1711 ( .A(n_1567), .B(n_1712), .Y(n_1711) );
NAND3xp33_ASAP7_75t_L g1715 ( .A(n_1567), .B(n_1677), .C(n_1716), .Y(n_1715) );
NAND2xp5_ASAP7_75t_L g1732 ( .A(n_1567), .B(n_1599), .Y(n_1732) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1568), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1568 ( .A(n_1569), .B(n_1570), .Y(n_1568) );
AOI32xp33_ASAP7_75t_L g1586 ( .A1(n_1569), .A2(n_1587), .A3(n_1590), .B1(n_1594), .B2(n_1598), .Y(n_1586) );
OR2x2_ASAP7_75t_L g1595 ( .A(n_1569), .B(n_1596), .Y(n_1595) );
OR2x2_ASAP7_75t_L g1633 ( .A(n_1569), .B(n_1634), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1569), .B(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1570), .Y(n_1592) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1570), .B(n_1608), .Y(n_1647) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1570), .B(n_1585), .Y(n_1649) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1570), .B(n_1654), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1572), .Y(n_1570) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1572), .Y(n_1620) );
OAI211xp5_ASAP7_75t_L g1573 ( .A1(n_1574), .A2(n_1583), .B(n_1586), .C(n_1602), .Y(n_1573) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1581), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1576), .B(n_1639), .Y(n_1685) );
O2A1O1Ixp33_ASAP7_75t_L g1733 ( .A1(n_1576), .A2(n_1664), .B(n_1670), .C(n_1734), .Y(n_1733) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1576), .Y(n_1736) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1577), .B(n_1639), .Y(n_1638) );
AOI322xp5_ASAP7_75t_L g1707 ( .A1(n_1577), .A2(n_1623), .A3(n_1649), .B1(n_1695), .B2(n_1708), .C1(n_1710), .C2(n_1711), .Y(n_1707) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1578), .Y(n_1601) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1578), .Y(n_1631) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1580), .Y(n_1578) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1581), .Y(n_1728) );
NAND2xp5_ASAP7_75t_L g1706 ( .A(n_1582), .B(n_1588), .Y(n_1706) );
OR2x2_ASAP7_75t_L g1718 ( .A(n_1582), .B(n_1589), .Y(n_1718) );
AOI32xp33_ASAP7_75t_L g1742 ( .A1(n_1582), .A2(n_1587), .A3(n_1676), .B1(n_1677), .B2(n_1743), .Y(n_1742) );
NAND2xp5_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1585), .Y(n_1583) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1584), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1585), .B(n_1597), .Y(n_1604) );
AOI311xp33_ASAP7_75t_L g1690 ( .A1(n_1588), .A2(n_1691), .A3(n_1692), .B(n_1693), .C(n_1704), .Y(n_1690) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
OAI321xp33_ASAP7_75t_L g1641 ( .A1(n_1589), .A2(n_1642), .A3(n_1643), .B1(n_1645), .B2(n_1646), .C(n_1648), .Y(n_1641) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
NAND2xp5_ASAP7_75t_L g1591 ( .A(n_1592), .B(n_1593), .Y(n_1591) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
OR2x2_ASAP7_75t_L g1745 ( .A(n_1596), .B(n_1608), .Y(n_1745) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1634 ( .A(n_1597), .B(n_1626), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1597), .B(n_1640), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1599), .B(n_1626), .Y(n_1722) );
INVx2_ASAP7_75t_SL g1599 ( .A(n_1600), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1602 ( .A(n_1603), .B(n_1604), .Y(n_1602) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1603), .Y(n_1642) );
AOI221xp5_ASAP7_75t_L g1605 ( .A1(n_1606), .A2(n_1612), .B1(n_1614), .B2(n_1616), .C(n_1621), .Y(n_1605) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
OR2x2_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1609), .Y(n_1607) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1608), .B(n_1645), .Y(n_1676) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1608), .B(n_1667), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1608), .B(n_1620), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1705 ( .A(n_1610), .B(n_1640), .Y(n_1705) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1612), .Y(n_1668) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
INVxp67_ASAP7_75t_SL g1616 ( .A(n_1617), .Y(n_1616) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
A2O1A1Ixp33_ASAP7_75t_L g1621 ( .A1(n_1622), .A2(n_1624), .B(n_1628), .C(n_1629), .Y(n_1621) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1623), .Y(n_1622) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1626), .B(n_1627), .Y(n_1625) );
CKINVDCx14_ASAP7_75t_R g1741 ( .A(n_1627), .Y(n_1741) );
NAND2xp5_ASAP7_75t_L g1691 ( .A(n_1628), .B(n_1689), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1632), .Y(n_1629) );
NAND2xp5_ASAP7_75t_L g1724 ( .A(n_1630), .B(n_1725), .Y(n_1724) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
NAND2xp5_ASAP7_75t_L g1680 ( .A(n_1633), .B(n_1681), .Y(n_1680) );
AOI211xp5_ASAP7_75t_L g1635 ( .A1(n_1636), .A2(n_1638), .B(n_1641), .C(n_1652), .Y(n_1635) );
NAND3xp33_ASAP7_75t_L g1700 ( .A(n_1636), .B(n_1657), .C(n_1701), .Y(n_1700) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
A2O1A1Ixp33_ASAP7_75t_L g1693 ( .A1(n_1637), .A2(n_1694), .B(n_1696), .C(n_1700), .Y(n_1693) );
NOR2xp33_ASAP7_75t_L g1671 ( .A(n_1642), .B(n_1646), .Y(n_1671) );
OAI221xp5_ASAP7_75t_SL g1704 ( .A1(n_1642), .A2(n_1646), .B1(n_1705), .B2(n_1706), .C(n_1707), .Y(n_1704) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1645), .Y(n_1716) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
OAI21xp5_ASAP7_75t_L g1648 ( .A1(n_1649), .A2(n_1650), .B(n_1651), .Y(n_1648) );
NAND2xp5_ASAP7_75t_L g1735 ( .A(n_1650), .B(n_1736), .Y(n_1735) );
AOI221xp5_ASAP7_75t_L g1678 ( .A1(n_1651), .A2(n_1654), .B1(n_1679), .B2(n_1680), .C(n_1683), .Y(n_1678) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1651), .Y(n_1744) );
INVxp67_ASAP7_75t_SL g1652 ( .A(n_1653), .Y(n_1652) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
AND2x2_ASAP7_75t_L g1738 ( .A(n_1657), .B(n_1739), .Y(n_1738) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1658), .Y(n_1657) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1658), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_1659), .B(n_1660), .Y(n_1658) );
NAND4xp25_ASAP7_75t_L g1661 ( .A(n_1662), .B(n_1678), .C(n_1690), .D(n_1713), .Y(n_1661) );
CKINVDCx14_ASAP7_75t_R g1726 ( .A(n_1663), .Y(n_1726) );
OAI211xp5_ASAP7_75t_SL g1665 ( .A1(n_1666), .A2(n_1668), .B(n_1669), .C(n_1672), .Y(n_1665) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1670), .Y(n_1689) );
O2A1O1Ixp33_ASAP7_75t_L g1713 ( .A1(n_1670), .A2(n_1714), .B(n_1717), .C(n_1719), .Y(n_1713) );
NOR2xp33_ASAP7_75t_L g1673 ( .A(n_1674), .B(n_1675), .Y(n_1673) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1688), .Y(n_1725) );
O2A1O1Ixp33_ASAP7_75t_L g1719 ( .A1(n_1694), .A2(n_1705), .B(n_1720), .C(n_1721), .Y(n_1719) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
NAND2xp5_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1698), .Y(n_1696) );
O2A1O1Ixp33_ASAP7_75t_L g1729 ( .A1(n_1697), .A2(n_1730), .B(n_1733), .C(n_1737), .Y(n_1729) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
INVxp67_ASAP7_75t_SL g1714 ( .A(n_1715), .Y(n_1714) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
A2O1A1Ixp33_ASAP7_75t_L g1740 ( .A1(n_1718), .A2(n_1726), .B(n_1741), .C(n_1742), .Y(n_1740) );
INVxp67_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
AOI31xp33_ASAP7_75t_L g1723 ( .A1(n_1724), .A2(n_1726), .A3(n_1727), .B(n_1728), .Y(n_1723) );
INVxp67_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1732), .Y(n_1731) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
NOR2xp33_ASAP7_75t_L g1743 ( .A(n_1744), .B(n_1745), .Y(n_1743) );
BUFx2_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
HB1xp67_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
AOI22xp33_ASAP7_75t_SL g1788 ( .A1(n_1760), .A2(n_1789), .B1(n_1790), .B2(n_1791), .Y(n_1788) );
NAND2xp5_ASAP7_75t_SL g1763 ( .A(n_1764), .B(n_1765), .Y(n_1763) );
OAI21xp5_ASAP7_75t_L g1766 ( .A1(n_1767), .A2(n_1770), .B(n_1774), .Y(n_1766) );
AOI21xp5_ASAP7_75t_L g1778 ( .A1(n_1779), .A2(n_1792), .B(n_1793), .Y(n_1778) );
NAND2xp5_ASAP7_75t_SL g1779 ( .A(n_1780), .B(n_1788), .Y(n_1779) );
INVx1_ASAP7_75t_L g1783 ( .A(n_1784), .Y(n_1783) );
INVxp67_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
OAI211xp5_ASAP7_75t_L g1795 ( .A1(n_1796), .A2(n_1797), .B(n_1798), .C(n_1799), .Y(n_1795) );
CKINVDCx20_ASAP7_75t_R g1803 ( .A(n_1804), .Y(n_1803) );
CKINVDCx20_ASAP7_75t_R g1804 ( .A(n_1805), .Y(n_1804) );
INVx3_ASAP7_75t_L g1805 ( .A(n_1806), .Y(n_1805) );
INVxp33_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
HB1xp67_ASAP7_75t_L g1811 ( .A(n_1812), .Y(n_1811) );
INVx2_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
OR2x2_ASAP7_75t_L g1813 ( .A(n_1814), .B(n_1835), .Y(n_1813) );
AOI21xp5_ASAP7_75t_L g1815 ( .A1(n_1816), .A2(n_1821), .B(n_1822), .Y(n_1815) );
NAND2xp5_ASAP7_75t_L g1822 ( .A(n_1823), .B(n_1826), .Y(n_1822) );
AOI22xp5_ASAP7_75t_L g1830 ( .A1(n_1831), .A2(n_1832), .B1(n_1833), .B2(n_1834), .Y(n_1830) );
NAND3xp33_ASAP7_75t_SL g1835 ( .A(n_1836), .B(n_1838), .C(n_1841), .Y(n_1835) );
NOR2xp33_ASAP7_75t_SL g1841 ( .A(n_1842), .B(n_1845), .Y(n_1841) );
HB1xp67_ASAP7_75t_L g1860 ( .A(n_1861), .Y(n_1860) );
BUFx3_ASAP7_75t_L g1861 ( .A(n_1862), .Y(n_1861) );
BUFx3_ASAP7_75t_L g1862 ( .A(n_1863), .Y(n_1862) );
HB1xp67_ASAP7_75t_L g1864 ( .A(n_1865), .Y(n_1864) );
HB1xp67_ASAP7_75t_L g1865 ( .A(n_1866), .Y(n_1865) );
OAI21xp5_ASAP7_75t_L g1866 ( .A1(n_1867), .A2(n_1868), .B(n_1869), .Y(n_1866) );
INVx1_ASAP7_75t_L g1869 ( .A(n_1870), .Y(n_1869) );
endmodule