module fake_jpeg_25566_n_103 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_103);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_103;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_52),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_0),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_51),
.A2(n_35),
.B1(n_44),
.B2(n_41),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_42),
.B1(n_45),
.B2(n_3),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_35),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_39),
.C(n_43),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_7),
.C(n_8),
.Y(n_77)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_0),
.CON(n_64),
.SN(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_75)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_1),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_14),
.B(n_31),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_13),
.B(n_15),
.C(n_17),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_2),
.B(n_3),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_2),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_4),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_75),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_5),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_9),
.B1(n_57),
.B2(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_72),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_20),
.B1(n_10),
.B2(n_11),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_71),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_85),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_19),
.B1(n_21),
.B2(n_24),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_77),
.B(n_30),
.C(n_34),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_91),
.B(n_85),
.Y(n_95)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_90),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_75),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_84),
.C(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_95),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_82),
.Y(n_97)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_81),
.CI(n_89),
.CON(n_98),
.SN(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_96),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_98),
.B(n_87),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_78),
.C(n_98),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_87),
.C(n_27),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_57),
.Y(n_103)
);


endmodule