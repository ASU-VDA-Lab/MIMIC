module fake_ariane_1515_n_1957 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1957);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1957;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_204),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_81),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_147),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_136),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_80),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_50),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_24),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_29),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_162),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_54),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_9),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_12),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_39),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_38),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_66),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_5),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_4),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_44),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_194),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_11),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_137),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_64),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_96),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_112),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_58),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_173),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_161),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_97),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_50),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_201),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_123),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_171),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_0),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_179),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_2),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_89),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_156),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_14),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_86),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_26),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_55),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_159),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_88),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_67),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_183),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_178),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_111),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_207),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_21),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_148),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_37),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_73),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_110),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_27),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_141),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_16),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_119),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_195),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_151),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_76),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_106),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_193),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_37),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_69),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_71),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_48),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_19),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_167),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_90),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_116),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_76),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_113),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_94),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_160),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_73),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_144),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_2),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_185),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_69),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_79),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_63),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_189),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_127),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_181),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_99),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_64),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_129),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_77),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_70),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_191),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_21),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_142),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_4),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_150),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_24),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_135),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_29),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_27),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_176),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_188),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_205),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_153),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_203),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_107),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_43),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_199),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_84),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_169),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_100),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_6),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_7),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_154),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_139),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_68),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_36),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_43),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_71),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_140),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_126),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_28),
.Y(n_336)
);

BUFx8_ASAP7_75t_SL g337 ( 
.A(n_33),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_30),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_133),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_18),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_3),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_172),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_91),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_164),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_62),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_83),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_47),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_33),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_102),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_145),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_18),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_163),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_197),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_124),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_186),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_128),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_59),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_52),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_53),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_157),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_47),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_58),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_168),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_11),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_70),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_166),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_39),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_118),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_40),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_1),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_42),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_12),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_132),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_57),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_62),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_59),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_60),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_65),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_105),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_45),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_152),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_114),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_35),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_66),
.Y(n_384)
);

BUFx8_ASAP7_75t_SL g385 ( 
.A(n_35),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_15),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_22),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_146),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_54),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_28),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_7),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_158),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_75),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_36),
.Y(n_394)
);

INVxp33_ASAP7_75t_R g395 ( 
.A(n_32),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_5),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_52),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_120),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_0),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_31),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_174),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_25),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_55),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_15),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_8),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_93),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_53),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_104),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_63),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_14),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_403),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_1),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_337),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_R g414 ( 
.A(n_216),
.B(n_253),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_403),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_385),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_403),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_292),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_243),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_212),
.B(n_3),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_316),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_254),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_212),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_335),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_224),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_224),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_254),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_213),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_224),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_213),
.B(n_8),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_348),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_270),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_270),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_223),
.B(n_9),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_223),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_228),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_228),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_357),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_304),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_231),
.B(n_10),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_309),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_396),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_309),
.B(n_10),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_305),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_397),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_231),
.B(n_235),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_235),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_305),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_372),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_372),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_240),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_386),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_240),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_244),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_244),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_383),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_258),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_258),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_326),
.B(n_13),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_263),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_263),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_383),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_273),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_273),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_278),
.B(n_13),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_278),
.B(n_289),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_217),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_289),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_405),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_308),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_304),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_308),
.B(n_16),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_304),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_310),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_218),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_221),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_329),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_225),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_310),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_226),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_227),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_229),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_312),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_232),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_312),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_219),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_329),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_317),
.B(n_17),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_329),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_234),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_243),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_237),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_260),
.B(n_17),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_342),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_358),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_317),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_318),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_326),
.B(n_19),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_342),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_342),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_243),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_241),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_234),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_318),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_249),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_219),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_243),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_257),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_375),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_325),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_375),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_268),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_375),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_415),
.B(n_325),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_488),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_418),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_439),
.B(n_245),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_488),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_493),
.B(n_339),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_415),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_488),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_417),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_497),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_417),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_488),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_508),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_421),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_411),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_505),
.B(n_245),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_411),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_425),
.B(n_245),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_508),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_423),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_423),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_446),
.B(n_339),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_484),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_428),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_428),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_435),
.Y(n_542)
);

NOR2x1_ASAP7_75t_L g543 ( 
.A(n_439),
.B(n_322),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_432),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_435),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_436),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_437),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_437),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_467),
.B(n_350),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_447),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_426),
.B(n_380),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_447),
.B(n_209),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_451),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_451),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_453),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_453),
.B(n_454),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_495),
.B(n_336),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_454),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_455),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_455),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_457),
.B(n_209),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_457),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_458),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_458),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_461),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_495),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_461),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_462),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_462),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_464),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_464),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_465),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_465),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_486),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_469),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_469),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_471),
.B(n_350),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_471),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_476),
.B(n_360),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_476),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_481),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_481),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_485),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_485),
.Y(n_585)
);

AND2x2_ASAP7_75t_SL g586 ( 
.A(n_443),
.B(n_238),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_487),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_429),
.B(n_380),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_487),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_431),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_498),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_498),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_499),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_499),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_506),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_506),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_512),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_427),
.A2(n_378),
.B1(n_336),
.B2(n_276),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_512),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_537),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_521),
.B(n_468),
.Y(n_601)
);

INVx6_ASAP7_75t_L g602 ( 
.A(n_519),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_537),
.Y(n_603)
);

AND2x2_ASAP7_75t_SL g604 ( 
.A(n_586),
.B(n_443),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_537),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_586),
.B(n_477),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g607 ( 
.A(n_539),
.B(n_440),
.C(n_434),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_537),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_567),
.B(n_419),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_526),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_537),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_586),
.A2(n_558),
.B1(n_567),
.B2(n_550),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_537),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_537),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_567),
.B(n_478),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_568),
.Y(n_616)
);

INVxp33_ASAP7_75t_L g617 ( 
.A(n_526),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_540),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_540),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_540),
.Y(n_620)
);

AND2x2_ASAP7_75t_SL g621 ( 
.A(n_567),
.B(n_238),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_589),
.B(n_480),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_539),
.B(n_422),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_540),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_589),
.B(n_482),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_590),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_540),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_558),
.B(n_460),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_540),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_558),
.A2(n_420),
.B1(n_430),
.B2(n_452),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_589),
.B(n_483),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_540),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_558),
.A2(n_441),
.B1(n_459),
.B2(n_460),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_558),
.B(n_500),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_548),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_561),
.B(n_494),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_548),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_548),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_548),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_548),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_548),
.Y(n_641)
);

INVxp33_ASAP7_75t_SL g642 ( 
.A(n_518),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_575),
.B(n_504),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_548),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_532),
.Y(n_645)
);

AND2x2_ASAP7_75t_SL g646 ( 
.A(n_538),
.B(n_275),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_554),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_532),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_557),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_554),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_554),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_538),
.B(n_466),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_554),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_575),
.B(n_507),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_543),
.B(n_510),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_554),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_568),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_554),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_543),
.B(n_433),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_554),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_534),
.B(n_492),
.Y(n_661)
);

CKINVDCx11_ASAP7_75t_R g662 ( 
.A(n_558),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_598),
.B(n_444),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_561),
.B(n_473),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_522),
.B(n_360),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_560),
.Y(n_666)
);

NOR3xp33_ASAP7_75t_L g667 ( 
.A(n_550),
.B(n_490),
.C(n_474),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_530),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_560),
.Y(n_669)
);

INVxp67_ASAP7_75t_SL g670 ( 
.A(n_557),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_534),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_598),
.B(n_448),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_544),
.A2(n_500),
.B1(n_449),
.B2(n_456),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_560),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_519),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_552),
.B(n_450),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_560),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_560),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_560),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_560),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_552),
.B(n_472),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_563),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_563),
.Y(n_683)
);

AOI22x1_ASAP7_75t_L g684 ( 
.A1(n_522),
.A2(n_260),
.B1(n_280),
.B2(n_265),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_568),
.B(n_475),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_588),
.B(n_463),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_563),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_563),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_563),
.B(n_247),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_563),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_563),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_566),
.B(n_247),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_566),
.Y(n_693)
);

AOI21x1_ASAP7_75t_L g694 ( 
.A1(n_516),
.A2(n_412),
.B(n_366),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_566),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_566),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_588),
.B(n_395),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_566),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_566),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_SL g700 ( 
.A1(n_578),
.A2(n_395),
.B1(n_279),
.B2(n_283),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_566),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_592),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_592),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_519),
.A2(n_479),
.B1(n_491),
.B2(n_489),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_519),
.B(n_414),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_592),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_568),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_577),
.B(n_514),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_553),
.B(n_503),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_577),
.B(n_496),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_577),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_536),
.B(n_501),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_592),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_577),
.B(n_502),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_595),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_592),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_595),
.B(n_509),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_595),
.B(n_407),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_578),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_580),
.B(n_222),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_592),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_536),
.B(n_380),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_592),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_525),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_580),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_516),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_529),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_541),
.B(n_363),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_541),
.A2(n_280),
.B1(n_260),
.B2(n_222),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_553),
.A2(n_272),
.B1(n_291),
.B2(n_287),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_546),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_546),
.B(n_363),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_529),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_553),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_542),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_547),
.A2(n_280),
.B1(n_327),
.B2(n_311),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_529),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_547),
.B(n_511),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_549),
.B(n_413),
.Y(n_739)
);

INVx4_ASAP7_75t_SL g740 ( 
.A(n_553),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_L g741 ( 
.A(n_549),
.B(n_247),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_525),
.Y(n_742)
);

BUFx2_ASAP7_75t_L g743 ( 
.A(n_553),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_527),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_551),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_527),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_551),
.B(n_513),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_559),
.B(n_515),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_735),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_L g750 ( 
.A(n_643),
.B(n_416),
.C(n_265),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_610),
.B(n_424),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_712),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_735),
.Y(n_753)
);

AND2x2_ASAP7_75t_SL g754 ( 
.A(n_621),
.B(n_275),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_724),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_738),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_621),
.B(n_559),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_726),
.B(n_569),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_719),
.B(n_569),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_602),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_SL g761 ( 
.A(n_642),
.B(n_438),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_719),
.B(n_571),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_621),
.A2(n_599),
.B1(n_573),
.B2(n_576),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_735),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_725),
.B(n_571),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_604),
.B(n_573),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_724),
.Y(n_767)
);

INVx8_ASAP7_75t_L g768 ( 
.A(n_628),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_742),
.Y(n_769)
);

BUFx5_ASAP7_75t_L g770 ( 
.A(n_665),
.Y(n_770)
);

AND2x6_ASAP7_75t_L g771 ( 
.A(n_634),
.B(n_576),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_742),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_604),
.B(n_579),
.Y(n_773)
);

AO221x1_ASAP7_75t_L g774 ( 
.A1(n_673),
.A2(n_662),
.B1(n_743),
.B2(n_734),
.C(n_256),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_626),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_628),
.A2(n_582),
.B1(n_583),
.B2(n_579),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_612),
.A2(n_599),
.B1(n_583),
.B2(n_584),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_744),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_744),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_725),
.B(n_582),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_L g781 ( 
.A(n_731),
.B(n_584),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_746),
.Y(n_782)
);

OR2x6_ASAP7_75t_L g783 ( 
.A(n_697),
.B(n_542),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_646),
.B(n_585),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_646),
.A2(n_587),
.B1(n_593),
.B2(n_585),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_649),
.B(n_587),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_634),
.B(n_593),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_670),
.B(n_594),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_654),
.B(n_686),
.C(n_676),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_718),
.B(n_594),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_652),
.A2(n_597),
.B1(n_596),
.B2(n_555),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_739),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_646),
.B(n_616),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_616),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_746),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_747),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_718),
.B(n_596),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_745),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_652),
.B(n_597),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_667),
.B(n_545),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_606),
.B(n_545),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_671),
.B(n_545),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_671),
.B(n_555),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_731),
.B(n_555),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_616),
.B(n_556),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_603),
.A2(n_564),
.B(n_556),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_642),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_600),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_709),
.A2(n_442),
.B1(n_470),
.B2(n_445),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_715),
.B(n_708),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_607),
.A2(n_556),
.B1(n_565),
.B2(n_564),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_739),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_715),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_608),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_748),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_634),
.A2(n_565),
.B1(n_570),
.B2(n_564),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_623),
.B(n_565),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_608),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_657),
.B(n_570),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_707),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_685),
.B(n_570),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_602),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_611),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_611),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_707),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_602),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_710),
.B(n_572),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_602),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_661),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_722),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_714),
.B(n_572),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_661),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_657),
.B(n_574),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_664),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_645),
.Y(n_835)
);

OR2x6_ASAP7_75t_L g836 ( 
.A(n_697),
.B(n_574),
.Y(n_836)
);

NAND2xp33_ASAP7_75t_L g837 ( 
.A(n_622),
.B(n_581),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_628),
.A2(n_591),
.B1(n_581),
.B2(n_562),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_L g839 ( 
.A(n_625),
.B(n_591),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_645),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_L g841 ( 
.A(n_623),
.B(n_591),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_628),
.A2(n_562),
.B1(n_553),
.B2(n_388),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_708),
.B(n_531),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_657),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_668),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_615),
.B(n_531),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_665),
.A2(n_562),
.B1(n_553),
.B2(n_533),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_648),
.A2(n_562),
.B1(n_553),
.B2(n_388),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_648),
.B(n_533),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_613),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_619),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_631),
.B(n_553),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_609),
.B(n_562),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_619),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_717),
.B(n_293),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_681),
.B(n_251),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_629),
.Y(n_857)
);

AOI221xp5_ASAP7_75t_L g858 ( 
.A1(n_630),
.A2(n_338),
.B1(n_347),
.B2(n_351),
.C(n_251),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_711),
.B(n_636),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_681),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_711),
.B(n_366),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_SL g862 ( 
.A(n_711),
.B(n_267),
.Y(n_862)
);

OAI22x1_ASAP7_75t_SL g863 ( 
.A1(n_697),
.A2(n_374),
.B1(n_410),
.B2(n_409),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_605),
.B(n_368),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_601),
.B(n_208),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_655),
.B(n_295),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_728),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_629),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_732),
.A2(n_281),
.B(n_267),
.C(n_282),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_720),
.B(n_562),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_637),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_675),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_659),
.B(n_302),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_675),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_720),
.B(n_562),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_617),
.B(n_407),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_675),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_663),
.B(n_307),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_697),
.B(n_281),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_720),
.B(n_562),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_603),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_614),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_605),
.B(n_356),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_605),
.B(n_356),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_665),
.A2(n_720),
.B1(n_684),
.B2(n_729),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_672),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_605),
.B(n_247),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_605),
.B(n_247),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_614),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_637),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_639),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_704),
.B(n_407),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_665),
.B(n_230),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_633),
.B(n_705),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_665),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_618),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_730),
.B(n_734),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_639),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_665),
.B(n_230),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_635),
.B(n_313),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_618),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_620),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_650),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_721),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_620),
.Y(n_905)
);

INVx4_ASAP7_75t_L g906 ( 
.A(n_740),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_624),
.Y(n_907)
);

CKINVDCx16_ASAP7_75t_R g908 ( 
.A(n_743),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_677),
.B(n_247),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_624),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_736),
.B(n_311),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_721),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_756),
.A2(n_700),
.B(n_297),
.C(n_314),
.Y(n_913)
);

CKINVDCx10_ASAP7_75t_R g914 ( 
.A(n_761),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_810),
.B(n_635),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_758),
.B(n_635),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_906),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_SL g918 ( 
.A(n_789),
.B(n_638),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_752),
.B(n_638),
.Y(n_919)
);

CKINVDCx8_ASAP7_75t_R g920 ( 
.A(n_807),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_859),
.A2(n_632),
.B(n_627),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_841),
.B(n_638),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_754),
.B(n_677),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_781),
.A2(n_632),
.B(n_627),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_805),
.A2(n_833),
.B(n_819),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_867),
.B(n_669),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_754),
.A2(n_741),
.B(n_695),
.C(n_698),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_796),
.A2(n_741),
.B1(n_695),
.B2(n_698),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_805),
.A2(n_641),
.B(n_640),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_819),
.A2(n_641),
.B(n_640),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_815),
.B(n_669),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_759),
.B(n_669),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_833),
.A2(n_647),
.B(n_644),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_775),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_837),
.A2(n_647),
.B(n_644),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_770),
.B(n_677),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_762),
.B(n_695),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_834),
.B(n_698),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_765),
.B(n_723),
.Y(n_939)
);

OAI21xp33_ASAP7_75t_L g940 ( 
.A1(n_855),
.A2(n_332),
.B(n_331),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_886),
.B(n_723),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_839),
.A2(n_788),
.B(n_786),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_804),
.A2(n_674),
.B(n_651),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_793),
.A2(n_852),
.B(n_797),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_793),
.A2(n_674),
.B(n_651),
.Y(n_945)
);

AO22x1_ASAP7_75t_L g946 ( 
.A1(n_892),
.A2(n_341),
.B1(n_345),
.B2(n_340),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_780),
.B(n_723),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_790),
.A2(n_679),
.B(n_678),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_778),
.A2(n_687),
.B1(n_690),
.B2(n_680),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_821),
.B(n_680),
.Y(n_950)
);

OAI21xp33_ASAP7_75t_L g951 ( 
.A1(n_855),
.A2(n_361),
.B(n_359),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_853),
.A2(n_690),
.B(n_687),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_799),
.A2(n_696),
.B(n_693),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_800),
.A2(n_696),
.B(n_693),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_906),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_770),
.B(n_677),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_SL g957 ( 
.A1(n_861),
.A2(n_713),
.B(n_706),
.C(n_703),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_860),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_766),
.A2(n_702),
.B1(n_703),
.B2(n_706),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_846),
.A2(n_713),
.B(n_702),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_782),
.A2(n_795),
.B1(n_767),
.B2(n_769),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_821),
.B(n_650),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_795),
.A2(n_682),
.B1(n_653),
.B2(n_660),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_827),
.B(n_831),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_770),
.B(n_776),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_846),
.A2(n_660),
.B(n_653),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_784),
.A2(n_682),
.B(n_666),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_792),
.B(n_407),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_827),
.B(n_666),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_801),
.A2(n_688),
.B(n_683),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_801),
.A2(n_683),
.B(n_688),
.C(n_691),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_904),
.Y(n_972)
);

AOI221xp5_ASAP7_75t_L g973 ( 
.A1(n_858),
.A2(n_362),
.B1(n_330),
.B2(n_376),
.C(n_321),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_784),
.A2(n_699),
.B(n_691),
.Y(n_974)
);

OAI21xp33_ASAP7_75t_L g975 ( 
.A1(n_813),
.A2(n_369),
.B(n_365),
.Y(n_975)
);

BUFx8_ASAP7_75t_L g976 ( 
.A(n_845),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_757),
.A2(n_701),
.B(n_699),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_831),
.A2(n_716),
.B(n_701),
.C(n_689),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_760),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_904),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_770),
.B(n_677),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_755),
.Y(n_982)
);

OR2x6_ASAP7_75t_L g983 ( 
.A(n_768),
.B(n_783),
.Y(n_983)
);

AND2x6_ASAP7_75t_L g984 ( 
.A(n_874),
.B(n_716),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_772),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_829),
.A2(n_832),
.B(n_766),
.C(n_773),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_779),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_843),
.B(n_727),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_835),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_773),
.A2(n_689),
.B1(n_692),
.B2(n_733),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_808),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_770),
.B(n_656),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_806),
.A2(n_694),
.B(n_733),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_770),
.B(n_656),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_840),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_887),
.A2(n_694),
.B(n_520),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_757),
.A2(n_861),
.B(n_844),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_760),
.Y(n_998)
);

NOR2x2_ASAP7_75t_L g999 ( 
.A(n_783),
.B(n_327),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_817),
.B(n_684),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_912),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_830),
.B(n_737),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_849),
.B(n_737),
.Y(n_1003)
);

AO21x1_ASAP7_75t_L g1004 ( 
.A1(n_883),
.A2(n_692),
.B(n_297),
.Y(n_1004)
);

INVx11_ASAP7_75t_L g1005 ( 
.A(n_771),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_763),
.B(n_737),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_791),
.A2(n_658),
.B(n_656),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_802),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_794),
.A2(n_658),
.B(n_656),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_808),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_894),
.B(n_737),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_794),
.A2(n_658),
.B(n_656),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_844),
.A2(n_658),
.B(n_737),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_812),
.B(n_282),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_749),
.A2(n_520),
.B(n_517),
.Y(n_1015)
);

OAI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_900),
.A2(n_377),
.B(n_370),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_895),
.B(n_740),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_749),
.A2(n_520),
.B(n_517),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_881),
.A2(n_528),
.B(n_517),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_753),
.A2(n_528),
.B(n_211),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_887),
.A2(n_528),
.B(n_321),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_751),
.B(n_314),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_783),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_798),
.B(n_330),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_803),
.Y(n_1025)
);

AOI21x1_ASAP7_75t_L g1026 ( 
.A1(n_888),
.A2(n_347),
.B(n_338),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_809),
.B(n_351),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_882),
.A2(n_364),
.B(n_362),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_912),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_885),
.A2(n_771),
.B1(n_774),
.B2(n_878),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_753),
.B(n_764),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_764),
.A2(n_896),
.B(n_889),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_750),
.A2(n_376),
.B(n_364),
.C(n_367),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_836),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_901),
.A2(n_214),
.B(n_210),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_777),
.B(n_367),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_902),
.A2(n_389),
.B(n_371),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_811),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_822),
.B(n_740),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_905),
.A2(n_389),
.B(n_371),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_771),
.B(n_822),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_907),
.A2(n_220),
.B(n_215),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_785),
.A2(n_393),
.B1(n_402),
.B2(n_394),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_856),
.A2(n_400),
.B(n_399),
.C(n_333),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_771),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_874),
.B(n_740),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_771),
.B(n_400),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_910),
.A2(n_236),
.B(n_233),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_885),
.B(n_219),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_826),
.B(n_387),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_872),
.B(n_333),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_828),
.B(n_390),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_876),
.B(n_391),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_878),
.B(n_404),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_838),
.B(n_877),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_836),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_908),
.B(n_399),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_L g1058 ( 
.A1(n_888),
.A2(n_524),
.B(n_523),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_820),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_814),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_825),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_814),
.A2(n_242),
.B(n_239),
.Y(n_1062)
);

BUFx12f_ASAP7_75t_L g1063 ( 
.A(n_879),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_866),
.A2(n_256),
.B(n_219),
.C(n_535),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_818),
.A2(n_824),
.B(n_823),
.Y(n_1065)
);

INVxp67_ASAP7_75t_L g1066 ( 
.A(n_787),
.Y(n_1066)
);

NOR2xp67_ASAP7_75t_L g1067 ( 
.A(n_866),
.B(n_246),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_842),
.B(n_219),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_816),
.B(n_256),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_824),
.A2(n_306),
.B(n_252),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_L g1071 ( 
.A1(n_909),
.A2(n_884),
.B(n_883),
.Y(n_1071)
);

OAI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_900),
.A2(n_873),
.B(n_862),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_768),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_897),
.A2(n_871),
.B1(n_857),
.B2(n_903),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_850),
.A2(n_315),
.B(n_255),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_851),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_870),
.B(n_256),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_863),
.Y(n_1078)
);

NOR3xp33_ASAP7_75t_L g1079 ( 
.A(n_873),
.B(n_354),
.C(n_290),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_909),
.A2(n_868),
.B(n_903),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_884),
.A2(n_524),
.B(n_523),
.Y(n_1081)
);

BUFx12f_ASAP7_75t_SL g1082 ( 
.A(n_865),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_869),
.Y(n_1083)
);

AO21x1_ASAP7_75t_L g1084 ( 
.A1(n_864),
.A2(n_247),
.B(n_529),
.Y(n_1084)
);

AOI21x1_ASAP7_75t_L g1085 ( 
.A1(n_864),
.A2(n_524),
.B(n_523),
.Y(n_1085)
);

AND2x2_ASAP7_75t_SL g1086 ( 
.A(n_847),
.B(n_256),
.Y(n_1086)
);

INVx4_ASAP7_75t_L g1087 ( 
.A(n_854),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_893),
.A2(n_535),
.B(n_529),
.C(n_320),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_964),
.A2(n_868),
.B(n_854),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_1054),
.A2(n_899),
.B(n_875),
.C(n_880),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_934),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_982),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1054),
.B(n_857),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_918),
.A2(n_847),
.B(n_898),
.C(n_891),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1086),
.A2(n_898),
.B1(n_891),
.B2(n_890),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1038),
.B(n_911),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_934),
.Y(n_1097)
);

CKINVDCx8_ASAP7_75t_R g1098 ( 
.A(n_914),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1072),
.A2(n_890),
.B(n_871),
.C(n_23),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_958),
.B(n_848),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_1079),
.B(n_535),
.C(n_529),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1086),
.A2(n_319),
.B1(n_250),
.B2(n_408),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_SL g1103 ( 
.A1(n_920),
.A2(n_379),
.B1(n_274),
.B2(n_271),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1081),
.A2(n_535),
.B(n_529),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_942),
.A2(n_524),
.B(n_523),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_944),
.A2(n_524),
.B(n_523),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1008),
.B(n_20),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_950),
.A2(n_524),
.B(n_523),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1079),
.A2(n_535),
.B(n_323),
.C(n_303),
.Y(n_1109)
);

AOI33xp33_ASAP7_75t_L g1110 ( 
.A1(n_1022),
.A2(n_20),
.A3(n_22),
.B1(n_23),
.B2(n_25),
.B3(n_30),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_1045),
.B(n_248),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_961),
.A2(n_985),
.B1(n_987),
.B2(n_919),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_983),
.B(n_535),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_925),
.A2(n_328),
.B(n_261),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_1088),
.A2(n_1084),
.A3(n_1074),
.B(n_971),
.Y(n_1115)
);

INVx3_ASAP7_75t_SL g1116 ( 
.A(n_999),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_976),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1033),
.A2(n_31),
.B(n_32),
.C(n_34),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_986),
.A2(n_535),
.B(n_324),
.C(n_301),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_958),
.B(n_259),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_965),
.A2(n_524),
.B(n_523),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_976),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_989),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1063),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_940),
.A2(n_34),
.B(n_38),
.C(n_40),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_955),
.Y(n_1126)
);

NAND2x1p5_ASAP7_75t_L g1127 ( 
.A(n_1045),
.B(n_78),
.Y(n_1127)
);

O2A1O1Ixp5_ASAP7_75t_L g1128 ( 
.A1(n_965),
.A2(n_247),
.B(n_42),
.C(n_44),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1073),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1025),
.B(n_41),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_946),
.B(n_41),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_962),
.A2(n_300),
.B(n_401),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1073),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_1073),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_951),
.A2(n_406),
.B(n_398),
.C(n_392),
.Y(n_1135)
);

INVxp67_ASAP7_75t_SL g1136 ( 
.A(n_1049),
.Y(n_1136)
);

AND2x2_ASAP7_75t_SL g1137 ( 
.A(n_1030),
.B(n_1045),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1045),
.B(n_262),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_969),
.A2(n_298),
.B(n_381),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1014),
.B(n_45),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_991),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_997),
.A2(n_382),
.B(n_373),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_919),
.B(n_1066),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1067),
.A2(n_1028),
.B(n_1040),
.C(n_1037),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1016),
.A2(n_355),
.B(n_353),
.C(n_352),
.Y(n_1145)
);

BUFx10_ASAP7_75t_L g1146 ( 
.A(n_1050),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1010),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_995),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_952),
.A2(n_288),
.B(n_346),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1057),
.Y(n_1150)
);

INVx5_ASAP7_75t_L g1151 ( 
.A(n_984),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1049),
.A2(n_349),
.B(n_344),
.C(n_343),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1053),
.B(n_46),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1073),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1058),
.A2(n_247),
.B(n_130),
.Y(n_1155)
);

AOI22x1_ASAP7_75t_L g1156 ( 
.A1(n_948),
.A2(n_334),
.B1(n_299),
.B2(n_296),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1059),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1066),
.B(n_46),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_968),
.B(n_48),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1060),
.Y(n_1160)
);

OAI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_1043),
.A2(n_294),
.B(n_286),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1030),
.A2(n_285),
.B(n_284),
.C(n_277),
.Y(n_1162)
);

AO22x1_ASAP7_75t_L g1163 ( 
.A1(n_1027),
.A2(n_269),
.B1(n_266),
.B2(n_264),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1083),
.B(n_49),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1000),
.A2(n_49),
.B(n_51),
.C(n_56),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1023),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1036),
.B(n_51),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1050),
.B(n_56),
.Y(n_1168)
);

INVxp67_ASAP7_75t_SL g1169 ( 
.A(n_1006),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1061),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_960),
.A2(n_57),
.B(n_60),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_921),
.A2(n_61),
.B(n_65),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_931),
.A2(n_61),
.B1(n_67),
.B2(n_68),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_923),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1024),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_954),
.A2(n_72),
.B(n_74),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_979),
.B(n_82),
.Y(n_1177)
);

OAI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1052),
.A2(n_85),
.B(n_87),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_915),
.A2(n_92),
.B(n_95),
.C(n_98),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_975),
.B(n_101),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1034),
.Y(n_1181)
);

INVxp67_ASAP7_75t_L g1182 ( 
.A(n_1011),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_916),
.A2(n_103),
.B(n_108),
.C(n_115),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1032),
.A2(n_117),
.B(n_121),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1003),
.A2(n_122),
.B(n_131),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_928),
.A2(n_134),
.B1(n_138),
.B2(n_143),
.Y(n_1186)
);

OR2x6_ASAP7_75t_SL g1187 ( 
.A(n_1047),
.B(n_149),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1005),
.A2(n_155),
.B1(n_170),
.B2(n_175),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_926),
.A2(n_177),
.B1(n_184),
.B2(n_187),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_983),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1052),
.B(n_938),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_938),
.B(n_192),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_979),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_966),
.A2(n_202),
.B(n_206),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_978),
.A2(n_957),
.B(n_988),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_941),
.B(n_1082),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_998),
.B(n_955),
.Y(n_1197)
);

AOI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1085),
.A2(n_996),
.B(n_1071),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_917),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1055),
.A2(n_1044),
.B(n_953),
.C(n_927),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_998),
.Y(n_1201)
);

AO22x1_ASAP7_75t_L g1202 ( 
.A1(n_1078),
.A2(n_1056),
.B1(n_984),
.B2(n_998),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_973),
.B(n_972),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1076),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_932),
.A2(n_937),
.B1(n_939),
.B2(n_947),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_980),
.A2(n_1029),
.B1(n_1001),
.B2(n_1041),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_957),
.A2(n_945),
.B(n_935),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_917),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_983),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1087),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1087),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1051),
.A2(n_913),
.B1(n_1001),
.B2(n_1029),
.Y(n_1212)
);

OAI21xp33_ASAP7_75t_L g1213 ( 
.A1(n_1035),
.A2(n_1048),
.B(n_1042),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_984),
.Y(n_1214)
);

BUFx10_ASAP7_75t_L g1215 ( 
.A(n_984),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_984),
.B(n_1002),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1026),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_959),
.A2(n_949),
.B1(n_1007),
.B2(n_922),
.Y(n_1218)
);

AO21x1_ASAP7_75t_L g1219 ( 
.A1(n_1077),
.A2(n_981),
.B(n_956),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_943),
.A2(n_974),
.B(n_967),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1069),
.A2(n_1031),
.B1(n_1039),
.B2(n_1068),
.Y(n_1221)
);

OA22x2_ASAP7_75t_L g1222 ( 
.A1(n_1080),
.A2(n_990),
.B1(n_1031),
.B2(n_1046),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_977),
.A2(n_929),
.B(n_930),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1077),
.B(n_1046),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1069),
.A2(n_1068),
.B1(n_936),
.B2(n_956),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_963),
.B(n_970),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1021),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1064),
.A2(n_1088),
.B(n_1075),
.C(n_1070),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1065),
.B(n_933),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1062),
.B(n_1017),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_936),
.B(n_981),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_993),
.A2(n_1004),
.B(n_1020),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1017),
.B(n_924),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_992),
.B(n_994),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_992),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1190),
.B(n_994),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1098),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1144),
.A2(n_1019),
.B(n_1013),
.C(n_1015),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_1125),
.B(n_1018),
.C(n_1009),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1187),
.A2(n_1012),
.B1(n_1168),
.B2(n_1131),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1191),
.A2(n_1143),
.B1(n_1112),
.B2(n_1100),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1205),
.A2(n_1218),
.B(n_1195),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1091),
.B(n_1175),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1195),
.A2(n_1207),
.B(n_1220),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1207),
.A2(n_1220),
.B(n_1226),
.Y(n_1245)
);

NAND3xp33_ASAP7_75t_L g1246 ( 
.A(n_1125),
.B(n_1118),
.C(n_1165),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1108),
.A2(n_1093),
.B(n_1192),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1117),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1099),
.A2(n_1178),
.B(n_1162),
.C(n_1180),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1092),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1202),
.B(n_1124),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1118),
.A2(n_1200),
.B(n_1173),
.C(n_1167),
.Y(n_1252)
);

NAND2xp33_ASAP7_75t_L g1253 ( 
.A(n_1151),
.B(n_1109),
.Y(n_1253)
);

CKINVDCx11_ASAP7_75t_R g1254 ( 
.A(n_1122),
.Y(n_1254)
);

AOI21xp33_ASAP7_75t_L g1255 ( 
.A1(n_1102),
.A2(n_1099),
.B(n_1161),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_SL g1256 ( 
.A(n_1151),
.B(n_1137),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1198),
.Y(n_1257)
);

OAI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1174),
.A2(n_1140),
.B1(n_1159),
.B2(n_1203),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1153),
.A2(n_1164),
.B1(n_1212),
.B2(n_1097),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1129),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1150),
.B(n_1163),
.Y(n_1261)
);

AO32x2_ASAP7_75t_L g1262 ( 
.A1(n_1095),
.A2(n_1206),
.A3(n_1186),
.B1(n_1189),
.B2(n_1169),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1089),
.A2(n_1223),
.B(n_1106),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1106),
.A2(n_1155),
.B(n_1121),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1157),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_1166),
.B(n_1181),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1116),
.B(n_1120),
.Y(n_1267)
);

AOI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1222),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1170),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_SL g1270 ( 
.A1(n_1090),
.A2(n_1130),
.B(n_1107),
.C(n_1094),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1116),
.Y(n_1271)
);

NOR2xp67_ASAP7_75t_L g1272 ( 
.A(n_1151),
.B(n_1199),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1146),
.B(n_1123),
.Y(n_1273)
);

AOI211x1_ASAP7_75t_L g1274 ( 
.A1(n_1171),
.A2(n_1176),
.B(n_1172),
.C(n_1158),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1103),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1233),
.A2(n_1194),
.B(n_1217),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1165),
.A2(n_1128),
.B(n_1171),
.C(n_1176),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1213),
.A2(n_1216),
.B(n_1151),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1196),
.B(n_1129),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1129),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1194),
.A2(n_1217),
.B(n_1184),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1193),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1101),
.A2(n_1114),
.B(n_1132),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1224),
.C(n_1139),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1184),
.A2(n_1228),
.B(n_1230),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1133),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1169),
.A2(n_1136),
.B(n_1225),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_SL g1288 ( 
.A(n_1126),
.B(n_1154),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1148),
.B(n_1110),
.Y(n_1289)
);

NOR2xp67_ASAP7_75t_SL g1290 ( 
.A(n_1126),
.B(n_1133),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1228),
.A2(n_1234),
.B(n_1149),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1149),
.A2(n_1185),
.B(n_1132),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1139),
.A2(n_1172),
.B(n_1183),
.C(n_1179),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1152),
.A2(n_1145),
.B(n_1135),
.Y(n_1294)
);

BUFx5_ASAP7_75t_L g1295 ( 
.A(n_1215),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1185),
.A2(n_1119),
.B(n_1179),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1133),
.Y(n_1297)
);

AO21x1_ASAP7_75t_L g1298 ( 
.A1(n_1183),
.A2(n_1136),
.B(n_1177),
.Y(n_1298)
);

BUFx12f_ASAP7_75t_L g1299 ( 
.A(n_1154),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1221),
.A2(n_1208),
.B1(n_1199),
.B2(n_1182),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1208),
.A2(n_1214),
.B(n_1197),
.Y(n_1301)
);

AO22x2_ASAP7_75t_L g1302 ( 
.A1(n_1204),
.A2(n_1160),
.B1(n_1147),
.B2(n_1141),
.Y(n_1302)
);

INVx5_ASAP7_75t_L g1303 ( 
.A(n_1215),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1096),
.A2(n_1111),
.B(n_1138),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1127),
.A2(n_1210),
.B(n_1211),
.Y(n_1305)
);

O2A1O1Ixp5_ASAP7_75t_SL g1306 ( 
.A1(n_1201),
.A2(n_1209),
.B(n_1188),
.C(n_1115),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1134),
.B(n_1154),
.Y(n_1307)
);

OAI21xp33_ASAP7_75t_L g1308 ( 
.A1(n_1156),
.A2(n_1127),
.B(n_1235),
.Y(n_1308)
);

NOR2xp67_ASAP7_75t_SL g1309 ( 
.A(n_1193),
.B(n_1235),
.Y(n_1309)
);

AOI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1113),
.A2(n_1105),
.B(n_1104),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1113),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1115),
.B(n_860),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1144),
.A2(n_756),
.B(n_815),
.C(n_796),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_789),
.C(n_1093),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1144),
.A2(n_756),
.B(n_815),
.C(n_796),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1091),
.B(n_860),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1191),
.A2(n_754),
.B1(n_796),
.B2(n_756),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1129),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1122),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1190),
.B(n_1073),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1091),
.B(n_860),
.Y(n_1323)
);

OAI21xp33_ASAP7_75t_L g1324 ( 
.A1(n_1168),
.A2(n_1054),
.B(n_796),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_SL g1325 ( 
.A1(n_1112),
.A2(n_986),
.B(n_1099),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1198),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1098),
.Y(n_1327)
);

AOI31xp67_ASAP7_75t_L g1328 ( 
.A1(n_1222),
.A2(n_1226),
.A3(n_1227),
.B(n_1229),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1092),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_SL g1330 ( 
.A1(n_1144),
.A2(n_1191),
.B(n_1168),
.C(n_1109),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_SL g1332 ( 
.A1(n_1144),
.A2(n_1191),
.B(n_1168),
.C(n_1109),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_789),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1198),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1124),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1091),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1191),
.A2(n_754),
.B1(n_796),
.B2(n_756),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1091),
.B(n_958),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1190),
.B(n_1073),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_789),
.C(n_1093),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1105),
.A2(n_1104),
.B(n_1106),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1091),
.B(n_1097),
.Y(n_1342)
);

O2A1O1Ixp5_ASAP7_75t_SL g1343 ( 
.A1(n_1231),
.A2(n_1217),
.B(n_1226),
.C(n_1182),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1092),
.Y(n_1345)
);

O2A1O1Ixp5_ASAP7_75t_SL g1346 ( 
.A1(n_1231),
.A2(n_1217),
.B(n_1226),
.C(n_1182),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1091),
.B(n_860),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_789),
.Y(n_1350)
);

AO21x1_ASAP7_75t_L g1351 ( 
.A1(n_1099),
.A2(n_1054),
.B(n_1168),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1098),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_789),
.C(n_1093),
.Y(n_1353)
);

INVx3_ASAP7_75t_SL g1354 ( 
.A(n_1117),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1091),
.B(n_958),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1091),
.B(n_1097),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1357)
);

AOI221x1_ASAP7_75t_L g1358 ( 
.A1(n_1178),
.A2(n_1144),
.B1(n_1171),
.B2(n_1162),
.C(n_1176),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1168),
.A2(n_761),
.B1(n_815),
.B2(n_796),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1129),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_789),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_SL g1363 ( 
.A1(n_1112),
.A2(n_986),
.B(n_1099),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1198),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1124),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1092),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1129),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1198),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_SL g1370 ( 
.A1(n_1144),
.A2(n_1191),
.B(n_1168),
.C(n_1109),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1198),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1091),
.B(n_860),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1198),
.Y(n_1374)
);

INVx3_ASAP7_75t_SL g1375 ( 
.A(n_1117),
.Y(n_1375)
);

AOI21xp33_ASAP7_75t_L g1376 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_796),
.Y(n_1376)
);

NAND3x1_ASAP7_75t_L g1377 ( 
.A(n_1164),
.B(n_1196),
.C(n_1131),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1219),
.A2(n_1108),
.A3(n_1088),
.B(n_1084),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1144),
.A2(n_756),
.B(n_815),
.C(n_796),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1091),
.Y(n_1381)
);

AO31x2_ASAP7_75t_L g1382 ( 
.A1(n_1219),
.A2(n_1108),
.A3(n_1088),
.B(n_1084),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_789),
.C(n_1093),
.Y(n_1384)
);

AOI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1105),
.A2(n_1104),
.B(n_1106),
.Y(n_1385)
);

NAND3x1_ASAP7_75t_L g1386 ( 
.A(n_1164),
.B(n_1196),
.C(n_1131),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1097),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1198),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1205),
.A2(n_964),
.B(n_1072),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1091),
.B(n_860),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1091),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1144),
.A2(n_756),
.B(n_815),
.C(n_796),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1190),
.B(n_1073),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1286),
.Y(n_1394)
);

INVx4_ASAP7_75t_L g1395 ( 
.A(n_1299),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1324),
.A2(n_1246),
.B1(n_1258),
.B2(n_1376),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1324),
.A2(n_1246),
.B1(n_1259),
.B2(n_1361),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1259),
.A2(n_1333),
.B1(n_1350),
.B2(n_1241),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1250),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1260),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1327),
.Y(n_1401)
);

INVx8_ASAP7_75t_L g1402 ( 
.A(n_1320),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1314),
.A2(n_1384),
.B1(n_1353),
.B2(n_1340),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1318),
.A2(n_1337),
.B1(n_1242),
.B2(n_1331),
.Y(n_1404)
);

BUFx12f_ASAP7_75t_L g1405 ( 
.A(n_1237),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1265),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1256),
.A2(n_1240),
.B1(n_1325),
.B2(n_1363),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1269),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1329),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1352),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1317),
.A2(n_1357),
.B1(n_1368),
.B2(n_1344),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_SL g1412 ( 
.A(n_1365),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1351),
.A2(n_1256),
.B1(n_1359),
.B2(n_1261),
.Y(n_1413)
);

CKINVDCx11_ASAP7_75t_R g1414 ( 
.A(n_1354),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1312),
.B(n_1321),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1289),
.A2(n_1275),
.B1(n_1255),
.B2(n_1240),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1358),
.A2(n_1383),
.B1(n_1379),
.B2(n_1389),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1260),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1348),
.A2(n_1371),
.B1(n_1362),
.B2(n_1349),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1266),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1243),
.A2(n_1283),
.B1(n_1267),
.B2(n_1251),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1266),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1252),
.A2(n_1274),
.B1(n_1392),
.B2(n_1315),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1345),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1366),
.Y(n_1425)
);

BUFx2_ASAP7_75t_SL g1426 ( 
.A(n_1338),
.Y(n_1426)
);

BUFx8_ASAP7_75t_L g1427 ( 
.A(n_1387),
.Y(n_1427)
);

BUFx8_ASAP7_75t_L g1428 ( 
.A(n_1355),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1254),
.Y(n_1429)
);

BUFx12f_ASAP7_75t_L g1430 ( 
.A(n_1248),
.Y(n_1430)
);

CKINVDCx11_ASAP7_75t_R g1431 ( 
.A(n_1375),
.Y(n_1431)
);

BUFx8_ASAP7_75t_L g1432 ( 
.A(n_1273),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1302),
.Y(n_1433)
);

BUFx12f_ASAP7_75t_L g1434 ( 
.A(n_1266),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1302),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1342),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1381),
.A2(n_1316),
.B1(n_1323),
.B2(n_1390),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1336),
.B(n_1391),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1356),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1347),
.A2(n_1373),
.B1(n_1251),
.B2(n_1294),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1311),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1251),
.A2(n_1300),
.B1(n_1291),
.B2(n_1271),
.Y(n_1442)
);

INVx8_ASAP7_75t_L g1443 ( 
.A(n_1303),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1253),
.A2(n_1287),
.B1(n_1386),
.B2(n_1377),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1236),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1236),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1328),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1298),
.A2(n_1308),
.B1(n_1296),
.B2(n_1287),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1308),
.A2(n_1304),
.B1(n_1292),
.B2(n_1393),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1307),
.Y(n_1450)
);

BUFx4_ASAP7_75t_R g1451 ( 
.A(n_1295),
.Y(n_1451)
);

INVx5_ASAP7_75t_L g1452 ( 
.A(n_1319),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1322),
.A2(n_1393),
.B1(n_1339),
.B2(n_1279),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1274),
.A2(n_1380),
.B1(n_1313),
.B2(n_1249),
.Y(n_1454)
);

OAI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1247),
.A2(n_1272),
.B1(n_1268),
.B2(n_1245),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1239),
.A2(n_1277),
.B1(n_1295),
.B2(n_1285),
.Y(n_1456)
);

BUFx2_ASAP7_75t_SL g1457 ( 
.A(n_1360),
.Y(n_1457)
);

BUFx8_ASAP7_75t_L g1458 ( 
.A(n_1367),
.Y(n_1458)
);

BUFx12f_ASAP7_75t_L g1459 ( 
.A(n_1367),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1284),
.A2(n_1293),
.B1(n_1244),
.B2(n_1239),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1367),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1263),
.A2(n_1272),
.B1(n_1330),
.B2(n_1332),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1280),
.A2(n_1297),
.B1(n_1282),
.B2(n_1301),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1370),
.A2(n_1339),
.B1(n_1309),
.B2(n_1290),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1295),
.A2(n_1288),
.B1(n_1278),
.B2(n_1305),
.Y(n_1465)
);

BUFx4_ASAP7_75t_R g1466 ( 
.A(n_1295),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1276),
.A2(n_1281),
.B1(n_1264),
.B2(n_1270),
.Y(n_1467)
);

CKINVDCx11_ASAP7_75t_R g1468 ( 
.A(n_1306),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1257),
.A2(n_1364),
.B1(n_1374),
.B2(n_1372),
.Y(n_1469)
);

INVx8_ASAP7_75t_L g1470 ( 
.A(n_1343),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1346),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1326),
.A2(n_1369),
.B1(n_1388),
.B2(n_1334),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1262),
.A2(n_1378),
.B1(n_1382),
.B2(n_1238),
.Y(n_1473)
);

BUFx8_ASAP7_75t_SL g1474 ( 
.A(n_1310),
.Y(n_1474)
);

BUFx12f_ASAP7_75t_L g1475 ( 
.A(n_1262),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1262),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1341),
.A2(n_1385),
.B1(n_1378),
.B2(n_1382),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1382),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1324),
.A2(n_809),
.B1(n_1054),
.B2(n_754),
.Y(n_1479)
);

INVx8_ASAP7_75t_L g1480 ( 
.A(n_1286),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1241),
.A2(n_754),
.B1(n_1340),
.B2(n_1314),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1324),
.A2(n_809),
.B1(n_1054),
.B2(n_754),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1246),
.A2(n_754),
.B1(n_1137),
.B2(n_1086),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1286),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1327),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1241),
.B(n_1169),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1250),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1250),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1250),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1250),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1250),
.Y(n_1491)
);

BUFx5_ASAP7_75t_L g1492 ( 
.A(n_1236),
.Y(n_1492)
);

CKINVDCx11_ASAP7_75t_R g1493 ( 
.A(n_1327),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1250),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1246),
.A2(n_754),
.B1(n_1137),
.B2(n_1086),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1327),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1250),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1250),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1241),
.B(n_1169),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1250),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1335),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1266),
.Y(n_1502)
);

CKINVDCx11_ASAP7_75t_R g1503 ( 
.A(n_1327),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1338),
.B(n_1355),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1335),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1324),
.A2(n_809),
.B1(n_1054),
.B2(n_754),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1324),
.A2(n_809),
.B1(n_1054),
.B2(n_754),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1338),
.B(n_1355),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1324),
.A2(n_809),
.B1(n_1054),
.B2(n_754),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1327),
.Y(n_1510)
);

CKINVDCx11_ASAP7_75t_R g1511 ( 
.A(n_1327),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1246),
.A2(n_754),
.B1(n_1027),
.B2(n_1324),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1327),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1246),
.A2(n_754),
.B1(n_1027),
.B2(n_1324),
.Y(n_1514)
);

OAI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1259),
.A2(n_1241),
.B1(n_1246),
.B2(n_1318),
.Y(n_1515)
);

AOI21xp33_ASAP7_75t_L g1516 ( 
.A1(n_1252),
.A2(n_1350),
.B(n_1333),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1250),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1324),
.A2(n_809),
.B1(n_1054),
.B2(n_754),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1246),
.A2(n_754),
.B1(n_1137),
.B2(n_1086),
.Y(n_1519)
);

BUFx4f_ASAP7_75t_SL g1520 ( 
.A(n_1320),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1447),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1504),
.B(n_1508),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1415),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1415),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1474),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1467),
.A2(n_1460),
.B(n_1477),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1476),
.B(n_1486),
.Y(n_1527)
);

AO21x2_ASAP7_75t_L g1528 ( 
.A1(n_1417),
.A2(n_1477),
.B(n_1455),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1486),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1499),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1499),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1460),
.A2(n_1411),
.B(n_1469),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1399),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1406),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1475),
.A2(n_1481),
.B1(n_1403),
.B2(n_1404),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1408),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1398),
.B(n_1515),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1515),
.B(n_1436),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1409),
.Y(n_1539)
);

BUFx2_ASAP7_75t_SL g1540 ( 
.A(n_1452),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1424),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1425),
.B(n_1487),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1488),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1433),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1439),
.B(n_1397),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1489),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1490),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1491),
.B(n_1494),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1411),
.A2(n_1472),
.B(n_1462),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1471),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1420),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1435),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1478),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1438),
.B(n_1426),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1497),
.Y(n_1555)
);

AO21x2_ASAP7_75t_L g1556 ( 
.A1(n_1417),
.A2(n_1455),
.B(n_1442),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1498),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1500),
.Y(n_1558)
);

OA21x2_ASAP7_75t_L g1559 ( 
.A1(n_1448),
.A2(n_1473),
.B(n_1516),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1462),
.A2(n_1448),
.B(n_1449),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1517),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1441),
.Y(n_1562)
);

AO21x2_ASAP7_75t_L g1563 ( 
.A1(n_1442),
.A2(n_1516),
.B(n_1404),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1492),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1445),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1446),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1492),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1470),
.Y(n_1568)
);

OR2x6_ASAP7_75t_L g1569 ( 
.A(n_1443),
.B(n_1481),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1492),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1422),
.B(n_1502),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1403),
.A2(n_1396),
.B(n_1419),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1449),
.A2(n_1465),
.B(n_1454),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1416),
.B(n_1437),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1470),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1470),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1450),
.Y(n_1577)
);

AO21x2_ASAP7_75t_L g1578 ( 
.A1(n_1454),
.A2(n_1463),
.B(n_1423),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1437),
.B(n_1440),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1407),
.B(n_1416),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1423),
.A2(n_1413),
.B(n_1464),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1407),
.B(n_1483),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1419),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1456),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1440),
.B(n_1427),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1479),
.A2(n_1509),
.B(n_1506),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1483),
.B(n_1495),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1456),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1468),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1463),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1512),
.A2(n_1514),
.B(n_1482),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1434),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1444),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1505),
.B(n_1501),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1444),
.Y(n_1595)
);

AO21x2_ASAP7_75t_L g1596 ( 
.A1(n_1495),
.A2(n_1519),
.B(n_1421),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1421),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1451),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1514),
.B(n_1428),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1466),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1400),
.B(n_1418),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1507),
.A2(n_1518),
.B1(n_1428),
.B2(n_1432),
.Y(n_1602)
);

INVx4_ASAP7_75t_L g1603 ( 
.A(n_1443),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1461),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1453),
.A2(n_1443),
.B(n_1452),
.Y(n_1605)
);

CKINVDCx14_ASAP7_75t_R g1606 ( 
.A(n_1493),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_SL g1607 ( 
.A(n_1457),
.B(n_1459),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1458),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1412),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1394),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1592),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1572),
.A2(n_1395),
.B(n_1429),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1592),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1537),
.A2(n_1485),
.B(n_1510),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1558),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1527),
.B(n_1402),
.Y(n_1616)
);

AND2x2_ASAP7_75t_SL g1617 ( 
.A(n_1587),
.B(n_1484),
.Y(n_1617)
);

AO32x2_ASAP7_75t_L g1618 ( 
.A1(n_1551),
.A2(n_1520),
.A3(n_1402),
.B1(n_1431),
.B2(n_1414),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1529),
.B(n_1480),
.Y(n_1619)
);

NAND4xp25_ASAP7_75t_L g1620 ( 
.A(n_1535),
.B(n_1511),
.C(n_1503),
.D(n_1496),
.Y(n_1620)
);

NAND3xp33_ASAP7_75t_L g1621 ( 
.A(n_1583),
.B(n_1401),
.C(n_1513),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1577),
.B(n_1480),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1558),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1583),
.A2(n_1430),
.B(n_1405),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1598),
.B(n_1410),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1558),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1538),
.B(n_1588),
.C(n_1584),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1581),
.A2(n_1580),
.B(n_1582),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1554),
.B(n_1522),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1598),
.B(n_1600),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1581),
.A2(n_1580),
.B(n_1582),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1533),
.B(n_1534),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1542),
.B(n_1548),
.Y(n_1633)
);

A2O1A1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1587),
.A2(n_1586),
.B(n_1574),
.C(n_1599),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1563),
.A2(n_1556),
.B(n_1578),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1530),
.B(n_1531),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1563),
.A2(n_1556),
.B(n_1578),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1571),
.B(n_1601),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_SL g1639 ( 
.A1(n_1585),
.A2(n_1607),
.B(n_1589),
.Y(n_1639)
);

AOI22x1_ASAP7_75t_SL g1640 ( 
.A1(n_1525),
.A2(n_1608),
.B1(n_1606),
.B2(n_1610),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1588),
.B(n_1574),
.C(n_1589),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1536),
.B(n_1539),
.Y(n_1642)
);

OAI211xp5_ASAP7_75t_L g1643 ( 
.A1(n_1589),
.A2(n_1550),
.B(n_1579),
.C(n_1595),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1602),
.A2(n_1593),
.B(n_1595),
.C(n_1597),
.Y(n_1644)
);

AO32x2_ASAP7_75t_L g1645 ( 
.A1(n_1551),
.A2(n_1603),
.A3(n_1544),
.B1(n_1545),
.B2(n_1559),
.Y(n_1645)
);

NOR2x1_ASAP7_75t_SL g1646 ( 
.A(n_1569),
.B(n_1540),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1525),
.B(n_1604),
.Y(n_1647)
);

AOI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1597),
.A2(n_1593),
.B1(n_1523),
.B2(n_1524),
.C(n_1555),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1594),
.B(n_1609),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1573),
.A2(n_1525),
.B(n_1560),
.C(n_1590),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1541),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1525),
.B(n_1604),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1591),
.A2(n_1569),
.B1(n_1608),
.B2(n_1559),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1591),
.A2(n_1569),
.B1(n_1608),
.B2(n_1559),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1543),
.Y(n_1655)
);

NAND4xp25_ASAP7_75t_L g1656 ( 
.A(n_1550),
.B(n_1575),
.C(n_1568),
.D(n_1576),
.Y(n_1656)
);

AO32x2_ASAP7_75t_L g1657 ( 
.A1(n_1603),
.A2(n_1544),
.A3(n_1559),
.B1(n_1596),
.B2(n_1591),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1592),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1549),
.A2(n_1526),
.B(n_1532),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1546),
.Y(n_1660)
);

A2O1A1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1590),
.A2(n_1532),
.B(n_1526),
.C(n_1550),
.Y(n_1661)
);

AO32x2_ASAP7_75t_L g1662 ( 
.A1(n_1603),
.A2(n_1544),
.A3(n_1596),
.B1(n_1591),
.B2(n_1552),
.Y(n_1662)
);

CKINVDCx8_ASAP7_75t_R g1663 ( 
.A(n_1540),
.Y(n_1663)
);

AOI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1547),
.A2(n_1557),
.B1(n_1561),
.B2(n_1562),
.C(n_1596),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1628),
.A2(n_1528),
.B1(n_1566),
.B2(n_1565),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1633),
.B(n_1528),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1646),
.B(n_1564),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1615),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1623),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1626),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1639),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1636),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1635),
.B(n_1550),
.Y(n_1673)
);

INVxp67_ASAP7_75t_SL g1674 ( 
.A(n_1637),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1659),
.B(n_1638),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1645),
.B(n_1521),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1645),
.B(n_1521),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1664),
.B(n_1568),
.Y(n_1678)
);

NOR2x1_ASAP7_75t_L g1679 ( 
.A(n_1656),
.B(n_1568),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1651),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1655),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1645),
.B(n_1521),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1657),
.B(n_1521),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1660),
.B(n_1650),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1657),
.B(n_1567),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1662),
.Y(n_1686)
);

BUFx2_ASAP7_75t_SL g1687 ( 
.A(n_1663),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1632),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1642),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1662),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1662),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1647),
.Y(n_1692)
);

INVxp67_ASAP7_75t_L g1693 ( 
.A(n_1619),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1661),
.B(n_1570),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1648),
.B(n_1575),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1680),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1683),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1672),
.B(n_1629),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1680),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1678),
.A2(n_1695),
.B(n_1674),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1666),
.B(n_1653),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1671),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1681),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1666),
.B(n_1654),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1671),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1692),
.B(n_1630),
.Y(n_1706)
);

OAI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1665),
.A2(n_1628),
.B1(n_1631),
.B2(n_1634),
.C(n_1627),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1683),
.Y(n_1708)
);

NOR3xp33_ASAP7_75t_SL g1709 ( 
.A(n_1673),
.B(n_1620),
.C(n_1621),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1672),
.B(n_1654),
.Y(n_1710)
);

NOR3xp33_ASAP7_75t_L g1711 ( 
.A(n_1673),
.B(n_1621),
.C(n_1620),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1675),
.B(n_1630),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1675),
.B(n_1652),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1668),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1665),
.A2(n_1631),
.B1(n_1627),
.B2(n_1643),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1684),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1671),
.Y(n_1717)
);

AO21x2_ASAP7_75t_L g1718 ( 
.A1(n_1674),
.A2(n_1641),
.B(n_1644),
.Y(n_1718)
);

INVx5_ASAP7_75t_L g1719 ( 
.A(n_1676),
.Y(n_1719)
);

NAND2x1_ASAP7_75t_L g1720 ( 
.A(n_1679),
.B(n_1625),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1695),
.A2(n_1641),
.B1(n_1617),
.B2(n_1612),
.Y(n_1721)
);

INVx4_ASAP7_75t_L g1722 ( 
.A(n_1667),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1668),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1669),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1693),
.B(n_1658),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1679),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1684),
.B(n_1616),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1670),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1686),
.A2(n_1624),
.B1(n_1612),
.B2(n_1553),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1719),
.B(n_1676),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1714),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1719),
.B(n_1677),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1716),
.B(n_1678),
.Y(n_1733)
);

INVx4_ASAP7_75t_L g1734 ( 
.A(n_1717),
.Y(n_1734)
);

INVx4_ASAP7_75t_L g1735 ( 
.A(n_1717),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1698),
.B(n_1688),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1725),
.B(n_1640),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1719),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1714),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1712),
.B(n_1713),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1723),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1696),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1697),
.B(n_1677),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1696),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1697),
.B(n_1682),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1698),
.B(n_1689),
.Y(n_1746)
);

NOR2x1p5_ASAP7_75t_L g1747 ( 
.A(n_1720),
.B(n_1622),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1722),
.B(n_1694),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1708),
.B(n_1685),
.Y(n_1749)
);

INVx3_ASAP7_75t_SL g1750 ( 
.A(n_1717),
.Y(n_1750)
);

NOR2x1_ASAP7_75t_L g1751 ( 
.A(n_1720),
.B(n_1687),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1700),
.B(n_1685),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1723),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1724),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1699),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1724),
.Y(n_1756)
);

NOR2x1_ASAP7_75t_L g1757 ( 
.A(n_1726),
.B(n_1687),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1722),
.B(n_1694),
.Y(n_1758)
);

OR2x6_ASAP7_75t_L g1759 ( 
.A(n_1701),
.B(n_1605),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1749),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1748),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1731),
.Y(n_1762)
);

AOI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1752),
.A2(n_1707),
.B1(n_1711),
.B2(n_1710),
.C(n_1709),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1740),
.B(n_1702),
.Y(n_1764)
);

OR2x6_ASAP7_75t_L g1765 ( 
.A(n_1738),
.B(n_1605),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1740),
.B(n_1702),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1749),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1731),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1742),
.B(n_1728),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1739),
.Y(n_1770)
);

INVxp67_ASAP7_75t_L g1771 ( 
.A(n_1742),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1749),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1743),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1739),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1743),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1752),
.A2(n_1718),
.B1(n_1715),
.B2(n_1701),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1744),
.B(n_1728),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1741),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1743),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1744),
.B(n_1703),
.Y(n_1780)
);

OR2x2_ASAP7_75t_SL g1781 ( 
.A(n_1733),
.B(n_1717),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1741),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1753),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1755),
.B(n_1703),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1753),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1751),
.B(n_1705),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1751),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1747),
.B(n_1705),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1754),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1737),
.B(n_1727),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1757),
.B(n_1717),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1754),
.Y(n_1792)
);

NAND2x1p5_ASAP7_75t_L g1793 ( 
.A(n_1757),
.B(n_1717),
.Y(n_1793)
);

OR2x6_ASAP7_75t_L g1794 ( 
.A(n_1738),
.B(n_1686),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1747),
.B(n_1748),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1736),
.B(n_1710),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1748),
.B(n_1721),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1748),
.B(n_1722),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1745),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1750),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1756),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1758),
.B(n_1706),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1756),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1745),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1762),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1762),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1768),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1764),
.B(n_1750),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1763),
.B(n_1733),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1800),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1768),
.Y(n_1811)
);

NAND2x1_ASAP7_75t_L g1812 ( 
.A(n_1787),
.B(n_1738),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1764),
.B(n_1750),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1760),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1770),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1781),
.Y(n_1816)
);

NOR2x1_ASAP7_75t_L g1817 ( 
.A(n_1791),
.B(n_1734),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1770),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1761),
.B(n_1795),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1766),
.B(n_1758),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1760),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1774),
.Y(n_1822)
);

AND2x2_ASAP7_75t_SL g1823 ( 
.A(n_1776),
.B(n_1734),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1774),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1778),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1766),
.B(n_1758),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1778),
.Y(n_1827)
);

NAND2xp67_ASAP7_75t_L g1828 ( 
.A(n_1788),
.B(n_1730),
.Y(n_1828)
);

INVx1_ASAP7_75t_SL g1829 ( 
.A(n_1800),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1760),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1802),
.B(n_1758),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1790),
.B(n_1727),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1782),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1796),
.B(n_1746),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1802),
.B(n_1734),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1795),
.B(n_1734),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1782),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1761),
.B(n_1787),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1786),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1771),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1797),
.B(n_1735),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1805),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1805),
.Y(n_1843)
);

AOI21xp33_ASAP7_75t_L g1844 ( 
.A1(n_1809),
.A2(n_1763),
.B(n_1794),
.Y(n_1844)
);

OAI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1816),
.A2(n_1715),
.B1(n_1721),
.B2(n_1704),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1832),
.B(n_1771),
.Y(n_1846)
);

NAND2x1_ASAP7_75t_L g1847 ( 
.A(n_1816),
.B(n_1761),
.Y(n_1847)
);

AND3x2_ASAP7_75t_L g1848 ( 
.A(n_1840),
.B(n_1614),
.C(n_1786),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1823),
.A2(n_1787),
.B(n_1793),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1823),
.A2(n_1718),
.B1(n_1729),
.B2(n_1759),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_R g1851 ( 
.A(n_1810),
.B(n_1761),
.Y(n_1851)
);

OAI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1823),
.A2(n_1793),
.B(n_1788),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1806),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1806),
.Y(n_1854)
);

NAND3xp33_ASAP7_75t_L g1855 ( 
.A(n_1841),
.B(n_1785),
.C(n_1783),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1807),
.Y(n_1856)
);

NOR4xp25_ASAP7_75t_SL g1857 ( 
.A(n_1807),
.B(n_1781),
.C(n_1803),
.D(n_1801),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1808),
.B(n_1793),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1829),
.B(n_1796),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1829),
.B(n_1839),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1820),
.B(n_1798),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1839),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1808),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1811),
.Y(n_1864)
);

INVxp67_ASAP7_75t_SL g1865 ( 
.A(n_1814),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1820),
.A2(n_1767),
.B1(n_1772),
.B2(n_1732),
.Y(n_1866)
);

NOR2x1_ASAP7_75t_L g1867 ( 
.A(n_1812),
.B(n_1735),
.Y(n_1867)
);

OAI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1834),
.A2(n_1794),
.B1(n_1765),
.B2(n_1614),
.C(n_1690),
.Y(n_1868)
);

OAI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1834),
.A2(n_1794),
.B1(n_1765),
.B2(n_1691),
.C(n_1690),
.Y(n_1869)
);

NOR2x1_ASAP7_75t_L g1870 ( 
.A(n_1860),
.B(n_1847),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1859),
.B(n_1767),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1857),
.A2(n_1812),
.B(n_1838),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1865),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1865),
.Y(n_1874)
);

INVx1_ASAP7_75t_SL g1875 ( 
.A(n_1851),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1862),
.B(n_1826),
.Y(n_1876)
);

NAND2xp33_ASAP7_75t_L g1877 ( 
.A(n_1863),
.B(n_1817),
.Y(n_1877)
);

O2A1O1Ixp33_ASAP7_75t_L g1878 ( 
.A1(n_1844),
.A2(n_1818),
.B(n_1837),
.C(n_1811),
.Y(n_1878)
);

NOR3xp33_ASAP7_75t_L g1879 ( 
.A(n_1862),
.B(n_1821),
.C(n_1814),
.Y(n_1879)
);

OAI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1850),
.A2(n_1704),
.B1(n_1794),
.B2(n_1759),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1861),
.B(n_1826),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1846),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1842),
.Y(n_1883)
);

INVxp67_ASAP7_75t_SL g1884 ( 
.A(n_1867),
.Y(n_1884)
);

INVx1_ASAP7_75t_SL g1885 ( 
.A(n_1848),
.Y(n_1885)
);

OAI211xp5_ASAP7_75t_L g1886 ( 
.A1(n_1852),
.A2(n_1817),
.B(n_1837),
.C(n_1818),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1843),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1853),
.Y(n_1888)
);

AOI32xp33_ASAP7_75t_L g1889 ( 
.A1(n_1845),
.A2(n_1868),
.A3(n_1869),
.B1(n_1848),
.B2(n_1866),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1854),
.Y(n_1890)
);

AOI211xp5_ASAP7_75t_L g1891 ( 
.A1(n_1849),
.A2(n_1822),
.B(n_1815),
.C(n_1824),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1881),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1873),
.Y(n_1893)
);

NOR4xp25_ASAP7_75t_L g1894 ( 
.A(n_1878),
.B(n_1864),
.C(n_1856),
.D(n_1855),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1876),
.B(n_1814),
.Y(n_1895)
);

CKINVDCx14_ASAP7_75t_R g1896 ( 
.A(n_1876),
.Y(n_1896)
);

OAI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1872),
.A2(n_1838),
.B(n_1858),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1885),
.A2(n_1821),
.B1(n_1830),
.B2(n_1833),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1882),
.B(n_1879),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1875),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1874),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1870),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1890),
.B(n_1819),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1871),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1883),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1904),
.Y(n_1906)
);

AOI21xp33_ASAP7_75t_L g1907 ( 
.A1(n_1904),
.A2(n_1878),
.B(n_1887),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1895),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1900),
.B(n_1884),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1894),
.A2(n_1872),
.B(n_1877),
.Y(n_1910)
);

AND4x1_ASAP7_75t_L g1911 ( 
.A(n_1903),
.B(n_1891),
.C(n_1888),
.D(n_1813),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1896),
.B(n_1889),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1899),
.Y(n_1913)
);

NOR4xp25_ASAP7_75t_L g1914 ( 
.A(n_1902),
.B(n_1886),
.C(n_1880),
.D(n_1821),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1892),
.B(n_1767),
.Y(n_1915)
);

NAND4xp25_ASAP7_75t_L g1916 ( 
.A(n_1903),
.B(n_1886),
.C(n_1819),
.D(n_1838),
.Y(n_1916)
);

OAI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1897),
.A2(n_1838),
.B(n_1819),
.Y(n_1917)
);

OAI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1914),
.A2(n_1898),
.B1(n_1902),
.B2(n_1893),
.C(n_1901),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1907),
.A2(n_1898),
.B1(n_1893),
.B2(n_1905),
.C(n_1830),
.Y(n_1919)
);

OAI211xp5_ASAP7_75t_SL g1920 ( 
.A1(n_1910),
.A2(n_1912),
.B(n_1909),
.C(n_1917),
.Y(n_1920)
);

O2A1O1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1913),
.A2(n_1794),
.B(n_1822),
.C(n_1833),
.Y(n_1921)
);

OAI211xp5_ASAP7_75t_L g1922 ( 
.A1(n_1916),
.A2(n_1836),
.B(n_1813),
.C(n_1835),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1915),
.B(n_1772),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1911),
.B(n_1819),
.Y(n_1924)
);

OAI321xp33_ASAP7_75t_L g1925 ( 
.A1(n_1906),
.A2(n_1830),
.A3(n_1836),
.B1(n_1794),
.B2(n_1815),
.C(n_1825),
.Y(n_1925)
);

NOR2x1_ASAP7_75t_L g1926 ( 
.A(n_1908),
.B(n_1824),
.Y(n_1926)
);

NOR2xp67_ASAP7_75t_L g1927 ( 
.A(n_1925),
.B(n_1913),
.Y(n_1927)
);

O2A1O1Ixp5_ASAP7_75t_SL g1928 ( 
.A1(n_1924),
.A2(n_1825),
.B(n_1827),
.C(n_1785),
.Y(n_1928)
);

OAI21xp33_ASAP7_75t_L g1929 ( 
.A1(n_1920),
.A2(n_1828),
.B(n_1835),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1923),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1919),
.B(n_1735),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1918),
.A2(n_1827),
.B1(n_1772),
.B2(n_1773),
.C(n_1804),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1926),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1922),
.B(n_1831),
.Y(n_1934)
);

OAI211xp5_ASAP7_75t_L g1935 ( 
.A1(n_1921),
.A2(n_1735),
.B(n_1831),
.C(n_1798),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1927),
.B(n_1828),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1933),
.B(n_1783),
.Y(n_1937)
);

OAI211xp5_ASAP7_75t_SL g1938 ( 
.A1(n_1929),
.A2(n_1804),
.B(n_1773),
.C(n_1775),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1930),
.B(n_1773),
.Y(n_1939)
);

NOR2x1_ASAP7_75t_L g1940 ( 
.A(n_1931),
.B(n_1789),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1934),
.B(n_1775),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1939),
.B(n_1935),
.Y(n_1942)
);

NAND2x1p5_ASAP7_75t_L g1943 ( 
.A(n_1937),
.B(n_1940),
.Y(n_1943)
);

OAI211xp5_ASAP7_75t_L g1944 ( 
.A1(n_1936),
.A2(n_1932),
.B(n_1938),
.C(n_1941),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1942),
.B(n_1775),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1945),
.Y(n_1946)
);

AOI311xp33_ASAP7_75t_L g1947 ( 
.A1(n_1946),
.A2(n_1944),
.A3(n_1943),
.B(n_1928),
.C(n_1789),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1946),
.A2(n_1804),
.B1(n_1779),
.B2(n_1799),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1948),
.A2(n_1784),
.B(n_1780),
.Y(n_1949)
);

OAI22x1_ASAP7_75t_L g1950 ( 
.A1(n_1947),
.A2(n_1799),
.B1(n_1779),
.B2(n_1649),
.Y(n_1950)
);

AO22x2_ASAP7_75t_L g1951 ( 
.A1(n_1950),
.A2(n_1779),
.B1(n_1799),
.B2(n_1803),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1949),
.A2(n_1784),
.B(n_1780),
.Y(n_1952)
);

OAI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1952),
.A2(n_1624),
.B(n_1769),
.Y(n_1953)
);

OAI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1953),
.A2(n_1951),
.B1(n_1769),
.B2(n_1777),
.Y(n_1954)
);

CKINVDCx20_ASAP7_75t_R g1955 ( 
.A(n_1954),
.Y(n_1955)
);

AOI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1955),
.A2(n_1801),
.B1(n_1792),
.B2(n_1777),
.C(n_1755),
.Y(n_1956)
);

AOI211xp5_ASAP7_75t_L g1957 ( 
.A1(n_1956),
.A2(n_1618),
.B(n_1611),
.C(n_1613),
.Y(n_1957)
);


endmodule