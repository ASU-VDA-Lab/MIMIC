module fake_jpeg_18465_n_175 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_127;
wire n_76;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_7),
.B(n_2),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_20),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_22),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_33),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_0),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_0),
.B(n_1),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_1),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_82),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_83),
.B1(n_60),
.B2(n_70),
.Y(n_109)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_84),
.B1(n_64),
.B2(n_71),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_97),
.B1(n_85),
.B2(n_98),
.Y(n_122)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_91),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_86),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_57),
.C(n_65),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_125),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_123),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_97),
.B1(n_62),
.B2(n_93),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_122),
.B1(n_128),
.B2(n_129),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_92),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_56),
.Y(n_134)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_95),
.B1(n_79),
.B2(n_58),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_72),
.B1(n_78),
.B2(n_66),
.Y(n_129)
);

OAI22x1_ASAP7_75t_SL g130 ( 
.A1(n_118),
.A2(n_58),
.B1(n_79),
.B2(n_77),
.Y(n_130)
);

OAI22x1_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_137),
.B1(n_4),
.B2(n_5),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_67),
.B(n_59),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_134),
.B(n_3),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_73),
.B1(n_55),
.B2(n_61),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_139),
.B1(n_6),
.B2(n_9),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_142),
.Y(n_151)
);

AO21x2_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_63),
.B(n_77),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_80),
.B1(n_75),
.B2(n_74),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_143),
.Y(n_145)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_68),
.C(n_76),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_116),
.B1(n_76),
.B2(n_51),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_150),
.B1(n_137),
.B2(n_9),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_149),
.B(n_6),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_51),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_153),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_158),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_137),
.B1(n_15),
.B2(n_18),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_159),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_162),
.B1(n_157),
.B2(n_154),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_144),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_151),
.C(n_157),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_161),
.B1(n_145),
.B2(n_26),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_14),
.B(n_24),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_170)
);

O2A1O1Ixp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_34),
.B(n_35),
.C(n_38),
.Y(n_171)
);

OAI21x1_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_43),
.B(n_45),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_46),
.B(n_47),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_48),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_50),
.B(n_137),
.Y(n_175)
);


endmodule