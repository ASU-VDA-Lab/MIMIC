module real_jpeg_3705_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_0),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_3),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_3),
.A2(n_32),
.B1(n_38),
.B2(n_114),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_114),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_3),
.A2(n_75),
.B1(n_76),
.B2(n_114),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_4),
.A2(n_27),
.B1(n_29),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_4),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_4),
.A2(n_32),
.B1(n_38),
.B2(n_84),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_84),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_4),
.A2(n_75),
.B1(n_76),
.B2(n_84),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_5),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_26),
.B1(n_32),
.B2(n_38),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_5),
.A2(n_26),
.B1(n_75),
.B2(n_76),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_6),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_136),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_6),
.A2(n_32),
.B1(n_38),
.B2(n_136),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_6),
.A2(n_75),
.B1(n_76),
.B2(n_136),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_32),
.B1(n_38),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_7),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_67),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_7),
.A2(n_67),
.B1(n_75),
.B2(n_76),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_8),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_8),
.A2(n_32),
.B1(n_38),
.B2(n_175),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_175),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_8),
.A2(n_75),
.B1(n_76),
.B2(n_175),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_9),
.Y(n_346)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_20),
.B(n_344),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g345 ( 
.A(n_13),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_14),
.A2(n_32),
.B1(n_38),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_64),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_14),
.A2(n_64),
.B1(n_75),
.B2(n_76),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_16),
.B(n_42),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_16),
.B(n_57),
.C(n_59),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_16),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_16),
.B(n_56),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_16),
.B(n_72),
.C(n_75),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_16),
.A2(n_58),
.B1(n_59),
.B2(n_210),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_16),
.B(n_107),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_16),
.B(n_93),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_16),
.A2(n_32),
.B1(n_38),
.B2(n_210),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_17),
.A2(n_27),
.B1(n_29),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_17),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_17),
.A2(n_41),
.B1(n_75),
.B2(n_76),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_17),
.A2(n_32),
.B1(n_38),
.B2(n_41),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_46),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_44),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_43),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_23),
.B(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_24),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_24),
.B(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_40),
.B2(n_42),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_25),
.A2(n_30),
.B1(n_42),
.B2(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_27),
.A2(n_85),
.B(n_210),
.C(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_27),
.B(n_210),
.Y(n_211)
);

AOI32xp33_ASAP7_75t_L g222 ( 
.A1(n_27),
.A2(n_35),
.A3(n_38),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_40),
.B(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_30),
.B(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_30),
.A2(n_42),
.B1(n_135),
.B2(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_31),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_31),
.A2(n_83),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_31),
.B(n_113),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_31),
.A2(n_85),
.B1(n_86),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_31),
.A2(n_111),
.B(n_296),
.Y(n_295)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_31)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_38),
.B1(n_57),
.B2(n_61),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_32),
.B(n_200),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_SL g224 ( 
.A(n_32),
.B(n_36),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

OAI21x1_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_339),
.B(n_341),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_327),
.B(n_338),
.Y(n_47)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_151),
.B(n_324),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_139),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_115),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_51),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_51),
.B(n_115),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_51),
.B(n_140),
.Y(n_326)
);

FAx1_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_80),
.CI(n_96),
.CON(n_51),
.SN(n_51)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_52),
.A2(n_53),
.B(n_68),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_68),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_65),
.B1(n_66),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_54),
.A2(n_63),
.B1(n_65),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_54),
.A2(n_65),
.B1(n_90),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_54),
.A2(n_65),
.B1(n_183),
.B2(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_54),
.A2(n_275),
.B(n_276),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_54),
.A2(n_214),
.B(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_55),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_55),
.A2(n_56),
.B(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_56),
.B(n_172),
.Y(n_276)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_59),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_59),
.B(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_65),
.A2(n_132),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_65),
.A2(n_171),
.B(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_69),
.A2(n_74),
.B1(n_78),
.B2(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_69),
.A2(n_195),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_69),
.A2(n_74),
.B1(n_193),
.B2(n_243),
.Y(n_277)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_70),
.A2(n_93),
.B1(n_101),
.B2(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_70),
.A2(n_93),
.B1(n_130),
.B2(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_70),
.A2(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_70),
.B(n_196),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_74),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_74),
.A2(n_217),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_75),
.B(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_87),
.B2(n_95),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_81),
.A2(n_82),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g150 ( 
.A(n_82),
.B(n_88),
.C(n_92),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_82),
.B(n_143),
.C(n_150),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_134),
.B(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_91),
.A2(n_92),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_92),
.B(n_144),
.C(n_148),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_93),
.B(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_103),
.B(n_110),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_98),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_99),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_103),
.B1(n_110),
.B2(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_107),
.B(n_108),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_104),
.A2(n_107),
.B1(n_127),
.B2(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_104),
.A2(n_210),
.B(n_237),
.Y(n_257)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_105),
.A2(n_106),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_105),
.B(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_105),
.A2(n_106),
.B1(n_190),
.B2(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_105),
.A2(n_235),
.B(n_236),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_105),
.A2(n_106),
.B1(n_235),
.B2(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_106),
.A2(n_189),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_106),
.B(n_204),
.Y(n_237)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_107),
.A2(n_203),
.B(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_131),
.C(n_133),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_124),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_125),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_133),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_138),
.B(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_139),
.A2(n_325),
.B(n_326),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_145),
.Y(n_333)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_149),
.Y(n_331)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_176),
.B(n_323),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_153),
.B(n_156),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_162),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_157),
.B(n_160),
.Y(n_321)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_162),
.B(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_169),
.C(n_173),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_163),
.A2(n_164),
.B1(n_311),
.B2(n_313),
.Y(n_310)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_165),
.B(n_167),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_168),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_173),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_174),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_318),
.B(n_322),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_287),
.B(n_315),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_229),
.B(n_286),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_205),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_180),
.B(n_205),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_191),
.C(n_197),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_181),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_185),
.C(n_188),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_191),
.B(n_197),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_219),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_206),
.B(n_220),
.C(n_228),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_212),
.B2(n_218),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_207),
.B(n_213),
.C(n_215),
.Y(n_300)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_228),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_221),
.B(n_226),
.Y(n_291)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_281),
.B(n_285),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_270),
.B(n_280),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_252),
.B(n_269),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_246),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_246),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_238),
.B1(n_244),
.B2(n_245),
.Y(n_233)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_241),
.C(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_263),
.B(n_268),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_258),
.B(n_262),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_261),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_260),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_266),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_272),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_277),
.C(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_302),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_301),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_301),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_298),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_299),
.C(n_300),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_293),
.C(n_297),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_297),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_314),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_314),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_308),
.C(n_310),
.Y(n_319)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_311),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_320),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_337),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_337),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_336),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_334),
.C(n_336),
.Y(n_340)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_340),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);


endmodule