module fake_jpeg_14072_n_111 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_2),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_51),
.Y(n_55)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_49),
.B1(n_38),
.B2(n_41),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_38),
.B1(n_37),
.B2(n_42),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_3),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_1),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_78),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_77),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_63),
.B1(n_56),
.B2(n_6),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_4),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_4),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_22),
.B(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_5),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_85),
.B(n_73),
.Y(n_99)
);

AO22x1_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_15),
.B1(n_16),
.B2(n_20),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_96),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_69),
.B(n_25),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_94),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_70),
.B(n_26),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_86),
.C(n_84),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_91),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_108),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_103),
.A3(n_105),
.B1(n_97),
.B2(n_89),
.C1(n_102),
.C2(n_83),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_88),
.Y(n_111)
);


endmodule