module real_aes_6208_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_746;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g571 ( .A1(n_0), .A2(n_171), .B(n_572), .C(n_575), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_1), .B(n_517), .Y(n_576) );
INVx1_ASAP7_75t_L g117 ( .A(n_2), .Y(n_117) );
INVx1_ASAP7_75t_L g205 ( .A(n_3), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_4), .B(n_163), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_5), .A2(n_486), .B(n_511), .Y(n_510) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_6), .A2(n_148), .B(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_7), .A2(n_37), .B1(n_157), .B2(n_235), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_8), .A2(n_106), .B1(n_119), .B2(n_769), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_9), .B(n_148), .Y(n_174) );
AND2x6_ASAP7_75t_L g172 ( .A(n_10), .B(n_173), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_11), .A2(n_172), .B(n_476), .C(n_478), .Y(n_475) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_12), .A2(n_457), .B1(n_750), .B2(n_751), .C1(n_760), .C2(n_764), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_13), .B(n_38), .Y(n_118) );
INVx1_ASAP7_75t_L g153 ( .A(n_14), .Y(n_153) );
INVx1_ASAP7_75t_L g198 ( .A(n_15), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_16), .B(n_161), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_17), .B(n_163), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_18), .B(n_149), .Y(n_210) );
AO32x2_ASAP7_75t_L g232 ( .A1(n_19), .A2(n_148), .A3(n_178), .B1(n_189), .B2(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_20), .B(n_157), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_21), .B(n_149), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_22), .A2(n_57), .B1(n_157), .B2(n_235), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g257 ( .A1(n_23), .A2(n_85), .B1(n_157), .B2(n_161), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_24), .B(n_157), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_25), .A2(n_189), .B(n_476), .C(n_537), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_26), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_26), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_27), .A2(n_189), .B(n_476), .C(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_28), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_29), .B(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_30), .A2(n_486), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_31), .B(n_191), .Y(n_229) );
INVx2_ASAP7_75t_L g159 ( .A(n_32), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_33), .A2(n_488), .B(n_496), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_34), .B(n_157), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_35), .B(n_191), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_36), .B(n_243), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_39), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_40), .B(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_41), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_42), .A2(n_81), .B1(n_756), .B2(n_757), .Y(n_755) );
CKINVDCx16_ASAP7_75t_R g757 ( .A(n_42), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_43), .B(n_163), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_44), .B(n_486), .Y(n_503) );
OAI22xp5_ASAP7_75t_SL g137 ( .A1(n_45), .A2(n_82), .B1(n_138), .B2(n_139), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_45), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_46), .A2(n_488), .B(n_490), .C(n_496), .Y(n_487) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_47), .A2(n_755), .B1(n_758), .B2(n_759), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_47), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_48), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g573 ( .A(n_49), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_50), .A2(n_94), .B1(n_235), .B2(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g491 ( .A(n_51), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_52), .B(n_157), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_53), .B(n_157), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_54), .A2(n_128), .B1(n_129), .B2(n_132), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_54), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_55), .B(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_56), .B(n_169), .Y(n_168) );
AOI22xp33_ASAP7_75t_SL g214 ( .A1(n_58), .A2(n_62), .B1(n_157), .B2(n_161), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_59), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_60), .B(n_157), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_61), .B(n_157), .Y(n_240) );
INVx1_ASAP7_75t_L g173 ( .A(n_63), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_64), .B(n_486), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_65), .B(n_517), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_66), .A2(n_169), .B(n_201), .C(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_67), .B(n_157), .Y(n_206) );
INVx1_ASAP7_75t_L g152 ( .A(n_68), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_69), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_70), .B(n_163), .Y(n_527) );
AO32x2_ASAP7_75t_L g253 ( .A1(n_71), .A2(n_148), .A3(n_189), .B1(n_254), .B2(n_258), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_72), .B(n_164), .Y(n_479) );
INVx1_ASAP7_75t_L g184 ( .A(n_73), .Y(n_184) );
INVx1_ASAP7_75t_L g224 ( .A(n_74), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g570 ( .A(n_75), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_76), .B(n_493), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_77), .A2(n_476), .B(n_496), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_78), .B(n_161), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_79), .Y(n_512) );
INVx1_ASAP7_75t_L g112 ( .A(n_80), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_81), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_82), .Y(n_139) );
OAI22xp5_ASAP7_75t_SL g458 ( .A1(n_82), .A2(n_139), .B1(n_140), .B2(n_450), .Y(n_458) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_83), .A2(n_90), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_83), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_84), .B(n_492), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_86), .B(n_235), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_87), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_88), .B(n_161), .Y(n_228) );
INVx2_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_90), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_91), .B(n_188), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_92), .B(n_161), .Y(n_160) );
OR2x2_ASAP7_75t_L g114 ( .A(n_93), .B(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g461 ( .A(n_93), .B(n_116), .Y(n_461) );
INVx2_ASAP7_75t_L g749 ( .A(n_93), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_95), .A2(n_104), .B1(n_161), .B2(n_162), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_96), .B(n_486), .Y(n_523) );
INVx1_ASAP7_75t_L g526 ( .A(n_97), .Y(n_526) );
INVxp67_ASAP7_75t_L g515 ( .A(n_98), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_99), .B(n_161), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g472 ( .A(n_101), .Y(n_472) );
INVx1_ASAP7_75t_L g550 ( .A(n_102), .Y(n_550) );
AND2x2_ASAP7_75t_L g498 ( .A(n_103), .B(n_191), .Y(n_498) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx6p67_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g770 ( .A(n_109), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_113), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_SL g125 ( .A(n_114), .Y(n_125) );
INVx2_ASAP7_75t_L g454 ( .A(n_114), .Y(n_454) );
NOR2x2_ASAP7_75t_L g766 ( .A(n_115), .B(n_749), .Y(n_766) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g748 ( .A(n_116), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
OA21x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_124), .B(n_455), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g768 ( .A(n_122), .Y(n_768) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B(n_451), .Y(n_124) );
XOR2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_133), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_131), .B(n_215), .Y(n_554) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B1(n_140), .B2(n_450), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g450 ( .A(n_140), .Y(n_450) );
NAND2x1p5_ASAP7_75t_L g140 ( .A(n_141), .B(n_374), .Y(n_140) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_332), .Y(n_141) );
NOR4xp25_ASAP7_75t_L g142 ( .A(n_143), .B(n_272), .C(n_308), .D(n_322), .Y(n_142) );
OAI221xp5_ASAP7_75t_SL g143 ( .A1(n_144), .A2(n_216), .B1(n_248), .B2(n_259), .C(n_263), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_144), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_192), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_175), .Y(n_146) );
AND2x2_ASAP7_75t_L g269 ( .A(n_147), .B(n_176), .Y(n_269) );
INVx3_ASAP7_75t_L g277 ( .A(n_147), .Y(n_277) );
AND2x2_ASAP7_75t_L g331 ( .A(n_147), .B(n_195), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_147), .B(n_194), .Y(n_367) );
AND2x2_ASAP7_75t_L g425 ( .A(n_147), .B(n_287), .Y(n_425) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_154), .B(n_174), .Y(n_147) );
INVx4_ASAP7_75t_L g215 ( .A(n_148), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_148), .A2(n_503), .B(n_504), .Y(n_502) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_148), .Y(n_509) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_150), .B(n_151), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_166), .B(n_172), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_160), .B(n_163), .Y(n_155) );
INVx3_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_157), .Y(n_552) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g235 ( .A(n_158), .Y(n_235) );
BUFx3_ASAP7_75t_L g256 ( .A(n_158), .Y(n_256) );
AND2x6_ASAP7_75t_L g476 ( .A(n_158), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g162 ( .A(n_159), .Y(n_162) );
INVx1_ASAP7_75t_L g170 ( .A(n_159), .Y(n_170) );
INVx2_ASAP7_75t_L g199 ( .A(n_161), .Y(n_199) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g171 ( .A(n_163), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_163), .A2(n_181), .B(n_182), .Y(n_180) );
O2A1O1Ixp5_ASAP7_75t_SL g222 ( .A1(n_163), .A2(n_223), .B(n_224), .C(n_225), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_163), .B(n_515), .Y(n_514) );
INVx5_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g254 ( .A1(n_164), .A2(n_188), .B1(n_255), .B2(n_257), .Y(n_254) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
INVx1_ASAP7_75t_L g243 ( .A(n_165), .Y(n_243) );
AND2x2_ASAP7_75t_L g474 ( .A(n_165), .B(n_170), .Y(n_474) );
INVx1_ASAP7_75t_L g477 ( .A(n_165), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_171), .Y(n_166) );
INVx2_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_171), .A2(n_185), .B(n_205), .C(n_206), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_171), .A2(n_188), .B1(n_213), .B2(n_214), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_171), .A2(n_188), .B1(n_234), .B2(n_236), .Y(n_233) );
BUFx3_ASAP7_75t_L g189 ( .A(n_172), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g196 ( .A1(n_172), .A2(n_197), .B(n_204), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_172), .A2(n_222), .B(n_226), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_172), .A2(n_239), .B(n_244), .Y(n_238) );
NAND2x1p5_ASAP7_75t_L g473 ( .A(n_172), .B(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_L g486 ( .A(n_172), .B(n_474), .Y(n_486) );
INVx4_ASAP7_75t_SL g497 ( .A(n_172), .Y(n_497) );
AND2x2_ASAP7_75t_L g260 ( .A(n_175), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g274 ( .A(n_175), .B(n_195), .Y(n_274) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_176), .B(n_195), .Y(n_289) );
AND2x2_ASAP7_75t_L g301 ( .A(n_176), .B(n_277), .Y(n_301) );
OR2x2_ASAP7_75t_L g303 ( .A(n_176), .B(n_261), .Y(n_303) );
AND2x2_ASAP7_75t_L g338 ( .A(n_176), .B(n_261), .Y(n_338) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_176), .Y(n_383) );
INVx1_ASAP7_75t_L g391 ( .A(n_176), .Y(n_391) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_179), .B(n_190), .Y(n_176) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_177), .A2(n_196), .B(n_207), .Y(n_195) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_178), .B(n_482), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_183), .B(n_189), .Y(n_179) );
O2A1O1Ixp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .C(n_187), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_185), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_187), .A2(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx4_ASAP7_75t_L g574 ( .A(n_188), .Y(n_574) );
NAND3xp33_ASAP7_75t_L g211 ( .A(n_189), .B(n_212), .C(n_215), .Y(n_211) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_191), .A2(n_221), .B(n_229), .Y(n_220) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_191), .A2(n_238), .B(n_247), .Y(n_237) );
INVx2_ASAP7_75t_L g258 ( .A(n_191), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_191), .A2(n_485), .B(n_487), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_191), .A2(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g543 ( .A(n_191), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g308 ( .A1(n_192), .A2(n_309), .B1(n_313), .B2(n_317), .C(n_318), .Y(n_308) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g268 ( .A(n_193), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_208), .Y(n_193) );
INVx2_ASAP7_75t_L g267 ( .A(n_194), .Y(n_267) );
AND2x2_ASAP7_75t_L g320 ( .A(n_194), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g339 ( .A(n_194), .B(n_277), .Y(n_339) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g402 ( .A(n_195), .B(n_277), .Y(n_402) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .C(n_201), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_199), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_199), .A2(n_506), .B(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_201), .A2(n_550), .B(n_551), .C(n_552), .Y(n_549) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_202), .A2(n_227), .B(n_228), .Y(n_226) );
INVx4_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g493 ( .A(n_203), .Y(n_493) );
AND2x2_ASAP7_75t_L g324 ( .A(n_208), .B(n_269), .Y(n_324) );
OAI322xp33_ASAP7_75t_L g392 ( .A1(n_208), .A2(n_348), .A3(n_393), .B1(n_395), .B2(n_398), .C1(n_400), .C2(n_404), .Y(n_392) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2x1_ASAP7_75t_L g275 ( .A(n_209), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g288 ( .A(n_209), .Y(n_288) );
AND2x2_ASAP7_75t_L g397 ( .A(n_209), .B(n_277), .Y(n_397) );
AND2x2_ASAP7_75t_L g429 ( .A(n_209), .B(n_301), .Y(n_429) );
OR2x2_ASAP7_75t_L g432 ( .A(n_209), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
INVx1_ASAP7_75t_L g262 ( .A(n_210), .Y(n_262) );
AO21x1_ASAP7_75t_L g261 ( .A1(n_212), .A2(n_215), .B(n_262), .Y(n_261) );
AO21x2_ASAP7_75t_L g470 ( .A1(n_215), .A2(n_471), .B(n_481), .Y(n_470) );
INVx3_ASAP7_75t_L g517 ( .A(n_215), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_215), .B(n_529), .Y(n_528) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_215), .A2(n_547), .B(n_554), .Y(n_546) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_230), .Y(n_217) );
INVx1_ASAP7_75t_L g445 ( .A(n_218), .Y(n_445) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g250 ( .A(n_219), .B(n_237), .Y(n_250) );
INVx2_ASAP7_75t_L g285 ( .A(n_219), .Y(n_285) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g307 ( .A(n_220), .Y(n_307) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_220), .Y(n_315) );
OR2x2_ASAP7_75t_L g439 ( .A(n_220), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g264 ( .A(n_230), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g304 ( .A(n_230), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g356 ( .A(n_230), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
AND2x2_ASAP7_75t_L g251 ( .A(n_231), .B(n_252), .Y(n_251) );
NOR2xp67_ASAP7_75t_L g311 ( .A(n_231), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g365 ( .A(n_231), .B(n_253), .Y(n_365) );
OR2x2_ASAP7_75t_L g373 ( .A(n_231), .B(n_307), .Y(n_373) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
BUFx2_ASAP7_75t_L g282 ( .A(n_232), .Y(n_282) );
AND2x2_ASAP7_75t_L g292 ( .A(n_232), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g316 ( .A(n_232), .B(n_237), .Y(n_316) );
AND2x2_ASAP7_75t_L g380 ( .A(n_232), .B(n_253), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_237), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_237), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g293 ( .A(n_237), .Y(n_293) );
INVx1_ASAP7_75t_L g298 ( .A(n_237), .Y(n_298) );
AND2x2_ASAP7_75t_L g310 ( .A(n_237), .B(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_237), .Y(n_388) );
INVx1_ASAP7_75t_L g440 ( .A(n_237), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_242), .Y(n_239) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
AND2x2_ASAP7_75t_L g417 ( .A(n_249), .B(n_326), .Y(n_417) );
INVx2_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g344 ( .A(n_251), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g443 ( .A(n_251), .B(n_378), .Y(n_443) );
INVx1_ASAP7_75t_L g265 ( .A(n_252), .Y(n_265) );
AND2x2_ASAP7_75t_L g291 ( .A(n_252), .B(n_285), .Y(n_291) );
BUFx2_ASAP7_75t_L g350 ( .A(n_252), .Y(n_350) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_253), .Y(n_271) );
INVx1_ASAP7_75t_L g281 ( .A(n_253), .Y(n_281) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_256), .Y(n_495) );
INVx2_ASAP7_75t_L g575 ( .A(n_256), .Y(n_575) );
INVx1_ASAP7_75t_L g540 ( .A(n_258), .Y(n_540) );
NOR2xp67_ASAP7_75t_L g419 ( .A(n_259), .B(n_266), .Y(n_419) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AOI32xp33_ASAP7_75t_L g263 ( .A1(n_260), .A2(n_264), .A3(n_266), .B1(n_268), .B2(n_270), .Y(n_263) );
AND2x2_ASAP7_75t_L g403 ( .A(n_260), .B(n_276), .Y(n_403) );
AND2x2_ASAP7_75t_L g441 ( .A(n_260), .B(n_339), .Y(n_441) );
INVx1_ASAP7_75t_L g321 ( .A(n_261), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_265), .B(n_327), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_266), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_266), .B(n_269), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_266), .B(n_338), .Y(n_420) );
OR2x2_ASAP7_75t_L g434 ( .A(n_266), .B(n_303), .Y(n_434) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g361 ( .A(n_267), .B(n_269), .Y(n_361) );
OR2x2_ASAP7_75t_L g370 ( .A(n_267), .B(n_357), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_269), .B(n_320), .Y(n_342) );
INVx2_ASAP7_75t_L g357 ( .A(n_271), .Y(n_357) );
OR2x2_ASAP7_75t_L g372 ( .A(n_271), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g387 ( .A(n_271), .B(n_388), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g444 ( .A1(n_271), .A2(n_364), .B(n_445), .C(n_446), .Y(n_444) );
OAI321xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_278), .A3(n_283), .B1(n_286), .B2(n_290), .C(n_294), .Y(n_272) );
INVx1_ASAP7_75t_L g385 ( .A(n_273), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x2_ASAP7_75t_L g396 ( .A(n_274), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g348 ( .A(n_276), .Y(n_348) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_277), .B(n_391), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_278), .A2(n_416), .B1(n_418), .B2(n_420), .C(n_421), .Y(n_415) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
AND2x2_ASAP7_75t_L g353 ( .A(n_280), .B(n_327), .Y(n_353) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_281), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g326 ( .A(n_282), .Y(n_326) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_283), .A2(n_324), .B(n_369), .C(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g335 ( .A(n_285), .B(n_292), .Y(n_335) );
BUFx2_ASAP7_75t_L g345 ( .A(n_285), .Y(n_345) );
INVx1_ASAP7_75t_L g360 ( .A(n_285), .Y(n_360) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
OR2x2_ASAP7_75t_L g366 ( .A(n_288), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g449 ( .A(n_288), .Y(n_449) );
INVx1_ASAP7_75t_L g442 ( .A(n_289), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x2_ASAP7_75t_L g295 ( .A(n_291), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g399 ( .A(n_291), .B(n_316), .Y(n_399) );
INVx1_ASAP7_75t_L g328 ( .A(n_292), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_299), .B1(n_302), .B2(n_304), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_296), .B(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g364 ( .A(n_297), .B(n_365), .Y(n_364) );
BUFx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_SL g327 ( .A(n_298), .B(n_307), .Y(n_327) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g319 ( .A(n_301), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g329 ( .A(n_303), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_306), .A2(n_424), .B1(n_426), .B2(n_427), .C(n_428), .Y(n_423) );
INVx1_ASAP7_75t_L g312 ( .A(n_307), .Y(n_312) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_307), .Y(n_378) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_310), .B(n_429), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g318 ( .A1(n_311), .A2(n_316), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_314), .B(n_324), .Y(n_421) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g390 ( .A(n_315), .Y(n_390) );
AND2x2_ASAP7_75t_L g349 ( .A(n_316), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g438 ( .A(n_316), .Y(n_438) );
INVx1_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
INVx1_ASAP7_75t_L g409 ( .A(n_320), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_325), .B1(n_328), .B2(n_329), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_326), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g394 ( .A(n_327), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_327), .B(n_365), .Y(n_431) );
OR2x2_ASAP7_75t_L g404 ( .A(n_328), .B(n_357), .Y(n_404) );
INVx1_ASAP7_75t_L g343 ( .A(n_329), .Y(n_343) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_331), .B(n_382), .Y(n_381) );
NOR3xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_351), .C(n_362), .Y(n_332) );
OAI211xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B(n_340), .C(n_346), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_335), .A2(n_406), .B1(n_410), .B2(n_413), .C(n_415), .Y(n_405) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
AND2x2_ASAP7_75t_L g347 ( .A(n_338), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g401 ( .A(n_338), .B(n_402), .Y(n_401) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_339), .A2(n_387), .B(n_389), .C(n_391), .Y(n_386) );
INVx2_ASAP7_75t_L g433 ( .A(n_339), .Y(n_433) );
OAI21xp5_ASAP7_75t_SL g340 ( .A1(n_341), .A2(n_343), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g412 ( .A(n_345), .B(n_365), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
OAI21xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_354), .B(n_355), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI21xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_358), .B(n_361), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_356), .B(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_361), .B(n_448), .Y(n_447) );
OAI21xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B(n_368), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g389 ( .A(n_365), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND4x1_ASAP7_75t_L g374 ( .A(n_375), .B(n_405), .C(n_422), .D(n_444), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_392), .Y(n_375) );
OAI211xp5_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_381), .B(n_384), .C(n_386), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_380), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_391), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g426 ( .A(n_401), .Y(n_426) );
INVx2_ASAP7_75t_SL g414 ( .A(n_402), .Y(n_414) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g427 ( .A(n_412), .Y(n_427) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NOR2xp33_ASAP7_75t_SL g422 ( .A(n_423), .B(n_430), .Y(n_422) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
OAI221xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_432), .B1(n_434), .B2(n_435), .C(n_436), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_441), .B1(n_442), .B2(n_443), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_451), .B(n_456), .C(n_767), .Y(n_455) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_459), .B1(n_462), .B2(n_746), .Y(n_457) );
INVx1_ASAP7_75t_L g761 ( .A(n_458), .Y(n_761) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g762 ( .A(n_460), .Y(n_762) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI22xp5_ASAP7_75t_SL g760 ( .A1(n_463), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_760) );
OR3x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_644), .C(n_709), .Y(n_463) );
NAND4xp25_ASAP7_75t_SL g464 ( .A(n_465), .B(n_585), .C(n_611), .D(n_634), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_518), .B1(n_555), .B2(n_562), .C(n_577), .Y(n_465) );
CKINVDCx14_ASAP7_75t_R g466 ( .A(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_467), .A2(n_578), .B1(n_602), .B2(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_499), .Y(n_467) );
INVx1_ASAP7_75t_SL g638 ( .A(n_468), .Y(n_638) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_483), .Y(n_468) );
OR2x2_ASAP7_75t_L g560 ( .A(n_469), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g580 ( .A(n_469), .B(n_500), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_469), .B(n_508), .Y(n_593) );
AND2x2_ASAP7_75t_L g610 ( .A(n_469), .B(n_483), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_469), .B(n_558), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_469), .B(n_609), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_469), .B(n_499), .Y(n_731) );
AOI211xp5_ASAP7_75t_SL g742 ( .A1(n_469), .A2(n_648), .B(n_743), .C(n_744), .Y(n_742) );
INVx5_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_470), .B(n_500), .Y(n_614) );
AND2x2_ASAP7_75t_L g617 ( .A(n_470), .B(n_501), .Y(n_617) );
OR2x2_ASAP7_75t_L g662 ( .A(n_470), .B(n_500), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_470), .B(n_508), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_475), .Y(n_471) );
INVx5_ASAP7_75t_L g489 ( .A(n_476), .Y(n_489) );
INVx5_ASAP7_75t_SL g561 ( .A(n_483), .Y(n_561) );
AND2x2_ASAP7_75t_L g579 ( .A(n_483), .B(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_483), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g665 ( .A(n_483), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g697 ( .A(n_483), .B(n_508), .Y(n_697) );
OR2x2_ASAP7_75t_L g703 ( .A(n_483), .B(n_593), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_483), .B(n_653), .Y(n_712) );
OR2x6_ASAP7_75t_L g483 ( .A(n_484), .B(n_498), .Y(n_483) );
BUFx2_ASAP7_75t_L g535 ( .A(n_486), .Y(n_535) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_489), .A2(n_497), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_SL g569 ( .A1(n_489), .A2(n_497), .B(n_570), .C(n_571), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B(n_494), .C(n_495), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_492), .A2(n_495), .B(n_526), .C(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_508), .Y(n_499) );
AND2x2_ASAP7_75t_L g594 ( .A(n_500), .B(n_561), .Y(n_594) );
INVx1_ASAP7_75t_SL g607 ( .A(n_500), .Y(n_607) );
OR2x2_ASAP7_75t_L g642 ( .A(n_500), .B(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g648 ( .A(n_500), .B(n_508), .Y(n_648) );
AND2x2_ASAP7_75t_L g706 ( .A(n_500), .B(n_558), .Y(n_706) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_501), .B(n_561), .Y(n_633) );
INVx3_ASAP7_75t_L g558 ( .A(n_508), .Y(n_558) );
OR2x2_ASAP7_75t_L g599 ( .A(n_508), .B(n_561), .Y(n_599) );
AND2x2_ASAP7_75t_L g609 ( .A(n_508), .B(n_607), .Y(n_609) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_508), .Y(n_657) );
AND2x2_ASAP7_75t_L g666 ( .A(n_508), .B(n_580), .Y(n_666) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_516), .Y(n_508) );
OA21x2_ASAP7_75t_L g567 ( .A1(n_517), .A2(n_568), .B(n_576), .Y(n_567) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_518), .A2(n_683), .B1(n_685), .B2(n_687), .C(n_690), .Y(n_682) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_530), .Y(n_519) );
AND2x2_ASAP7_75t_L g656 ( .A(n_520), .B(n_637), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_520), .B(n_715), .Y(n_719) );
OR2x2_ASAP7_75t_L g740 ( .A(n_520), .B(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_520), .B(n_745), .Y(n_744) );
BUFx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx5_ASAP7_75t_L g587 ( .A(n_521), .Y(n_587) );
AND2x2_ASAP7_75t_L g664 ( .A(n_521), .B(n_532), .Y(n_664) );
AND2x2_ASAP7_75t_L g725 ( .A(n_521), .B(n_604), .Y(n_725) );
AND2x2_ASAP7_75t_L g738 ( .A(n_521), .B(n_558), .Y(n_738) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_544), .Y(n_530) );
AND2x4_ASAP7_75t_L g565 ( .A(n_531), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g583 ( .A(n_531), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
AND2x2_ASAP7_75t_L g659 ( .A(n_531), .B(n_637), .Y(n_659) );
AND2x2_ASAP7_75t_L g669 ( .A(n_531), .B(n_587), .Y(n_669) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_531), .Y(n_677) );
AND2x2_ASAP7_75t_L g689 ( .A(n_531), .B(n_567), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_531), .B(n_621), .Y(n_693) );
AND2x2_ASAP7_75t_L g730 ( .A(n_531), .B(n_725), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_531), .B(n_604), .Y(n_741) );
OR2x2_ASAP7_75t_L g743 ( .A(n_531), .B(n_679), .Y(n_743) );
INVx5_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g629 ( .A(n_532), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g639 ( .A(n_532), .B(n_584), .Y(n_639) );
AND2x2_ASAP7_75t_L g651 ( .A(n_532), .B(n_567), .Y(n_651) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_532), .Y(n_681) );
AND2x4_ASAP7_75t_L g715 ( .A(n_532), .B(n_566), .Y(n_715) );
OR2x6_ASAP7_75t_L g532 ( .A(n_533), .B(n_541), .Y(n_532) );
AOI21xp5_ASAP7_75t_SL g533 ( .A1(n_534), .A2(n_536), .B(n_540), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
BUFx2_ASAP7_75t_L g564 ( .A(n_544), .Y(n_564) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g604 ( .A(n_545), .Y(n_604) );
AND2x2_ASAP7_75t_L g637 ( .A(n_545), .B(n_567), .Y(n_637) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g584 ( .A(n_546), .B(n_567), .Y(n_584) );
BUFx2_ASAP7_75t_L g630 ( .A(n_546), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_553), .Y(n_547) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_557), .B(n_638), .Y(n_717) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_558), .B(n_580), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_558), .B(n_561), .Y(n_619) );
AND2x2_ASAP7_75t_L g674 ( .A(n_558), .B(n_610), .Y(n_674) );
AOI221xp5_ASAP7_75t_SL g611 ( .A1(n_559), .A2(n_612), .B1(n_620), .B2(n_622), .C(n_626), .Y(n_611) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g606 ( .A(n_560), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g647 ( .A(n_560), .B(n_648), .Y(n_647) );
OAI321xp33_ASAP7_75t_L g654 ( .A1(n_560), .A2(n_613), .A3(n_655), .B1(n_657), .B2(n_658), .C(n_660), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_561), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_564), .B(n_715), .Y(n_733) );
AND2x2_ASAP7_75t_L g620 ( .A(n_565), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_565), .B(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_566), .Y(n_596) );
AND2x2_ASAP7_75t_L g603 ( .A(n_566), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_566), .B(n_678), .Y(n_708) );
INVx1_ASAP7_75t_L g745 ( .A(n_566), .Y(n_745) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B(n_582), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_579), .A2(n_689), .B(n_738), .C(n_739), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_580), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_580), .B(n_618), .Y(n_684) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g627 ( .A(n_584), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_584), .B(n_587), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_584), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_584), .B(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B1(n_600), .B2(n_605), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g601 ( .A(n_587), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g624 ( .A(n_587), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g636 ( .A(n_587), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_587), .B(n_630), .Y(n_672) );
OR2x2_ASAP7_75t_L g679 ( .A(n_587), .B(n_604), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_587), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g729 ( .A(n_587), .B(n_715), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B1(n_595), .B2(n_597), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g635 ( .A(n_590), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_593), .A2(n_608), .B1(n_676), .B2(n_680), .Y(n_675) );
INVx1_ASAP7_75t_L g723 ( .A(n_594), .Y(n_723) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_598), .A2(n_635), .B1(n_638), .B2(n_639), .C(n_640), .Y(n_634) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g613 ( .A(n_599), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_603), .B(n_669), .Y(n_701) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_604), .Y(n_621) );
INVx1_ASAP7_75t_L g625 ( .A(n_604), .Y(n_625) );
NAND2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g643 ( .A(n_610), .Y(n_643) );
AND2x2_ASAP7_75t_L g652 ( .A(n_610), .B(n_653), .Y(n_652) );
NAND2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx2_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g696 ( .A(n_617), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_620), .A2(n_646), .B1(n_649), .B2(n_652), .C(n_654), .Y(n_645) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_624), .B(n_681), .Y(n_680) );
AOI21xp33_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_628), .B(n_631), .Y(n_626) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
CKINVDCx16_ASAP7_75t_R g728 ( .A(n_631), .Y(n_728) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
OR2x2_ASAP7_75t_L g670 ( .A(n_633), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g691 ( .A(n_636), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_636), .B(n_696), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_639), .B(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g644 ( .A(n_645), .B(n_663), .C(n_682), .D(n_695), .Y(n_644) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g653 ( .A(n_648), .Y(n_653) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g686 ( .A(n_657), .B(n_662), .Y(n_686) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B(n_667), .C(n_675), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g734 ( .A1(n_665), .A2(n_707), .B(n_735), .C(n_742), .Y(n_734) );
INVx1_ASAP7_75t_SL g694 ( .A(n_666), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B1(n_672), .B2(n_673), .Y(n_667) );
INVx1_ASAP7_75t_L g698 ( .A(n_672), .Y(n_698) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_678), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_678), .B(n_689), .Y(n_722) );
INVx2_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g699 ( .A(n_689), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B(n_694), .Y(n_690) );
INVxp33_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI322xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .A3(n_699), .B1(n_700), .B2(n_702), .C1(n_704), .C2(n_707), .Y(n_695) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND3xp33_ASAP7_75t_SL g709 ( .A(n_710), .B(n_727), .C(n_734), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_713), .B1(n_716), .B2(n_718), .C(n_720), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g726 ( .A(n_715), .Y(n_726) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_730), .B2(n_731), .C(n_732), .Y(n_727) );
NAND2xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g763 ( .A(n_747), .Y(n_763) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
CKINVDCx16_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
CKINVDCx16_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g758 ( .A(n_755), .Y(n_758) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx3_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
endmodule