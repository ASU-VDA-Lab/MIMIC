module real_jpeg_15321_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_0),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_0),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_0),
.B(n_581),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_20),
.B(n_587),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_1),
.B(n_588),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_2),
.B(n_68),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_2),
.B(n_142),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_2),
.B(n_181),
.Y(n_180)
);

NAND2x1_ASAP7_75t_L g205 ( 
.A(n_2),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_2),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_2),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_2),
.B(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_3),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_3),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_3),
.Y(n_299)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_4),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_4),
.Y(n_218)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_5),
.Y(n_116)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_5),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_5),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_5),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_5),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_5),
.Y(n_467)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_6),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_7),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_7),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_7),
.B(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_7),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_7),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_7),
.B(n_308),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_7),
.B(n_142),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_7),
.B(n_144),
.Y(n_448)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_8),
.Y(n_142)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

BUFx4f_ASAP7_75t_L g256 ( 
.A(n_8),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_8),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_9),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_9),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_9),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_9),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_9),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_9),
.B(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_9),
.B(n_493),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_10),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_10),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_10),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_10),
.B(n_55),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_10),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_10),
.B(n_152),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_10),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_10),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_11),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_11),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_11),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_11),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_11),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_11),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_11),
.B(n_206),
.Y(n_348)
);

AOI22x1_ASAP7_75t_L g149 ( 
.A1(n_12),
.A2(n_15),
.B1(n_150),
.B2(n_154),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_12),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_12),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_12),
.B(n_302),
.Y(n_301)
);

AOI31xp67_ASAP7_75t_L g377 ( 
.A1(n_12),
.A2(n_149),
.A3(n_378),
.B(n_381),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_12),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_12),
.B(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_12),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_12),
.B(n_480),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_13),
.Y(n_270)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_13),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_14),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_14),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_14),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_14),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_14),
.B(n_246),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_14),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_14),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_14),
.B(n_153),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_15),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_15),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_15),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_15),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_15),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_15),
.B(n_272),
.Y(n_271)
);

NAND2x1_ASAP7_75t_L g343 ( 
.A(n_15),
.B(n_344),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_15),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_16),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_16),
.Y(n_274)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_16),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_16),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g106 ( 
.A(n_18),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_575),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_124),
.B(n_574),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_77),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_24),
.B(n_77),
.Y(n_574)
);

BUFx24_ASAP7_75t_SL g589 ( 
.A(n_24),
.Y(n_589)
);

FAx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_43),
.CI(n_57),
.CON(n_24),
.SN(n_24)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_25),
.B(n_43),
.C(n_57),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.C(n_37),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_26),
.A2(n_32),
.B1(n_50),
.B2(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_SL g578 ( 
.A(n_26),
.B(n_45),
.C(n_52),
.Y(n_578)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_30),
.Y(n_87)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_31),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_67),
.C(n_72),
.Y(n_66)
);

AOI22x1_ASAP7_75t_L g119 ( 
.A1(n_32),
.A2(n_61),
.B1(n_72),
.B2(n_73),
.Y(n_119)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_36),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_52),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_45),
.A2(n_51),
.B1(n_580),
.B2(n_584),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_49),
.B(n_113),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_49),
.B(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_56),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.C(n_66),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_58),
.A2(n_59),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_62),
.B(n_66),
.Y(n_123)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XOR2x1_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_70),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_72),
.A2(n_73),
.B1(n_112),
.B2(n_335),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_108),
.C(n_112),
.Y(n_107)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_76),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_120),
.C(n_121),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_78),
.B(n_549),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_107),
.C(n_117),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_79),
.B(n_547),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_88),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_85),
.C(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_84),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_84),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_97),
.C(n_104),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_89),
.A2(n_90),
.B1(n_97),
.B2(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_96),
.Y(n_188)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_96),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_96),
.Y(n_333)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_98),
.Y(n_538)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_102),
.Y(n_225)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_102),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_104),
.B(n_537),
.Y(n_536)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_107),
.B(n_118),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_SL g541 ( 
.A(n_108),
.B(n_542),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_112),
.A2(n_254),
.B1(n_257),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_112),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_112),
.B(n_257),
.C(n_330),
.Y(n_543)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_116),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_120),
.B(n_121),
.Y(n_549)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21x1_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_529),
.B(n_569),
.Y(n_124)
);

AO21x2_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_362),
.B(n_526),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_323),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_277),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_128),
.B(n_277),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_201),
.Y(n_128)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_129),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_166),
.C(n_189),
.Y(n_129)
);

INVxp33_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_131),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_148),
.C(n_158),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_132),
.B(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g539 ( 
.A(n_133),
.B(n_245),
.C(n_355),
.Y(n_539)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_134),
.B(n_245),
.Y(n_352)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_139),
.C(n_143),
.Y(n_192)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_137),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_142),
.Y(n_295)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_148),
.A2(n_149),
.B1(n_158),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_158),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.C(n_165),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_159),
.A2(n_160),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_159),
.A2(n_160),
.B1(n_165),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_160),
.B(n_232),
.C(n_254),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_163),
.B(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_165),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_167),
.A2(n_190),
.B1(n_191),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_167),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_179),
.C(n_184),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_168),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.C(n_175),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_169),
.A2(n_175),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_169),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_169),
.B(n_429),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_171),
.Y(n_476)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_173),
.B(n_374),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_175),
.Y(n_376)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_177),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_179),
.A2(n_180),
.B1(n_184),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_184),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_194),
.C(n_198),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_194),
.A2(n_195),
.B1(n_390),
.B2(n_391),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_195),
.Y(n_389)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx8_ASAP7_75t_L g488 ( 
.A(n_200),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_250),
.B1(n_275),
.B2(n_276),
.Y(n_201)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_240),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_SL g325 ( 
.A(n_203),
.B(n_241),
.C(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_214),
.C(n_226),
.Y(n_203)
);

XNOR2x2_ASAP7_75t_SL g283 ( 
.A(n_204),
.B(n_284),
.Y(n_283)
);

XOR2x1_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_208),
.C(n_211),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_214),
.B(n_226),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.C(n_223),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_215),
.A2(n_223),
.B1(n_224),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_215),
.Y(n_322)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_218),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_219),
.B(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_223),
.B(n_409),
.C(n_411),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_223),
.A2(n_224),
.B1(n_409),
.B2(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_232),
.C(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_234),
.B1(n_235),
.B2(n_239),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_232),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_232),
.A2(n_239),
.B1(n_254),
.B2(n_257),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_233),
.Y(n_384)
);

INVx6_ASAP7_75t_L g481 ( 
.A(n_233),
.Y(n_481)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_242),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_243),
.B(n_249),
.C(n_357),
.Y(n_356)
);

XNOR2x1_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_245),
.Y(n_357)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_250),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_258),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_251),
.B(n_259),
.C(n_261),
.Y(n_358)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_254),
.Y(n_257)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_255),
.Y(n_447)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_256),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_262),
.B(n_267),
.C(n_271),
.Y(n_337)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_270),
.Y(n_347)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_275),
.B(n_360),
.C(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_283),
.C(n_285),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_283),
.Y(n_367)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_286),
.B(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_316),
.C(n_320),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_287),
.B(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.C(n_300),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2x1_ASAP7_75t_SL g416 ( 
.A(n_289),
.B(n_417),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_L g417 ( 
.A(n_292),
.B(n_300),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_297),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_293),
.B(n_297),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_307),
.C(n_311),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_301),
.A2(n_307),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_301),
.Y(n_405)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_307),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_307),
.A2(n_406),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_307),
.B(n_474),
.C(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2x1_ASAP7_75t_SL g403 ( 
.A(n_311),
.B(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_317),
.B(n_320),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_323),
.A2(n_527),
.B(n_528),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_359),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_324),
.B(n_359),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_325),
.B(n_328),
.C(n_349),
.Y(n_565)
);

XNOR2x1_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_349),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_336),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_329),
.B(n_337),
.C(n_338),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_334),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_332),
.Y(n_410)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_339),
.B(n_343),
.C(n_348),
.Y(n_544)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_348),
.Y(n_342)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2x1_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_358),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_356),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_351),
.B(n_356),
.C(n_563),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_353),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_358),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_420),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_368),
.C(n_397),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_365),
.B(n_369),
.Y(n_422)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.C(n_393),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_372),
.B(n_394),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_377),
.C(n_385),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_377),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_375),
.B(n_430),
.C(n_434),
.Y(n_453)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx6_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_400),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_389),
.C(n_390),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_386),
.B(n_515),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

XNOR2x1_ASAP7_75t_SL g460 ( 
.A(n_387),
.B(n_388),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_387),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_387),
.A2(n_478),
.B1(n_479),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NOR2x1_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_418),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_418),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_401),
.C(n_416),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_399),
.B(n_524),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_402),
.B(n_416),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_407),
.C(n_414),
.Y(n_402)
);

XOR2x1_ASAP7_75t_L g509 ( 
.A(n_403),
.B(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_408),
.B(n_415),
.Y(n_510)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_409),
.Y(n_456)
);

XOR2x2_ASAP7_75t_L g454 ( 
.A(n_411),
.B(n_455),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NAND3xp33_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.C(n_423),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_424),
.A2(n_521),
.B(n_525),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_506),
.B(n_520),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_468),
.B(n_505),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_451),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_427),
.B(n_451),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_436),
.C(n_445),
.Y(n_427)
);

XOR2x1_ASAP7_75t_SL g499 ( 
.A(n_428),
.B(n_500),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_434),
.Y(n_429)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_436),
.A2(n_437),
.B1(n_445),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_444),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_444),
.Y(n_472)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_445),
.Y(n_501)
);

AO22x1_ASAP7_75t_SL g445 ( 
.A1(n_446),
.A2(n_448),
.B1(n_449),
.B2(n_450),
.Y(n_445)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_446),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_448),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_448),
.B(n_449),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_450),
.B(n_492),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_457),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_453),
.B(n_454),
.C(n_519),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_457),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

MAJx2_ASAP7_75t_L g517 ( 
.A(n_458),
.B(n_460),
.C(n_461),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx6_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_498),
.B(n_504),
.Y(n_468)
);

OAI21x1_ASAP7_75t_SL g469 ( 
.A1(n_470),
.A2(n_482),
.B(n_497),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_477),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_477),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_472),
.Y(n_503)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_479),
.Y(n_490)
);

INVx6_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_483),
.A2(n_491),
.B(n_496),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_489),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_489),
.Y(n_496)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_502),
.Y(n_498)
);

NOR2xp67_ASAP7_75t_L g504 ( 
.A(n_499),
.B(n_502),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_507),
.B(n_518),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_518),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_509),
.B1(n_511),
.B2(n_512),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_513),
.C(n_517),
.Y(n_522)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_514),
.B1(n_516),
.B2(n_517),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_523),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_522),
.B(n_523),
.Y(n_525)
);

NOR3xp33_ASAP7_75t_SL g529 ( 
.A(n_530),
.B(n_550),
.C(n_564),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_530),
.A2(n_570),
.B(n_573),
.Y(n_569)
);

NOR2xp67_ASAP7_75t_R g530 ( 
.A(n_531),
.B(n_548),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_531),
.B(n_548),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_540),
.C(n_545),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_532),
.B(n_553),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_535),
.C(n_539),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_559),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_536),
.B(n_539),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_540),
.A2(n_545),
.B1(n_546),
.B2(n_554),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g554 ( 
.A(n_540),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_543),
.C(n_544),
.Y(n_540)
);

XNOR2x2_ASAP7_75t_SL g560 ( 
.A(n_541),
.B(n_561),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_543),
.B(n_544),
.Y(n_561)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_551),
.A2(n_571),
.B(n_572),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_552),
.B(n_555),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_552),
.B(n_555),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_560),
.C(n_562),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_557),
.A2(n_558),
.B1(n_560),
.B2(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_560),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_562),
.B(n_567),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_566),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_SL g571 ( 
.A(n_565),
.B(n_566),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_576),
.B(n_586),
.Y(n_575)
);

NOR2xp67_ASAP7_75t_R g576 ( 
.A(n_577),
.B(n_585),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_577),
.B(n_585),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_578),
.B(n_579),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_580),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_582),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);


endmodule