module fake_jpeg_7257_n_98 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_98);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_12),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_22),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_17),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_24),
.B1(n_13),
.B2(n_15),
.Y(n_41)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_16),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_22),
.B1(n_17),
.B2(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_33),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_33),
.B(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_13),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_19),
.B1(n_21),
.B2(n_20),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_28),
.B(n_27),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_54),
.B1(n_55),
.B2(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_28),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_32),
.B1(n_26),
.B2(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_21),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_60),
.B(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

OAI22x1_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_38),
.B1(n_27),
.B2(n_29),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_48),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_71),
.B1(n_74),
.B2(n_58),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_46),
.C(n_42),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_63),
.Y(n_80)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_53),
.C(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_15),
.Y(n_75)
);

BUFx24_ASAP7_75t_SL g76 ( 
.A(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_5),
.B(n_7),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_86),
.B(n_76),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_11),
.C(n_8),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_90),
.C(n_9),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_81),
.B(n_78),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_78),
.B(n_8),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_7),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_93),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_97),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_92),
.Y(n_97)
);


endmodule