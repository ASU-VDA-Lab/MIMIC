module fake_jpeg_14489_n_169 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_14),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_4),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_19),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_36),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_15),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_79),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx6p67_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_1),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_81),
.B1(n_70),
.B2(n_54),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_63),
.B1(n_51),
.B2(n_66),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_72),
.C(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_90),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_47),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_54),
.B1(n_70),
.B2(n_58),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_47),
.B1(n_62),
.B2(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

BUFx2_ASAP7_75t_SL g98 ( 
.A(n_91),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_105),
.Y(n_120)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_65),
.A3(n_55),
.B1(n_57),
.B2(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_69),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_107),
.Y(n_132)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_114),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_50),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_113),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_52),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_53),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_97),
.B(n_112),
.C(n_100),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_56),
.B1(n_49),
.B2(n_48),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_122),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_50),
.B(n_68),
.C(n_26),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_1),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_130),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_25),
.B(n_45),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_29),
.B(n_39),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_131),
.B(n_4),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_134),
.A2(n_2),
.B(n_3),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_145),
.B(n_120),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_142),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_146),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_119),
.B(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_124),
.B1(n_116),
.B2(n_128),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_144),
.B1(n_117),
.B2(n_119),
.Y(n_151)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_151),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_145),
.C(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_10),
.Y(n_152)
);

OAI322xp33_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_141),
.A3(n_12),
.B1(n_13),
.B2(n_11),
.C1(n_18),
.C2(n_27),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_121),
.C(n_31),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_139),
.C(n_17),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_157),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_156),
.B(n_148),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_139),
.C(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_160),
.C(n_158),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_158),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_37),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_44),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_153),
.Y(n_169)
);


endmodule