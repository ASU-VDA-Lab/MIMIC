module fake_netlist_5_2224_n_174 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_174);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_174;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_124;
wire n_136;
wire n_146;
wire n_86;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_123;
wire n_38;
wire n_139;
wire n_113;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_53;
wire n_160;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_77;
wire n_102;
wire n_106;
wire n_64;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_5),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_6),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_6),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NAND2x1p5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_50),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

OR2x6_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_14),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_44),
.B(n_53),
.C(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_37),
.B(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_48),
.Y(n_82)
);

INVxp67_ASAP7_75t_SL g83 ( 
.A(n_66),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_26),
.B(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_75),
.Y(n_88)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_69),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_74),
.B(n_71),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_69),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_73),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_71),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_62),
.B1(n_59),
.B2(n_69),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_62),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_85),
.B(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

AO21x2_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_78),
.B(n_61),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_97),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_103),
.C(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_104),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_94),
.B1(n_100),
.B2(n_59),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_101),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_122),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_107),
.B(n_111),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_109),
.B(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_101),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_124),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_89),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_89),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_56),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_108),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_61),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_134),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_64),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_132),
.Y(n_144)
);

OAI22x1_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_64),
.B1(n_126),
.B2(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

AND3x4_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_93),
.C(n_135),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_140),
.C(n_128),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_129),
.C(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_111),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_111),
.B1(n_95),
.B2(n_107),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_150),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_77),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

AND2x4_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_152),
.Y(n_162)
);

OR3x2_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_145),
.C(n_79),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_88),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_160),
.C(n_159),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_155),
.B1(n_160),
.B2(n_95),
.Y(n_167)
);

NOR4xp25_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_81),
.C(n_79),
.D(n_86),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

AOI31xp33_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_162),
.A3(n_161),
.B(n_165),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_162),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_86),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_SL g173 ( 
.A(n_169),
.B(n_105),
.C(n_113),
.Y(n_173)
);

OAI221xp5_ASAP7_75t_R g174 ( 
.A1(n_173),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.C(n_98),
.Y(n_174)
);


endmodule