module fake_netlist_5_778_n_18332 (n_924, n_977, n_2253, n_2417, n_2756, n_4706, n_2380, n_3241, n_3006, n_532, n_2327, n_1488, n_2899, n_790, n_3619, n_3541, n_3622, n_2395, n_2347, n_4963, n_4240, n_4508, n_2021, n_2391, n_5035, n_1960, n_2843, n_4, n_551, n_3615, n_2059, n_1466, n_1695, n_2487, n_3202, n_4977, n_3813, n_671, n_3341, n_3587, n_4128, n_3445, n_2001, n_4145, n_3785, n_5033, n_1462, n_4211, n_3448, n_3019, n_2096, n_877, n_3776, n_2530, n_4517, n_1696, n_2483, n_4425, n_4950, n_4988, n_1285, n_1860, n_4615, n_87, n_1107, n_1728, n_2076, n_668, n_301, n_2147, n_3010, n_2770, n_4131, n_2584, n_171, n_3188, n_3403, n_3624, n_3461, n_3082, n_2189, n_3796, n_1242, n_3283, n_519, n_2323, n_2597, n_3340, n_3277, n_281, n_2052, n_4499, n_4927, n_731, n_1314, n_1512, n_1490, n_317, n_569, n_3214, n_1517, n_2091, n_4311, n_3631, n_3806, n_4691, n_1449, n_4678, n_1566, n_2032, n_297, n_2587, n_156, n_219, n_157, n_3947, n_3490, n_600, n_223, n_1948, n_3868, n_3183, n_3437, n_3353, n_264, n_4203, n_3687, n_882, n_2384, n_3156, n_696, n_3376, n_646, n_5037, n_436, n_4468, n_3653, n_3702, n_1040, n_4976, n_2202, n_2648, n_5008, n_2159, n_2976, n_3876, n_2353, n_2439, n_4811, n_2276, n_2089, n_3420, n_72, n_1561, n_1165, n_1034, n_3361, n_4758, n_1600, n_521, n_845, n_528, n_4255, n_1796, n_395, n_553, n_901, n_4484, n_3668, n_4237, n_2934, n_1672, n_1880, n_3550, n_1626, n_637, n_144, n_2079, n_2238, n_96, n_1151, n_1405, n_1706, n_3418, n_342, n_4901, n_197, n_2859, n_1075, n_3395, n_4917, n_2863, n_2072, n_2738, n_2968, n_1585, n_2684, n_3593, n_1599, n_4421, n_4836, n_4020, n_2730, n_2251, n_3915, n_1377, n_4469, n_4414, n_190, n_4532, n_3339, n_228, n_283, n_3349, n_3735, n_2248, n_3007, n_1000, n_2622, n_2062, n_2668, n_1002, n_2100, n_310, n_3310, n_54, n_3487, n_2258, n_748, n_1058, n_1667, n_838, n_3983, n_332, n_1053, n_1224, n_4405, n_1926, n_1331, n_4195, n_279, n_1014, n_4969, n_1241, n_4504, n_1385, n_440, n_793, n_2776, n_4408, n_2140, n_2385, n_1819, n_4531, n_476, n_2987, n_1527, n_4567, n_4164, n_4234, n_345, n_4130, n_3611, n_2862, n_2175, n_2324, n_2606, n_3187, n_2828, n_182, n_4471, n_5031, n_407, n_3392, n_3975, n_3430, n_4444, n_3208, n_207, n_3331, n_2379, n_4983, n_2911, n_2154, n_4916, n_3649, n_4302, n_2514, n_4786, n_3257, n_1027, n_326, n_4160, n_2293, n_4051, n_2028, n_558, n_3009, n_1276, n_1412, n_3981, n_1199, n_352, n_1038, n_520, n_1841, n_154, n_2581, n_71, n_3224, n_4647, n_3752, n_870, n_1711, n_1891, n_434, n_3526, n_2546, n_965, n_3790, n_3491, n_935, n_817, n_1175, n_4613, n_4649, n_64, n_1888, n_1963, n_4795, n_2226, n_2891, n_4028, n_103, n_97, n_7, n_1690, n_3819, n_2449, n_431, n_1194, n_2297, n_4186, n_4731, n_1759, n_2177, n_3747, n_2227, n_4618, n_127, n_2190, n_3346, n_4742, n_2876, n_4099, n_452, n_3484, n_3620, n_1260, n_1746, n_2479, n_1464, n_4295, n_649, n_1444, n_4694, n_4533, n_3038, n_3068, n_2871, n_4244, n_4603, n_2943, n_4254, n_3143, n_3168, n_1680, n_4697, n_2607, n_3994, n_4190, n_4810, n_3317, n_1121, n_433, n_8, n_4391, n_949, n_3263, n_2582, n_4157, n_4283, n_4681, n_1001, n_1503, n_4638, n_1468, n_3455, n_3452, n_1510, n_1380, n_1994, n_1195, n_4707, n_2577, n_4527, n_2796, n_757, n_2342, n_106, n_4156, n_1851, n_4848, n_2937, n_3095, n_2805, n_1145, n_524, n_394, n_4918, n_1153, n_3856, n_741, n_2914, n_4898, n_1964, n_2869, n_4002, n_1163, n_1207, n_5010, n_2406, n_3623, n_2846, n_2925, n_3773, n_3918, n_2398, n_2857, n_4528, n_3932, n_4619, n_4673, n_940, n_3516, n_4822, n_2155, n_2516, n_3797, n_1596, n_2947, n_123, n_978, n_4299, n_4801, n_1474, n_1665, n_1269, n_3515, n_2886, n_267, n_2093, n_2473, n_1208, n_3287, n_3378, n_1431, n_4279, n_4769, n_4632, n_660, n_4294, n_1732, n_4125, n_4232, n_4949, n_374, n_2941, n_2457, n_4790, n_459, n_962, n_723, n_2536, n_1336, n_1758, n_2952, n_4847, n_3058, n_4365, n_1878, n_3505, n_4610, n_88, n_3730, n_4489, n_168, n_974, n_727, n_4967, n_957, n_4992, n_3001, n_303, n_3945, n_4542, n_2261, n_2729, n_3597, n_1612, n_2897, n_2077, n_4198, n_2909, n_4534, n_4500, n_5014, n_69, n_3185, n_1300, n_1127, n_3523, n_1785, n_2829, n_4597, n_4329, n_1006, n_4087, n_3811, n_1270, n_1664, n_3200, n_2231, n_2017, n_2604, n_4257, n_3453, n_322, n_2390, n_3213, n_1041, n_3077, n_1562, n_383, n_3474, n_3984, n_239, n_630, n_2151, n_55, n_2106, n_2716, n_4665, n_1913, n_1823, n_3679, n_3422, n_3888, n_4189, n_1875, n_1304, n_2803, n_1324, n_3707, n_1846, n_3429, n_1903, n_3849, n_3946, n_860, n_3229, n_4463, n_1805, n_429, n_4687, n_948, n_4670, n_4084, n_4703, n_4037, n_2922, n_83, n_3275, n_3499, n_2645, n_2727, n_560, n_340, n_3421, n_2240, n_2436, n_1552, n_3618, n_574, n_2593, n_3683, n_58, n_3642, n_3286, n_3808, n_824, n_359, n_1327, n_4763, n_1684, n_3590, n_366, n_815, n_4594, n_3424, n_1381, n_1037, n_2301, n_3583, n_3560, n_4076, n_4714, n_2419, n_3215, n_589, n_4776, n_2122, n_2512, n_4102, n_2786, n_3171, n_1437, n_645, n_238, n_3020, n_3677, n_3462, n_3468, n_1893, n_2910, n_222, n_1123, n_1467, n_2163, n_634, n_32, n_2254, n_1382, n_925, n_3546, n_424, n_2647, n_1311, n_1519, n_256, n_950, n_4443, n_4507, n_1811, n_2443, n_2624, n_3012, n_4575, n_380, n_419, n_3244, n_389, n_3130, n_3822, n_3569, n_912, n_136, n_86, n_968, n_4452, n_4348, n_619, n_376, n_4355, n_3494, n_515, n_351, n_885, n_2125, n_3771, n_683, n_3110, n_1057, n_1051, n_721, n_1157, n_3073, n_4572, n_22, n_802, n_4026, n_2265, n_4104, n_1608, n_4512, n_3554, n_38, n_4377, n_280, n_1305, n_3178, n_873, n_2334, n_690, n_33, n_4521, n_583, n_4488, n_2289, n_3051, n_302, n_1343, n_2783, n_2263, n_3750, n_2341, n_3632, n_4588, n_2733, n_1288, n_212, n_2785, n_2415, n_3299, n_4519, n_3715, n_972, n_3040, n_1938, n_1200, n_2499, n_3568, n_3737, n_1185, n_991, n_1967, n_576, n_1329, n_3255, n_4856, n_2997, n_4400, n_943, n_3326, n_3734, n_650, n_4778, n_286, n_2429, n_883, n_470, n_325, n_132, n_856, n_1793, n_4352, n_4441, n_918, n_4761, n_942, n_1804, n_189, n_4347, n_4095, n_3196, n_4593, n_2364, n_2533, n_3492, n_2780, n_4727, n_4568, n_195, n_2291, n_4043, n_1636, n_3601, n_1350, n_1865, n_2973, n_1096, n_2094, n_1575, n_2393, n_1697, n_3831, n_3801, n_225, n_2043, n_2751, n_192, n_4893, n_5032, n_1549, n_1934, n_4948, n_4000, n_655, n_3240, n_2025, n_1446, n_4406, n_2758, n_1458, n_472, n_1807, n_387, n_2618, n_398, n_2559, n_763, n_4748, n_2295, n_3931, n_1219, n_4010, n_2840, n_5017, n_1814, n_2822, n_4710, n_287, n_555, n_4607, n_4117, n_3636, n_1722, n_2441, n_1802, n_3083, n_4487, n_5001, n_2795, n_2981, n_2282, n_2800, n_4817, n_311, n_3380, n_2098, n_1296, n_3460, n_3409, n_3538, n_2068, n_4849, n_4867, n_445, n_2641, n_3198, n_1895, n_4728, n_588, n_789, n_4247, n_4933, n_107, n_4018, n_3900, n_1105, n_4902, n_4518, n_4409, n_4411, n_3872, n_4336, n_149, n_2270, n_4777, n_2653, n_836, n_2496, n_1908, n_2259, n_3877, n_458, n_2995, n_2494, n_3547, n_3977, n_1102, n_4052, n_3459, n_1499, n_4398, n_3155, n_2633, n_4954, n_2435, n_1392, n_1164, n_2097, n_4304, n_3911, n_1303, n_4431, n_4192, n_3736, n_4805, n_118, n_601, n_4885, n_253, n_1661, n_3565, n_172, n_4701, n_2575, n_861, n_1658, n_1904, n_1345, n_176, n_1899, n_1003, n_2067, n_2219, n_3533, n_2877, n_2148, n_393, n_4631, n_1726, n_3035, n_421, n_1657, n_768, n_1475, n_1725, n_1313, n_1136, n_1491, n_754, n_3639, n_708, n_735, n_2501, n_3079, n_4965, n_1915, n_1109, n_1310, n_2605, n_4747, n_1399, n_1979, n_193, n_2924, n_4111, n_808, n_2484, n_797, n_1025, n_4587, n_3731, n_2946, n_4538, n_435, n_766, n_541, n_1117, n_2754, n_687, n_1742, n_2489, n_536, n_2012, n_1291, n_4094, n_3503, n_2866, n_3561, n_1155, n_1418, n_1011, n_2917, n_2425, n_3536, n_3661, n_4150, n_827, n_4878, n_1703, n_1650, n_1137, n_3934, n_4985, n_3922, n_3846, n_318, n_2103, n_653, n_2160, n_2498, n_2697, n_850, n_3074, n_1999, n_2372, n_3673, n_3768, n_1372, n_2861, n_605, n_2630, n_3943, n_353, n_2430, n_493, n_2433, n_3293, n_4022, n_1531, n_840, n_1334, n_4852, n_2528, n_4869, n_4700, n_4035, n_2316, n_1898, n_3294, n_4426, n_554, n_3415, n_2284, n_2817, n_3139, n_2598, n_4601, n_2687, n_1120, n_198, n_1890, n_714, n_4220, n_1944, n_909, n_1497, n_3431, n_3169, n_3151, n_2078, n_3284, n_3070, n_4066, n_119, n_2884, n_4515, n_4351, n_3126, n_4403, n_1981, n_1663, n_1718, n_4509, n_4858, n_3700, n_509, n_147, n_1518, n_4223, n_1281, n_1889, n_209, n_1489, n_5025, n_2966, n_1376, n_2326, n_1569, n_2188, n_186, n_756, n_1429, n_4644, n_4456, n_399, n_2448, n_4346, n_3170, n_2748, n_3311, n_3272, n_2898, n_2717, n_1861, n_760, n_3628, n_3691, n_220, n_4235, n_1867, n_1945, n_3018, n_481, n_2573, n_4435, n_2939, n_3807, n_271, n_2447, n_4764, n_886, n_1221, n_167, n_2774, n_1707, n_853, n_4655, n_3161, n_377, n_4581, n_751, n_4827, n_2488, n_392, n_3477, n_2476, n_704, n_4399, n_2781, n_2778, n_771, n_4782, n_1520, n_4363, n_2887, n_1287, n_4864, n_1262, n_2691, n_1411, n_3054, n_4335, n_2526, n_2703, n_2167, n_3391, n_4259, n_56, n_2709, n_816, n_1536, n_4865, n_4056, n_1344, n_4564, n_1246, n_3840, n_1339, n_3518, n_2956, n_3733, n_328, n_2173, n_1842, n_871, n_3738, n_685, n_78, n_3464, n_2018, n_4526, n_1555, n_3245, n_4417, n_499, n_98, n_402, n_4899, n_796, n_2119, n_1502, n_2157, n_2552, n_1012, n_1, n_2453, n_4798, n_1525, n_740, n_3509, n_3352, n_3076, n_3535, n_2182, n_277, n_1061, n_3251, n_92, n_2931, n_1193, n_3118, n_3511, n_1226, n_3443, n_2146, n_1487, n_3644, n_3336, n_3935, n_781, n_542, n_3521, n_3562, n_3948, n_4750, n_1515, n_2918, n_3232, n_1673, n_27, n_2112, n_1739, n_2958, n_3114, n_3125, n_4981, n_2394, n_3612, n_2954, n_4835, n_4430, n_4081, n_1103, n_3132, n_4407, n_648, n_312, n_3951, n_4894, n_3238, n_3210, n_2036, n_3267, n_4995, n_480, n_425, n_695, n_37, n_3964, n_3772, n_229, n_1956, n_437, n_1642, n_2279, n_3373, n_4446, n_3884, n_0, n_3726, n_805, n_2525, n_2892, n_113, n_2907, n_3577, n_2820, n_269, n_2049, n_2273, n_2719, n_1741, n_1160, n_4057, n_4332, n_1258, n_4314, n_1074, n_3347, n_3216, n_1621, n_3809, n_2113, n_1448, n_4288, n_3567, n_1634, n_3939, n_4241, n_3321, n_3212, n_666, n_1433, n_2256, n_3152, n_319, n_2920, n_4265, n_1186, n_1018, n_2247, n_713, n_1622, n_166, n_1180, n_3705, n_2802, n_4705, n_3159, n_2268, n_3778, n_3304, n_1378, n_3912, n_1729, n_2739, n_469, n_2771, n_4604, n_549, n_3795, n_5020, n_4419, n_4477, n_3179, n_3256, n_667, n_2386, n_1501, n_3086, n_1007, n_2369, n_2927, n_4217, n_4395, n_2821, n_1099, n_2568, n_564, n_1738, n_3728, n_21, n_3064, n_3088, n_1021, n_4639, n_3713, n_3663, n_3246, n_2495, n_1535, n_1789, n_819, n_2302, n_951, n_247, n_1494, n_292, n_625, n_2069, n_417, n_3434, n_1806, n_933, n_1563, n_4227, n_26, n_4033, n_4289, n_2024, n_4780, n_755, n_4243, n_4982, n_530, n_4330, n_3695, n_556, n_2482, n_2677, n_3832, n_3987, n_902, n_4991, n_579, n_1698, n_2329, n_1098, n_2142, n_320, n_3332, n_1135, n_3048, n_3937, n_2203, n_4525, n_1243, n_101, n_3782, n_2978, n_2058, n_2458, n_4208, n_3786, n_371, n_2888, n_3638, n_1236, n_1633, n_4177, n_3763, n_2669, n_1778, n_2306, n_3022, n_4264, n_335, n_3087, n_3489, n_2566, n_343, n_308, n_2149, n_1078, n_3060, n_4276, n_3013, n_1984, n_2408, n_1877, n_3049, n_1723, n_339, n_4485, n_183, n_4626, n_1036, n_1097, n_347, n_798, n_2659, n_1414, n_290, n_4975, n_1852, n_578, n_344, n_3089, n_422, n_2470, n_3985, n_496, n_1391, n_670, n_4760, n_4652, n_4624, n_48, n_663, n_2551, n_1587, n_2682, n_813, n_1284, n_3440, n_1748, n_4569, n_2699, n_4897, n_888, n_2769, n_3542, n_3436, n_2615, n_3940, n_446, n_1064, n_858, n_2985, n_691, n_2753, n_363, n_1582, n_3637, n_2842, n_4523, n_1836, n_2868, n_3141, n_3164, n_3570, n_4919, n_4025, n_461, n_2712, n_3936, n_4503, n_3507, n_3821, n_2700, n_1211, n_3367, n_4464, n_907, n_3096, n_3496, n_4114, n_989, n_2544, n_2356, n_488, n_892, n_4556, n_2620, n_1581, n_4089, n_586, n_2919, n_4327, n_230, n_953, n_4218, n_2150, n_3146, n_2241, n_2757, n_963, n_1052, n_954, n_478, n_4353, n_2042, n_534, n_884, n_1754, n_1623, n_2921, n_2720, n_1854, n_4990, n_1856, n_143, n_4959, n_4161, n_237, n_832, n_1319, n_3992, n_2616, n_1906, n_4103, n_1387, n_4466, n_2262, n_2462, n_1532, n_18, n_3625, n_1156, n_794, n_2798, n_2945, n_2331, n_686, n_2837, n_847, n_4844, n_2979, n_3655, n_4688, n_4765, n_702, n_2548, n_822, n_2108, n_3640, n_4388, n_4206, n_1538, n_1779, n_4738, n_53, n_1369, n_3909, n_3207, n_3944, n_809, n_4434, n_4837, n_3042, n_1942, n_2510, n_4219, n_2804, n_3659, n_2120, n_411, n_414, n_5012, n_1293, n_1876, n_4620, n_36, n_1810, n_2813, n_4438, n_2009, n_2222, n_3510, n_28, n_3218, n_2667, n_11, n_3150, n_747, n_52, n_4325, n_1733, n_2413, n_615, n_851, n_843, n_705, n_3775, n_4133, n_678, n_4184, n_2518, n_2629, n_367, n_4481, n_3416, n_4379, n_2181, n_1829, n_547, n_4030, n_116, n_4490, n_3138, n_4397, n_1710, n_1128, n_2928, n_1734, n_4820, n_590, n_3770, n_1308, n_4938, n_4179, n_3469, n_372, n_677, n_2723, n_314, n_368, n_3220, n_4641, n_2539, n_100, n_3855, n_1008, n_2054, n_1559, n_4931, n_1765, n_3158, n_1744, n_2623, n_1617, n_295, n_133, n_3113, n_2718, n_3760, n_4078, n_1760, n_568, n_39, n_2856, n_1832, n_4146, n_4360, n_3666, n_3828, n_93, n_3288, n_4404, n_1509, n_1874, n_4787, n_2060, n_2613, n_1987, n_3667, n_878, n_1306, n_3703, n_4903, n_3558, n_2545, n_2787, n_906, n_919, n_4356, n_658, n_2061, n_4432, n_2378, n_1740, n_1586, n_4291, n_535, n_4386, n_9, n_4149, n_1492, n_592, n_1692, n_2982, n_2481, n_3545, n_2507, n_4019, n_2900, n_1095, n_1614, n_2339, n_457, n_4637, n_603, n_4935, n_4785, n_3426, n_3454, n_3820, n_3741, n_3410, n_2029, n_995, n_1609, n_396, n_1887, n_4413, n_1073, n_2346, n_662, n_3990, n_4493, n_218, n_3475, n_1215, n_1592, n_2882, n_1721, n_2338, n_3672, n_3197, n_3109, n_2721, n_1043, n_486, n_3002, n_337, n_3897, n_1159, n_3845, n_2081, n_299, n_4570, n_2156, n_4296, n_1820, n_5019, n_2418, n_2179, n_1416, n_1724, n_2521, n_3458, n_1420, n_1132, n_3330, n_4606, n_4774, n_2477, n_3887, n_4093, n_1486, n_4672, n_3519, n_4174, n_3374, n_3045, n_1870, n_309, n_2367, n_4766, n_84, n_2896, n_652, n_1365, n_4074, n_4600, n_1927, n_1349, n_4460, n_288, n_1031, n_3645, n_3223, n_3929, n_834, n_2255, n_2272, n_893, n_1965, n_1902, n_1941, n_3938, n_2878, n_504, n_874, n_3498, n_2015, n_1982, n_4110, n_3189, n_2066, n_993, n_3154, n_1551, n_545, n_450, n_2905, n_3965, n_3566, n_1217, n_2220, n_4349, n_628, n_3788, n_2410, n_4313, n_1084, n_970, n_1935, n_3366, n_1534, n_1351, n_2696, n_4863, n_1205, n_3242, n_495, n_3525, n_3486, n_2405, n_3995, n_2088, n_2953, n_4036, n_921, n_1795, n_2578, n_3483, n_128, n_1821, n_3894, n_3478, n_4015, n_3890, n_2740, n_2656, n_1080, n_1274, n_3524, n_5034, n_1708, n_426, n_562, n_1436, n_3549, n_1691, n_2092, n_2075, n_3658, n_1776, n_4807, n_2281, n_2131, n_3026, n_1757, n_890, n_1919, n_960, n_4230, n_3419, n_1290, n_1047, n_2053, n_1958, n_1252, n_348, n_3784, n_2969, n_3941, n_2864, n_3195, n_3190, n_1553, n_3678, n_2664, n_3456, n_444, n_1808, n_316, n_2266, n_2650, n_4428, n_146, n_5003, n_408, n_967, n_2731, n_3953, n_3166, n_4122, n_3976, n_1357, n_3979, n_4582, n_2998, n_4684, n_4840, n_3162, n_983, n_2760, n_3377, n_3749, n_3962, n_1826, n_2304, n_762, n_1283, n_17, n_2637, n_4384, n_4423, n_4096, n_2881, n_1203, n_3282, n_821, n_1763, n_3231, n_1966, n_321, n_4996, n_621, n_2475, n_4598, n_4478, n_507, n_2646, n_1605, n_1228, n_3920, n_4890, n_5027, n_3203, n_3866, n_2903, n_3921, n_828, n_779, n_4106, n_3717, n_2743, n_2675, n_1439, n_3052, n_945, n_3743, n_1932, n_4721, n_984, n_694, n_1983, n_4029, n_1594, n_900, n_3870, n_4496, n_3529, n_1147, n_1977, n_2153, n_13, n_4338, n_3094, n_2310, n_3952, n_2287, n_2860, n_2056, n_1470, n_1735, n_2318, n_833, n_2502, n_2504, n_4495, n_4762, n_2974, n_2901, n_1940, n_2793, n_3442, n_1201, n_1114, n_3998, n_2285, n_3147, n_4141, n_669, n_1176, n_1149, n_1020, n_211, n_1824, n_1917, n_3386, n_4107, n_3, n_4667, n_2325, n_178, n_2446, n_3488, n_1035, n_4547, n_2893, n_2588, n_2962, n_4004, n_661, n_4668, n_4953, n_3898, n_849, n_584, n_1786, n_50, n_430, n_4997, n_4274, n_2627, n_4759, n_1413, n_801, n_4467, n_2080, n_2377, n_2340, n_3552, n_875, n_357, n_3684, n_4735, n_3137, n_165, n_2361, n_1173, n_1603, n_969, n_1401, n_4113, n_1019, n_1998, n_4686, n_304, n_3759, n_4321, n_4342, n_2034, n_3933, n_3206, n_3966, n_1702, n_4183, n_778, n_1122, n_4068, n_4872, n_4233, n_3192, n_3764, n_4709, n_5038, n_2649, n_1187, n_1929, n_2807, n_2542, n_2313, n_489, n_1174, n_3324, n_3914, n_4625, n_2558, n_2063, n_3803, n_3742, n_2252, n_4819, n_1685, n_917, n_1714, n_1541, n_2576, n_4900, n_3390, n_1573, n_3746, n_2373, n_1713, n_3817, n_2745, n_1253, n_210, n_1737, n_774, n_2493, n_4930, n_1059, n_1133, n_4537, n_2885, n_5011, n_3318, n_4070, n_4282, n_3485, n_4180, n_665, n_3839, n_1440, n_3333, n_2845, n_4143, n_4659, n_2602, n_205, n_4579, n_4616, n_1496, n_1125, n_3014, n_2547, n_5023, n_1812, n_4105, n_232, n_2532, n_3791, n_2665, n_3905, n_427, n_3368, n_3530, n_1930, n_1955, n_2765, n_3329, n_2994, n_2401, n_3135, n_2003, n_1457, n_4895, n_3573, n_3148, n_2264, n_3534, n_1482, n_4275, n_1266, n_3970, n_3438, n_4098, n_872, n_594, n_200, n_1297, n_4789, n_1972, n_2806, n_1184, n_2184, n_985, n_3217, n_3404, n_3425, n_4055, n_2926, n_626, n_3540, n_3670, n_3973, n_2023, n_3249, n_2351, n_676, n_4442, n_4698, n_642, n_1602, n_194, n_1178, n_4779, n_2286, n_4966, n_503, n_2065, n_4017, n_3397, n_3740, n_620, n_1081, n_4418, n_2549, n_2705, n_2332, n_703, n_1318, n_780, n_2977, n_1454, n_3723, n_1227, n_3600, n_245, n_4134, n_1388, n_2836, n_672, n_581, n_1625, n_2130, n_898, n_3239, n_2773, n_3365, n_3476, n_3686, n_4913, n_1452, n_265, n_443, n_1791, n_2850, n_1747, n_4251, n_1817, n_3982, n_2654, n_4621, n_1326, n_3176, n_4559, n_2186, n_4368, n_4740, n_5007, n_3581, n_2562, n_4077, n_67, n_4642, n_1192, n_2221, n_1024, n_3576, n_1792, n_1564, n_1868, n_1613, n_4049, n_941, n_3862, n_68, n_3495, n_3879, n_2348, n_4724, n_1238, n_1772, n_282, n_752, n_1476, n_1108, n_2818, n_1100, n_3646, n_2129, n_3345, n_1395, n_4546, n_862, n_3584, n_3756, n_381, n_2889, n_390, n_5021, n_2772, n_1675, n_1924, n_4382, n_1554, n_3999, n_42, n_2844, n_2138, n_2260, n_1813, n_4833, n_3056, n_2345, n_1172, n_379, n_428, n_1341, n_3295, n_2382, n_4719, n_4178, n_3062, n_2317, n_3289, n_1973, n_786, n_1142, n_2579, n_1770, n_138, n_4228, n_4401, n_1756, n_1716, n_2788, n_2984, n_3364, n_1873, n_3201, n_221, n_622, n_1087, n_3472, n_2874, n_4605, n_4877, n_3235, n_4968, n_1272, n_104, n_5030, n_3949, n_3543, n_1247, n_591, n_3050, n_313, n_1478, n_3903, n_4834, n_1210, n_1364, n_2183, n_2742, n_3314, n_4158, n_2360, n_3254, n_369, n_4171, n_4045, n_598, n_1367, n_4562, n_3634, n_1460, n_2834, n_2531, n_517, n_413, n_5015, n_2702, n_2030, n_903, n_3115, n_4749, n_203, n_4390, n_4979, n_1404, n_1794, n_2234, n_4804, n_2209, n_4270, n_2797, n_1255, n_79, n_2321, n_722, n_3680, n_844, n_201, n_3497, n_40, n_1601, n_2940, n_2612, n_1495, n_4566, n_979, n_2841, n_3322, n_4576, n_846, n_2427, n_2505, n_76, n_4061, n_2070, n_3250, n_585, n_270, n_2594, n_1914, n_2335, n_2904, n_4767, n_4328, n_3004, n_3112, n_2349, n_1379, n_3874, n_4676, n_4544, n_2170, n_1091, n_641, n_3175, n_3522, n_4429, n_575, n_4591, n_3266, n_4646, n_1130, n_4563, n_4725, n_2210, n_4169, n_3247, n_3091, n_3066, n_246, n_2426, n_657, n_4320, n_4881, n_491, n_160, n_566, n_565, n_3613, n_3444, n_1181, n_1505, n_4012, n_651, n_4636, n_4584, n_807, n_3910, n_4711, n_835, n_3319, n_3335, n_99, n_3413, n_1969, n_4680, n_2044, n_1138, n_927, n_2689, n_3259, n_4191, n_4293, n_2010, n_3688, n_3016, n_1693, n_2599, n_904, n_3338, n_3414, n_1827, n_4671, n_4209, n_1271, n_1542, n_1423, n_1166, n_1751, n_1508, n_82, n_785, n_2200, n_3261, n_5026, n_1161, n_3863, n_3027, n_2746, n_1150, n_3127, n_226, n_1780, n_3732, n_4250, n_1055, n_3596, n_4699, n_111, n_3906, n_4127, n_880, n_3297, n_544, n_155, n_2683, n_1370, n_1360, n_2388, n_4292, n_3641, n_4577, n_4854, n_105, n_4202, n_5000, n_2853, n_1323, n_688, n_3766, n_1353, n_800, n_2880, n_1666, n_3350, n_2389, n_4165, n_4866, n_4038, n_4109, n_915, n_864, n_1264, n_447, n_4412, n_3407, n_3599, n_3621, n_1580, n_2244, n_3815, n_2257, n_497, n_1607, n_2538, n_2105, n_2, n_3163, n_1118, n_1686, n_947, n_373, n_3710, n_307, n_4155, n_1359, n_2031, n_3891, n_1230, n_4144, n_375, n_2165, n_929, n_3379, n_4374, n_3532, n_1124, n_1818, n_2127, n_1576, n_1104, n_1294, n_51, n_1257, n_1182, n_3531, n_2963, n_3834, n_4548, n_3258, n_24, n_4989, n_4622, n_1016, n_4315, n_2959, n_2047, n_1845, n_240, n_2193, n_2478, n_4816, n_231, n_1483, n_2983, n_227, n_3810, n_1289, n_94, n_2715, n_2085, n_1669, n_370, n_4483, n_2782, n_1670, n_2672, n_2651, n_4358, n_3656, n_2071, n_2561, n_2643, n_1374, n_4793, n_4168, n_3446, n_955, n_3028, n_4806, n_1146, n_4350, n_550, n_897, n_1428, n_1216, n_3836, n_3963, n_1872, n_3389, n_1931, n_4187, n_1070, n_4166, n_1030, n_3222, n_1071, n_1267, n_1801, n_1513, n_2970, n_2235, n_673, n_837, n_4937, n_3980, n_2791, n_680, n_1473, n_3755, n_4258, n_4498, n_1590, n_2174, n_2714, n_3563, n_2506, n_675, n_4064, n_4936, n_1556, n_184, n_1863, n_3841, n_114, n_2118, n_4770, n_2944, n_881, n_2407, n_4907, n_468, n_129, n_3262, n_1450, n_5018, n_4006, n_4861, n_1322, n_3690, n_889, n_2358, n_973, n_3716, n_1700, n_2833, n_4712, n_477, n_3191, n_3837, n_3193, n_1971, n_3252, n_2275, n_2855, n_3273, n_3544, n_4310, n_1523, n_1950, n_1447, n_2370, n_3954, n_3025, n_4674, n_4908, n_736, n_2750, n_3899, n_1278, n_4159, n_3714, n_49, n_3071, n_3739, n_593, n_4069, n_12, n_2784, n_3718, n_3092, n_3470, n_4862, n_2557, n_1248, n_70, n_289, n_4850, n_3781, n_4813, n_4912, n_2590, n_2330, n_2942, n_3106, n_1882, n_3328, n_944, n_3889, n_4256, n_4224, n_3508, n_4024, n_2218, n_2267, n_857, n_2636, n_1825, n_1951, n_1883, n_2759, n_4415, n_4702, n_4252, n_4457, n_971, n_117, n_404, n_1393, n_2319, n_596, n_3481, n_2808, n_2676, n_1709, n_2679, n_4491, n_266, n_2930, n_1838, n_3514, n_2777, n_2434, n_4132, n_2660, n_2611, n_4261, n_1660, n_4886, n_4090, n_2529, n_2698, n_1662, n_1481, n_4001, n_3047, n_868, n_2454, n_4371, n_914, n_4473, n_3120, n_4007, n_1743, n_4268, n_5028, n_1479, n_4480, n_2350, n_3895, n_4194, n_759, n_4824, n_1892, n_4120, n_4427, n_3745, n_806, n_2990, n_1766, n_324, n_1571, n_3119, n_4142, n_1189, n_4082, n_3479, n_4085, n_4073, n_4260, n_1649, n_4163, n_4439, n_2064, n_3867, n_4372, n_3500, n_3279, n_2621, n_5024, n_523, n_1537, n_4262, n_2671, n_1798, n_1790, n_4720, n_525, n_1647, n_4685, n_2563, n_43, n_2387, n_4334, n_1674, n_1830, n_2073, n_4511, n_139, n_4014, n_3144, n_4757, n_2913, n_2336, n_254, n_1233, n_1615, n_4175, n_2005, n_526, n_1916, n_293, n_244, n_4648, n_47, n_1333, n_5006, n_1443, n_946, n_1539, n_4892, n_3823, n_1866, n_4173, n_689, n_738, n_1624, n_4970, n_640, n_3816, n_1279, n_4108, n_4486, n_610, n_2960, n_1090, n_633, n_439, n_4627, n_758, n_2290, n_2045, n_3369, n_3783, n_2040, n_3199, n_3843, n_1049, n_2145, n_1639, n_1068, n_3030, n_2580, n_3685, n_4249, n_122, n_331, n_10, n_2039, n_4961, n_90, n_3753, n_2035, n_4718, n_3555, n_3579, n_2509, n_3236, n_4317, n_1362, n_4855, n_3969, n_2459, n_4154, n_152, n_3396, n_1445, n_4023, n_4420, n_1923, n_1017, n_2116, n_1434, n_1054, n_1828, n_2320, n_1045, n_2038, n_2137, n_4973, n_4640, n_2583, n_484, n_1033, n_4396, n_636, n_4367, n_2087, n_1009, n_109, n_454, n_1989, n_3818, n_2523, n_255, n_4387, n_4951, n_4453, n_4170, n_1578, n_3719, n_1959, n_3681, n_2737, n_1574, n_2399, n_4308, n_2812, n_473, n_2355, n_2133, n_1426, n_3830, n_2585, n_2725, n_614, n_3883, n_1355, n_2565, n_4152, n_773, n_208, n_142, n_743, n_4392, n_4660, n_3149, n_296, n_3268, n_4281, n_65, n_4661, n_4200, n_3614, n_2111, n_3301, n_3466, n_4962, n_1237, n_2595, n_761, n_3411, n_4958, n_329, n_4271, n_3586, n_1390, n_30, n_4071, n_4921, n_130, n_1980, n_3065, n_4361, n_1093, n_263, n_4614, n_1265, n_44, n_224, n_2681, n_3103, n_765, n_4945, n_2424, n_4922, n_4732, n_1015, n_1651, n_2775, n_4693, n_511, n_358, n_1101, n_77, n_1106, n_4326, n_3557, n_2230, n_4744, n_2851, n_4305, n_174, n_1455, n_767, n_2490, n_1407, n_441, n_4213, n_2849, n_3692, n_2204, n_365, n_4929, n_729, n_1961, n_4964, n_911, n_1430, n_4802, n_513, n_1354, n_4139, n_1044, n_3029, n_2508, n_4031, n_2416, n_623, n_3881, n_2461, n_490, n_2243, n_4583, n_233, n_572, n_4210, n_4666, n_2929, n_3751, n_2555, n_2662, n_1611, n_2368, n_2890, n_2554, n_3698, n_3927, n_1082, n_1840, n_4540, n_3961, n_716, n_1630, n_4891, n_391, n_701, n_1023, n_539, n_803, n_1092, n_3559, n_2661, n_2572, n_3993, n_4940, n_1056, n_3588, n_2308, n_4590, n_4830, n_4664, n_3860, n_1029, n_1206, n_3160, n_2191, n_2428, n_3847, n_4946, n_1346, n_4906, n_2158, n_3290, n_4663, n_1060, n_2824, n_3033, n_3298, n_248, n_2440, n_4883, n_1386, n_2923, n_1442, n_4162, n_3665, n_74, n_3264, n_2333, n_2916, n_483, n_4297, n_1632, n_1085, n_1066, n_3800, n_2403, n_4608, n_46, n_2792, n_2870, n_3991, n_378, n_1112, n_3134, n_4172, n_4791, n_4536, n_2463, n_4773, n_4497, n_2472, n_4611, n_4755, n_1768, n_2294, n_4960, n_455, n_2993, n_1719, n_3864, n_385, n_4658, n_2732, n_2309, n_2948, n_1560, n_4362, n_4306, n_2123, n_3209, n_3504, n_2037, n_2685, n_1953, n_4422, n_2589, n_1301, n_1363, n_3482, n_2233, n_1312, n_804, n_537, n_4555, n_2827, n_153, n_1504, n_3956, n_3572, n_250, n_992, n_4215, n_4280, n_3375, n_4047, n_260, n_842, n_2082, n_1643, n_3167, n_3423, n_2362, n_2609, n_1976, n_2223, n_3044, n_3854, n_2468, n_1610, n_1077, n_1422, n_3078, n_540, n_323, n_894, n_3253, n_4027, n_831, n_2280, n_4599, n_3363, n_4812, n_1511, n_234, n_3689, n_2020, n_4628, n_1881, n_988, n_2749, n_3451, n_4873, n_4657, n_2971, n_2311, n_3950, n_4458, n_4121, n_1616, n_4476, n_2298, n_4756, n_3869, n_4307, n_4860, n_4359, n_635, n_2303, n_2810, n_2747, n_1848, n_2126, n_4573, n_4118, n_4803, n_4079, n_15, n_4091, n_681, n_1638, n_2002, n_3712, n_2371, n_2935, n_830, n_3085, n_1655, n_749, n_2574, n_1134, n_1358, n_717, n_4316, n_939, n_3697, n_482, n_1232, n_734, n_2638, n_4044, n_4062, n_4524, n_4843, n_3971, n_1338, n_2016, n_1522, n_2949, n_2711, n_338, n_1653, n_1506, n_14, n_990, n_2867, n_1894, n_975, n_2794, n_567, n_3145, n_3124, n_4253, n_151, n_2608, n_2657, n_770, n_2852, n_2392, n_711, n_85, n_3517, n_1441, n_3100, n_2522, n_1834, n_3758, n_3356, n_2835, n_617, n_1572, n_1968, n_3269, n_1516, n_3506, n_1736, n_3605, n_2409, n_3402, n_217, n_4679, n_4115, n_726, n_4998, n_2988, n_1731, n_818, n_1970, n_2766, n_2201, n_2117, n_4167, n_1993, n_3835, n_2205, n_1335, n_1777, n_1957, n_3967, n_5016, n_1912, n_3401, n_3226, n_1410, n_707, n_3902, n_4730, n_937, n_2779, n_1584, n_487, n_3654, n_2164, n_2115, n_2232, n_1302, n_1774, n_4713, n_2811, n_3348, n_179, n_410, n_895, n_3358, n_2121, n_1803, n_4204, n_1543, n_1991, n_2224, n_732, n_4743, n_500, n_1067, n_3805, n_3825, n_148, n_3657, n_4924, n_3928, n_4859, n_2692, n_538, n_2008, n_4654, n_799, n_1213, n_4733, n_3792, n_4272, n_3974, n_3871, n_1753, n_2283, n_3278, n_89, n_1689, n_4269, n_4695, n_1855, n_869, n_401, n_3312, n_1352, n_2197, n_2199, n_3285, n_137, n_294, n_3968, n_2228, n_4704, n_4551, n_684, n_124, n_268, n_2421, n_2902, n_4957, n_664, n_2480, n_235, n_2363, n_643, n_4072, n_916, n_1115, n_4781, n_3606, n_5004, n_2550, n_467, n_4424, n_823, n_725, n_3055, n_3711, n_3315, n_3172, n_3292, n_4436, n_3878, n_4450, n_3553, n_719, n_4746, n_1683, n_1530, n_997, n_932, n_3131, n_1409, n_3850, n_788, n_4459, n_1268, n_2996, n_559, n_508, n_1320, n_4050, n_986, n_2315, n_3228, n_1317, n_2102, n_1063, n_4853, n_981, n_867, n_2422, n_134, n_2239, n_587, n_2950, n_3852, n_548, n_812, n_4520, n_518, n_2057, n_4008, n_905, n_782, n_3858, n_1901, n_4502, n_3032, n_4851, n_1330, n_31, n_3072, n_3081, n_3313, n_2710, n_1745, n_3924, n_769, n_4571, n_2006, n_934, n_1618, n_826, n_2343, n_3439, n_654, n_2535, n_4205, n_2726, n_570, n_4723, n_2799, n_4454, n_4229, n_1083, n_4739, n_2376, n_3017, n_787, n_2456, n_3904, n_2678, n_95, n_4838, n_2872, n_2451, n_522, n_4879, n_930, n_181, n_3926, n_1962, n_3996, n_4221, n_1577, n_2854, n_386, n_1701, n_4181, n_1550, n_2764, n_1498, n_4225, n_682, n_141, n_2567, n_3102, n_922, n_1648, n_4153, n_3627, n_4300, n_3551, n_432, n_1769, n_4783, n_839, n_2964, n_3769, n_2673, n_4530, n_4267, n_140, n_2292, n_3865, n_3859, n_3722, n_2442, n_928, n_1943, n_3117, n_3428, n_2961, n_3351, n_3527, n_236, n_1396, n_1348, n_2883, n_1752, n_4182, n_80, n_2912, n_35, n_1315, n_4825, n_4440, n_4549, n_1910, n_3955, n_462, n_4565, n_4039, n_3227, n_3300, n_4303, n_4574, n_471, n_4839, n_1028, n_4016, n_474, n_3435, n_3575, n_1546, n_595, n_632, n_4231, n_3165, n_4923, n_3652, n_4097, n_170, n_161, n_4083, n_1937, n_81, n_4461, n_3234, n_745, n_2381, n_3303, n_1654, n_3916, n_2569, n_3556, n_4101, n_2196, n_3591, n_4273, n_3024, n_3512, n_4939, n_4389, n_3930, n_4448, n_1325, n_1595, n_2161, n_2404, n_2083, n_2503, n_1540, n_1936, n_2027, n_453, n_403, n_2642, n_720, n_2500, n_1918, n_863, n_4831, n_2513, n_2695, n_3480, n_3057, n_3194, n_2414, n_1402, n_3662, n_4319, n_644, n_2229, n_1397, n_4596, n_2004, n_251, n_3694, n_2586, n_4726, n_1398, n_1879, n_4751, n_4222, n_1196, n_2274, n_2972, n_3225, n_334, n_811, n_175, n_4119, n_3799, n_4298, n_4474, n_1089, n_1004, n_242, n_2511, n_1681, n_3383, n_3585, n_2975, n_438, n_5029, n_2704, n_4214, n_4884, n_533, n_4366, n_1251, n_4009, n_278, n_4580, n_1263, n_611, n_1126, n_4129, n_4871, n_2617, n_4999, n_1859, n_1677, n_2955, n_4112, n_4337, n_4138, n_552, n_1528, n_1292, n_2520, n_1198, n_956, n_423, n_2134, n_4236, n_2185, n_3270, n_2143, n_5002, n_3595, n_1347, n_4238, n_1451, n_1022, n_1545, n_2374, n_173, n_859, n_1947, n_2114, n_3571, n_854, n_1799, n_2396, n_4734, n_674, n_1939, n_2486, n_516, n_4635, n_1152, n_3501, n_1869, n_4013, n_606, n_3039, n_275, n_2011, n_4242, n_6, n_4984, n_3851, n_2543, n_150, n_3036, n_1896, n_3180, n_191, n_1705, n_659, n_4561, n_2639, n_3325, n_3107, n_4021, n_3880, n_1261, n_938, n_3186, n_4955, n_1154, n_4501, n_3696, n_406, n_546, n_1280, n_3650, n_291, n_2761, n_257, n_3157, n_709, n_2537, n_2144, n_920, n_2515, n_2466, n_2652, n_2635, n_4197, n_4829, n_976, n_1949, n_1946, n_2936, n_775, n_1484, n_1328, n_4715, n_2141, n_4369, n_4543, n_2099, n_4941, n_1831, n_1598, n_4394, n_1850, n_163, n_243, n_1749, n_59, n_3101, n_3669, n_215, n_350, n_196, n_2663, n_1394, n_580, n_2693, n_3798, n_4065, n_4944, n_926, n_2180, n_2249, n_4135, n_1218, n_2632, n_475, n_1547, n_777, n_1755, n_415, n_485, n_958, n_2908, n_3744, n_4263, n_1862, n_1239, n_2915, n_2300, n_3291, n_4716, n_4942, n_164, n_2432, n_1521, n_3405, n_214, n_4745, n_2337, n_1167, n_1384, n_3907, n_923, n_4629, n_213, n_2932, n_2980, n_464, n_1069, n_3306, n_1784, n_4857, n_3136, n_4080, n_4226, n_4741, n_2101, n_1471, n_1986, n_4752, n_1750, n_1459, n_460, n_3986, n_4376, n_4753, n_571, n_4552, n_3885, n_2713, n_2644, n_1197, n_2951, n_3008, n_3709, n_1039, n_2214, n_34, n_2055, n_3427, n_4067, n_1403, n_4042, n_4176, n_4385, n_3320, n_5009, n_2688, n_1202, n_1463, n_3651, n_4333, n_3359, n_2865, n_349, n_2706, n_3676, n_4375, n_4788, n_4717, n_4986, n_3789, n_2152, n_3598, n_627, n_4815, n_4246, n_3580, n_2139, n_4609, n_91, n_2674, n_1565, n_4088, n_3682, n_4357, n_3371, n_1809, n_4462, n_4472, n_647, n_3433, n_1072, n_2305, n_2450, n_561, n_3447, n_3305, n_4148, n_4151, n_1712, n_3528, n_4373, n_4934, n_2322, n_2271, n_2625, n_4630, n_4643, n_4331, n_3989, n_4475, n_4846, n_3804, n_4344, n_1775, n_3296, n_1368, n_2762, n_4683, n_728, n_1162, n_272, n_1847, n_2767, n_2603, n_3116, n_1884, n_3602, n_2967, n_409, n_887, n_1905, n_2553, n_3706, n_2195, n_300, n_3923, n_931, n_599, n_4696, n_2626, n_3441, n_1978, n_1544, n_639, n_1629, n_2801, n_4011, n_4905, n_121, n_2763, n_360, n_2825, n_3643, n_4876, n_1997, n_3748, n_1477, n_3142, n_4278, n_1635, n_4623, n_187, n_4910, n_2690, n_4410, n_3370, n_2215, n_1259, n_4553, n_706, n_746, n_784, n_3978, n_110, n_4809, n_1244, n_1925, n_3660, n_1815, n_1788, n_2491, n_913, n_3833, n_865, n_61, n_697, n_1222, n_75, n_1679, n_4841, n_776, n_2022, n_3814, n_1415, n_2592, n_2838, n_4842, n_4911, n_4340, n_3513, n_3133, n_4645, n_1191, n_2992, n_3725, n_1833, n_4920, n_4972, n_2517, n_284, n_3128, n_744, n_629, n_2631, n_2178, n_1767, n_23, n_1529, n_2469, n_3355, n_604, n_2007, n_3917, n_3942, n_2736, n_3765, n_498, n_3000, n_252, n_624, n_1010, n_1231, n_739, n_1406, n_3108, n_3111, n_1837, n_1839, n_4557, n_4451, n_2875, n_936, n_1500, n_3844, n_3280, n_4054, n_3471, n_259, n_448, n_999, n_3205, n_2046, n_2848, n_2741, n_3003, n_3610, n_1933, n_1656, n_3564, n_1158, n_3988, n_563, n_3457, n_204, n_1678, n_4324, n_4821, n_1871, n_3630, n_3271, n_4771, n_908, n_4086, n_2412, n_4814, n_724, n_1781, n_2084, n_3648, n_3075, n_3173, n_4692, n_456, n_959, n_3031, n_3701, n_1773, n_3243, n_1169, n_45, n_2666, n_3385, n_2171, n_4708, n_2768, n_2314, n_4826, n_2420, n_3343, n_514, n_1079, n_1593, n_3767, n_442, n_2299, n_131, n_2540, n_2873, n_4589, n_4578, n_1640, n_2162, n_2847, n_1148, n_2051, n_3221, n_742, n_750, n_2168, n_2790, n_3629, n_3021, n_185, n_2359, n_3674, n_3502, n_3098, n_1383, n_5013, n_2312, n_3015, n_1171, n_1920, n_1065, n_4147, n_2048, n_3607, n_4925, n_1921, n_1309, n_4974, n_355, n_1800, n_1548, n_4932, n_1421, n_4510, n_2571, n_1286, n_1177, n_3276, n_3787, n_2124, n_613, n_1119, n_1240, n_3827, n_829, n_2519, n_3354, n_2724, n_4447, n_4285, n_4651, n_361, n_700, n_573, n_4818, n_4514, n_388, n_1366, n_4800, n_3960, n_3248, n_2277, n_1568, n_2110, n_274, n_582, n_1332, n_4433, n_2879, n_73, n_2474, n_19, n_2090, n_3153, n_512, n_1591, n_2033, n_4341, n_1682, n_4312, n_2628, n_3399, n_1249, n_1111, n_25, n_2132, n_2400, n_4633, n_609, n_3838, n_1909, n_4277, n_112, n_4140, n_3675, n_1140, n_891, n_3387, n_4662, n_3779, n_2464, n_2831, n_102, n_1456, n_4882, n_4993, n_2365, n_4832, n_4207, n_987, n_4545, n_3037, n_261, n_4868, n_1885, n_2452, n_3925, n_2176, n_1816, n_4059, n_2455, n_4595, n_1849, n_1131, n_2467, n_1094, n_2288, n_4063, n_346, n_1209, n_3592, n_4650, n_602, n_4888, n_1435, n_879, n_3394, n_4874, n_3793, n_16, n_4669, n_405, n_4339, n_1645, n_4041, n_2858, n_4060, n_996, n_2658, n_1717, n_2895, n_2128, n_3097, n_120, n_327, n_135, n_4541, n_3824, n_3388, n_4494, n_3059, n_3465, n_1316, n_4796, n_1438, n_3589, n_62, n_952, n_2534, n_1229, n_4799, n_3449, n_2694, n_2198, n_2610, n_2989, n_2789, n_4775, n_2216, n_531, n_1897, n_764, n_1424, n_162, n_2933, n_4381, n_4266, n_3886, n_4455, n_2328, n_199, n_4248, n_4754, n_4554, n_4845, n_3053, n_1299, n_3893, n_1141, n_2465, n_3548, n_4585, n_418, n_315, n_451, n_1699, n_3334, n_2541, n_4383, n_1139, n_57, n_397, n_1432, n_3875, n_4003, n_2402, n_4301, n_841, n_1050, n_4586, n_1954, n_4048, n_1844, n_3777, n_4784, n_2999, n_1644, n_4046, n_1974, n_2086, n_3537, n_3080, n_4199, n_2701, n_3362, n_1631, n_3105, n_1179, n_753, n_1048, n_4286, n_2556, n_2269, n_3274, n_3041, n_4470, n_2236, n_330, n_2816, n_692, n_820, n_1911, n_3616, n_2460, n_4058, n_3664, n_4188, n_1668, n_3913, n_3417, n_1143, n_1579, n_4034, n_1688, n_492, n_3327, n_4689, n_341, n_3067, n_2755, n_543, n_3237, n_1992, n_4402, n_4239, n_3400, n_449, n_4550, n_1214, n_1342, n_1400, n_3382, n_3574, n_2169, n_1557, n_4201, n_618, n_896, n_3316, n_356, n_3099, n_3704, n_2596, n_1730, n_3603, n_4123, n_2192, n_964, n_3633, n_4479, n_1373, n_2670, n_5, n_1646, n_1307, n_4416, n_3372, n_4539, n_814, n_2707, n_2471, n_1472, n_1671, n_3230, n_1062, n_3342, n_4682, n_3708, n_1204, n_3729, n_4978, n_4690, n_4437, n_3861, n_4736, n_3780, n_783, n_1928, n_1188, n_3957, n_3848, n_41, n_4284, n_2600, n_3919, n_336, n_3608, n_510, n_216, n_4513, n_3233, n_3829, n_3177, n_4053, n_2352, n_4040, n_2207, n_2619, n_2444, n_241, n_1110, n_3123, n_1088, n_3393, n_638, n_866, n_4887, n_4617, n_3520, n_2492, n_249, n_577, n_4005, n_1687, n_1637, n_4904, n_1419, n_693, n_4792, n_3578, n_3812, n_1886, n_1389, n_1256, n_4980, n_1465, n_4290, n_306, n_1375, n_3727, n_3774, n_3093, n_1843, n_3061, n_1597, n_1659, n_2431, n_1371, n_4956, n_2206, n_3182, n_2564, n_4947, n_876, n_4656, n_1190, n_3896, n_3958, n_3450, n_966, n_4729, n_4987, n_4971, n_1116, n_2000, n_1212, n_2074, n_206, n_3174, n_982, n_1453, n_2217, n_1183, n_3398, n_2307, n_3408, n_899, n_2722, n_2640, n_4823, n_4875, n_1628, n_3432, n_1514, n_1771, n_557, n_1005, n_607, n_679, n_710, n_3090, n_527, n_1168, n_2437, n_3762, n_2445, n_1427, n_108, n_1835, n_66, n_177, n_1988, n_1853, n_1356, n_1787, n_4137, n_2634, n_4529, n_910, n_4323, n_3034, n_2212, n_3972, n_125, n_529, n_126, n_202, n_3308, n_791, n_1533, n_5036, n_4772, n_3467, n_4322, n_1720, n_2830, n_4354, n_159, n_4653, n_2354, n_2246, n_4677, n_3901, n_715, n_1480, n_3757, n_3381, n_1782, n_2245, n_4909, n_1524, n_1485, n_115, n_810, n_2965, n_416, n_3635, n_5022, n_5005, n_1144, n_2814, n_1570, n_3882, n_3046, n_1170, n_305, n_2213, n_3826, n_3211, n_2211, n_2095, n_3121, n_4634, n_3337, n_2527, n_855, n_1461, n_3204, n_2136, n_1273, n_1822, n_4952, n_3005, n_1235, n_4380, n_980, n_698, n_3129, n_4126, n_1282, n_1783, n_2601, n_3043, n_998, n_3802, n_2375, n_4506, n_4880, n_1907, n_501, n_2686, n_2344, n_3892, n_4896, n_1417, n_1295, n_1985, n_2107, n_3219, n_2906, n_4943, n_382, n_2187, n_1762, n_1013, n_718, n_3023, n_4193, n_4075, n_3104, n_612, n_4737, n_3647, n_825, n_2819, n_506, n_737, n_3609, n_4136, n_1715, n_1952, n_4393, n_3720, n_4535, n_733, n_1922, n_2560, n_4522, n_4794, n_3959, n_63, n_792, n_3140, n_3724, n_298, n_2104, n_505, n_3011, n_4196, n_1425, n_4592, n_4675, n_3069, n_4370, n_1900, n_1620, n_3084, n_1727, n_2735, n_2497, n_3412, n_1995, n_2411, n_1046, n_3761, n_4889, n_2014, n_2986, n_1641, n_1361, n_3184, n_4828, n_4558, n_2172, n_4722, n_1129, n_158, n_3626, n_4768, n_4100, n_961, n_2250, n_276, n_1225, n_169, n_400, n_4092, n_3908, n_2423, n_3671, n_994, n_3344, n_2194, n_848, n_4465, n_3302, n_1223, n_2680, n_1567, n_3122, n_4808, n_3842, n_145, n_3265, n_1857, n_4482, n_2041, n_631, n_479, n_1797, n_2957, n_2357, n_1250, n_3309, n_608, n_772, n_3260, n_4926, n_3357, n_1589, n_4116, n_1086, n_2570, n_1858, n_1619, n_2815, n_3754, n_4612, n_1469, n_2744, n_4287, n_2397, n_384, n_2208, n_3063, n_3617, n_333, n_1298, n_1652, n_4516, n_3794, n_2809, n_2050, n_4505, n_1676, n_258, n_1113, n_29, n_1277, n_2591, n_188, n_3384, n_852, n_4602, n_4449, n_1864, n_463, n_502, n_466, n_420, n_1337, n_4445, n_699, n_1627, n_1245, n_4870, n_2438, n_465, n_2832, n_362, n_1321, n_1975, n_2296, n_273, n_3181, n_616, n_2278, n_4915, n_2135, n_3493, n_3323, n_2734, n_4914, n_1076, n_2823, n_1408, n_494, n_1761, n_730, n_354, n_795, n_4345, n_180, n_3281, n_656, n_3307, n_1606, n_1220, n_1694, n_4318, n_2485, n_2655, n_60, n_4185, n_4797, n_2366, n_1526, n_3997, n_1604, n_1275, n_4032, n_1764, n_3582, n_712, n_1583, n_2826, n_3539, n_1042, n_285, n_412, n_4343, n_1493, n_4212, n_4124, n_4492, n_2708, n_4994, n_4245, n_4364, n_4928, n_2225, n_1507, n_4378, n_2383, n_1996, n_597, n_3406, n_3604, n_3853, n_4216, n_2019, n_1340, n_1558, n_2166, n_2938, n_4309, n_3594, n_262, n_1704, n_3721, n_1254, n_1026, n_2026, n_1234, n_2109, n_364, n_2013, n_20, n_1990, n_1032, n_2614, n_2991, n_2242, n_2752, n_2894, n_3473, n_4560, n_2839, n_1588, n_2237, n_3463, n_3699, n_3360, n_2524, n_3873, n_3693, n_2728, n_3857, n_18332);

input n_924;
input n_977;
input n_2253;
input n_2417;
input n_2756;
input n_4706;
input n_2380;
input n_3241;
input n_3006;
input n_532;
input n_2327;
input n_1488;
input n_2899;
input n_790;
input n_3619;
input n_3541;
input n_3622;
input n_2395;
input n_2347;
input n_4963;
input n_4240;
input n_4508;
input n_2021;
input n_2391;
input n_5035;
input n_1960;
input n_2843;
input n_4;
input n_551;
input n_3615;
input n_2059;
input n_1466;
input n_1695;
input n_2487;
input n_3202;
input n_4977;
input n_3813;
input n_671;
input n_3341;
input n_3587;
input n_4128;
input n_3445;
input n_2001;
input n_4145;
input n_3785;
input n_5033;
input n_1462;
input n_4211;
input n_3448;
input n_3019;
input n_2096;
input n_877;
input n_3776;
input n_2530;
input n_4517;
input n_1696;
input n_2483;
input n_4425;
input n_4950;
input n_4988;
input n_1285;
input n_1860;
input n_4615;
input n_87;
input n_1107;
input n_1728;
input n_2076;
input n_668;
input n_301;
input n_2147;
input n_3010;
input n_2770;
input n_4131;
input n_2584;
input n_171;
input n_3188;
input n_3403;
input n_3624;
input n_3461;
input n_3082;
input n_2189;
input n_3796;
input n_1242;
input n_3283;
input n_519;
input n_2323;
input n_2597;
input n_3340;
input n_3277;
input n_281;
input n_2052;
input n_4499;
input n_4927;
input n_731;
input n_1314;
input n_1512;
input n_1490;
input n_317;
input n_569;
input n_3214;
input n_1517;
input n_2091;
input n_4311;
input n_3631;
input n_3806;
input n_4691;
input n_1449;
input n_4678;
input n_1566;
input n_2032;
input n_297;
input n_2587;
input n_156;
input n_219;
input n_157;
input n_3947;
input n_3490;
input n_600;
input n_223;
input n_1948;
input n_3868;
input n_3183;
input n_3437;
input n_3353;
input n_264;
input n_4203;
input n_3687;
input n_882;
input n_2384;
input n_3156;
input n_696;
input n_3376;
input n_646;
input n_5037;
input n_436;
input n_4468;
input n_3653;
input n_3702;
input n_1040;
input n_4976;
input n_2202;
input n_2648;
input n_5008;
input n_2159;
input n_2976;
input n_3876;
input n_2353;
input n_2439;
input n_4811;
input n_2276;
input n_2089;
input n_3420;
input n_72;
input n_1561;
input n_1165;
input n_1034;
input n_3361;
input n_4758;
input n_1600;
input n_521;
input n_845;
input n_528;
input n_4255;
input n_1796;
input n_395;
input n_553;
input n_901;
input n_4484;
input n_3668;
input n_4237;
input n_2934;
input n_1672;
input n_1880;
input n_3550;
input n_1626;
input n_637;
input n_144;
input n_2079;
input n_2238;
input n_96;
input n_1151;
input n_1405;
input n_1706;
input n_3418;
input n_342;
input n_4901;
input n_197;
input n_2859;
input n_1075;
input n_3395;
input n_4917;
input n_2863;
input n_2072;
input n_2738;
input n_2968;
input n_1585;
input n_2684;
input n_3593;
input n_1599;
input n_4421;
input n_4836;
input n_4020;
input n_2730;
input n_2251;
input n_3915;
input n_1377;
input n_4469;
input n_4414;
input n_190;
input n_4532;
input n_3339;
input n_228;
input n_283;
input n_3349;
input n_3735;
input n_2248;
input n_3007;
input n_1000;
input n_2622;
input n_2062;
input n_2668;
input n_1002;
input n_2100;
input n_310;
input n_3310;
input n_54;
input n_3487;
input n_2258;
input n_748;
input n_1058;
input n_1667;
input n_838;
input n_3983;
input n_332;
input n_1053;
input n_1224;
input n_4405;
input n_1926;
input n_1331;
input n_4195;
input n_279;
input n_1014;
input n_4969;
input n_1241;
input n_4504;
input n_1385;
input n_440;
input n_793;
input n_2776;
input n_4408;
input n_2140;
input n_2385;
input n_1819;
input n_4531;
input n_476;
input n_2987;
input n_1527;
input n_4567;
input n_4164;
input n_4234;
input n_345;
input n_4130;
input n_3611;
input n_2862;
input n_2175;
input n_2324;
input n_2606;
input n_3187;
input n_2828;
input n_182;
input n_4471;
input n_5031;
input n_407;
input n_3392;
input n_3975;
input n_3430;
input n_4444;
input n_3208;
input n_207;
input n_3331;
input n_2379;
input n_4983;
input n_2911;
input n_2154;
input n_4916;
input n_3649;
input n_4302;
input n_2514;
input n_4786;
input n_3257;
input n_1027;
input n_326;
input n_4160;
input n_2293;
input n_4051;
input n_2028;
input n_558;
input n_3009;
input n_1276;
input n_1412;
input n_3981;
input n_1199;
input n_352;
input n_1038;
input n_520;
input n_1841;
input n_154;
input n_2581;
input n_71;
input n_3224;
input n_4647;
input n_3752;
input n_870;
input n_1711;
input n_1891;
input n_434;
input n_3526;
input n_2546;
input n_965;
input n_3790;
input n_3491;
input n_935;
input n_817;
input n_1175;
input n_4613;
input n_4649;
input n_64;
input n_1888;
input n_1963;
input n_4795;
input n_2226;
input n_2891;
input n_4028;
input n_103;
input n_97;
input n_7;
input n_1690;
input n_3819;
input n_2449;
input n_431;
input n_1194;
input n_2297;
input n_4186;
input n_4731;
input n_1759;
input n_2177;
input n_3747;
input n_2227;
input n_4618;
input n_127;
input n_2190;
input n_3346;
input n_4742;
input n_2876;
input n_4099;
input n_452;
input n_3484;
input n_3620;
input n_1260;
input n_1746;
input n_2479;
input n_1464;
input n_4295;
input n_649;
input n_1444;
input n_4694;
input n_4533;
input n_3038;
input n_3068;
input n_2871;
input n_4244;
input n_4603;
input n_2943;
input n_4254;
input n_3143;
input n_3168;
input n_1680;
input n_4697;
input n_2607;
input n_3994;
input n_4190;
input n_4810;
input n_3317;
input n_1121;
input n_433;
input n_8;
input n_4391;
input n_949;
input n_3263;
input n_2582;
input n_4157;
input n_4283;
input n_4681;
input n_1001;
input n_1503;
input n_4638;
input n_1468;
input n_3455;
input n_3452;
input n_1510;
input n_1380;
input n_1994;
input n_1195;
input n_4707;
input n_2577;
input n_4527;
input n_2796;
input n_757;
input n_2342;
input n_106;
input n_4156;
input n_1851;
input n_4848;
input n_2937;
input n_3095;
input n_2805;
input n_1145;
input n_524;
input n_394;
input n_4918;
input n_1153;
input n_3856;
input n_741;
input n_2914;
input n_4898;
input n_1964;
input n_2869;
input n_4002;
input n_1163;
input n_1207;
input n_5010;
input n_2406;
input n_3623;
input n_2846;
input n_2925;
input n_3773;
input n_3918;
input n_2398;
input n_2857;
input n_4528;
input n_3932;
input n_4619;
input n_4673;
input n_940;
input n_3516;
input n_4822;
input n_2155;
input n_2516;
input n_3797;
input n_1596;
input n_2947;
input n_123;
input n_978;
input n_4299;
input n_4801;
input n_1474;
input n_1665;
input n_1269;
input n_3515;
input n_2886;
input n_267;
input n_2093;
input n_2473;
input n_1208;
input n_3287;
input n_3378;
input n_1431;
input n_4279;
input n_4769;
input n_4632;
input n_660;
input n_4294;
input n_1732;
input n_4125;
input n_4232;
input n_4949;
input n_374;
input n_2941;
input n_2457;
input n_4790;
input n_459;
input n_962;
input n_723;
input n_2536;
input n_1336;
input n_1758;
input n_2952;
input n_4847;
input n_3058;
input n_4365;
input n_1878;
input n_3505;
input n_4610;
input n_88;
input n_3730;
input n_4489;
input n_168;
input n_974;
input n_727;
input n_4967;
input n_957;
input n_4992;
input n_3001;
input n_303;
input n_3945;
input n_4542;
input n_2261;
input n_2729;
input n_3597;
input n_1612;
input n_2897;
input n_2077;
input n_4198;
input n_2909;
input n_4534;
input n_4500;
input n_5014;
input n_69;
input n_3185;
input n_1300;
input n_1127;
input n_3523;
input n_1785;
input n_2829;
input n_4597;
input n_4329;
input n_1006;
input n_4087;
input n_3811;
input n_1270;
input n_1664;
input n_3200;
input n_2231;
input n_2017;
input n_2604;
input n_4257;
input n_3453;
input n_322;
input n_2390;
input n_3213;
input n_1041;
input n_3077;
input n_1562;
input n_383;
input n_3474;
input n_3984;
input n_239;
input n_630;
input n_2151;
input n_55;
input n_2106;
input n_2716;
input n_4665;
input n_1913;
input n_1823;
input n_3679;
input n_3422;
input n_3888;
input n_4189;
input n_1875;
input n_1304;
input n_2803;
input n_1324;
input n_3707;
input n_1846;
input n_3429;
input n_1903;
input n_3849;
input n_3946;
input n_860;
input n_3229;
input n_4463;
input n_1805;
input n_429;
input n_4687;
input n_948;
input n_4670;
input n_4084;
input n_4703;
input n_4037;
input n_2922;
input n_83;
input n_3275;
input n_3499;
input n_2645;
input n_2727;
input n_560;
input n_340;
input n_3421;
input n_2240;
input n_2436;
input n_1552;
input n_3618;
input n_574;
input n_2593;
input n_3683;
input n_58;
input n_3642;
input n_3286;
input n_3808;
input n_824;
input n_359;
input n_1327;
input n_4763;
input n_1684;
input n_3590;
input n_366;
input n_815;
input n_4594;
input n_3424;
input n_1381;
input n_1037;
input n_2301;
input n_3583;
input n_3560;
input n_4076;
input n_4714;
input n_2419;
input n_3215;
input n_589;
input n_4776;
input n_2122;
input n_2512;
input n_4102;
input n_2786;
input n_3171;
input n_1437;
input n_645;
input n_238;
input n_3020;
input n_3677;
input n_3462;
input n_3468;
input n_1893;
input n_2910;
input n_222;
input n_1123;
input n_1467;
input n_2163;
input n_634;
input n_32;
input n_2254;
input n_1382;
input n_925;
input n_3546;
input n_424;
input n_2647;
input n_1311;
input n_1519;
input n_256;
input n_950;
input n_4443;
input n_4507;
input n_1811;
input n_2443;
input n_2624;
input n_3012;
input n_4575;
input n_380;
input n_419;
input n_3244;
input n_389;
input n_3130;
input n_3822;
input n_3569;
input n_912;
input n_136;
input n_86;
input n_968;
input n_4452;
input n_4348;
input n_619;
input n_376;
input n_4355;
input n_3494;
input n_515;
input n_351;
input n_885;
input n_2125;
input n_3771;
input n_683;
input n_3110;
input n_1057;
input n_1051;
input n_721;
input n_1157;
input n_3073;
input n_4572;
input n_22;
input n_802;
input n_4026;
input n_2265;
input n_4104;
input n_1608;
input n_4512;
input n_3554;
input n_38;
input n_4377;
input n_280;
input n_1305;
input n_3178;
input n_873;
input n_2334;
input n_690;
input n_33;
input n_4521;
input n_583;
input n_4488;
input n_2289;
input n_3051;
input n_302;
input n_1343;
input n_2783;
input n_2263;
input n_3750;
input n_2341;
input n_3632;
input n_4588;
input n_2733;
input n_1288;
input n_212;
input n_2785;
input n_2415;
input n_3299;
input n_4519;
input n_3715;
input n_972;
input n_3040;
input n_1938;
input n_1200;
input n_2499;
input n_3568;
input n_3737;
input n_1185;
input n_991;
input n_1967;
input n_576;
input n_1329;
input n_3255;
input n_4856;
input n_2997;
input n_4400;
input n_943;
input n_3326;
input n_3734;
input n_650;
input n_4778;
input n_286;
input n_2429;
input n_883;
input n_470;
input n_325;
input n_132;
input n_856;
input n_1793;
input n_4352;
input n_4441;
input n_918;
input n_4761;
input n_942;
input n_1804;
input n_189;
input n_4347;
input n_4095;
input n_3196;
input n_4593;
input n_2364;
input n_2533;
input n_3492;
input n_2780;
input n_4727;
input n_4568;
input n_195;
input n_2291;
input n_4043;
input n_1636;
input n_3601;
input n_1350;
input n_1865;
input n_2973;
input n_1096;
input n_2094;
input n_1575;
input n_2393;
input n_1697;
input n_3831;
input n_3801;
input n_225;
input n_2043;
input n_2751;
input n_192;
input n_4893;
input n_5032;
input n_1549;
input n_1934;
input n_4948;
input n_4000;
input n_655;
input n_3240;
input n_2025;
input n_1446;
input n_4406;
input n_2758;
input n_1458;
input n_472;
input n_1807;
input n_387;
input n_2618;
input n_398;
input n_2559;
input n_763;
input n_4748;
input n_2295;
input n_3931;
input n_1219;
input n_4010;
input n_2840;
input n_5017;
input n_1814;
input n_2822;
input n_4710;
input n_287;
input n_555;
input n_4607;
input n_4117;
input n_3636;
input n_1722;
input n_2441;
input n_1802;
input n_3083;
input n_4487;
input n_5001;
input n_2795;
input n_2981;
input n_2282;
input n_2800;
input n_4817;
input n_311;
input n_3380;
input n_2098;
input n_1296;
input n_3460;
input n_3409;
input n_3538;
input n_2068;
input n_4849;
input n_4867;
input n_445;
input n_2641;
input n_3198;
input n_1895;
input n_4728;
input n_588;
input n_789;
input n_4247;
input n_4933;
input n_107;
input n_4018;
input n_3900;
input n_1105;
input n_4902;
input n_4518;
input n_4409;
input n_4411;
input n_3872;
input n_4336;
input n_149;
input n_2270;
input n_4777;
input n_2653;
input n_836;
input n_2496;
input n_1908;
input n_2259;
input n_3877;
input n_458;
input n_2995;
input n_2494;
input n_3547;
input n_3977;
input n_1102;
input n_4052;
input n_3459;
input n_1499;
input n_4398;
input n_3155;
input n_2633;
input n_4954;
input n_2435;
input n_1392;
input n_1164;
input n_2097;
input n_4304;
input n_3911;
input n_1303;
input n_4431;
input n_4192;
input n_3736;
input n_4805;
input n_118;
input n_601;
input n_4885;
input n_253;
input n_1661;
input n_3565;
input n_172;
input n_4701;
input n_2575;
input n_861;
input n_1658;
input n_1904;
input n_1345;
input n_176;
input n_1899;
input n_1003;
input n_2067;
input n_2219;
input n_3533;
input n_2877;
input n_2148;
input n_393;
input n_4631;
input n_1726;
input n_3035;
input n_421;
input n_1657;
input n_768;
input n_1475;
input n_1725;
input n_1313;
input n_1136;
input n_1491;
input n_754;
input n_3639;
input n_708;
input n_735;
input n_2501;
input n_3079;
input n_4965;
input n_1915;
input n_1109;
input n_1310;
input n_2605;
input n_4747;
input n_1399;
input n_1979;
input n_193;
input n_2924;
input n_4111;
input n_808;
input n_2484;
input n_797;
input n_1025;
input n_4587;
input n_3731;
input n_2946;
input n_4538;
input n_435;
input n_766;
input n_541;
input n_1117;
input n_2754;
input n_687;
input n_1742;
input n_2489;
input n_536;
input n_2012;
input n_1291;
input n_4094;
input n_3503;
input n_2866;
input n_3561;
input n_1155;
input n_1418;
input n_1011;
input n_2917;
input n_2425;
input n_3536;
input n_3661;
input n_4150;
input n_827;
input n_4878;
input n_1703;
input n_1650;
input n_1137;
input n_3934;
input n_4985;
input n_3922;
input n_3846;
input n_318;
input n_2103;
input n_653;
input n_2160;
input n_2498;
input n_2697;
input n_850;
input n_3074;
input n_1999;
input n_2372;
input n_3673;
input n_3768;
input n_1372;
input n_2861;
input n_605;
input n_2630;
input n_3943;
input n_353;
input n_2430;
input n_493;
input n_2433;
input n_3293;
input n_4022;
input n_1531;
input n_840;
input n_1334;
input n_4852;
input n_2528;
input n_4869;
input n_4700;
input n_4035;
input n_2316;
input n_1898;
input n_3294;
input n_4426;
input n_554;
input n_3415;
input n_2284;
input n_2817;
input n_3139;
input n_2598;
input n_4601;
input n_2687;
input n_1120;
input n_198;
input n_1890;
input n_714;
input n_4220;
input n_1944;
input n_909;
input n_1497;
input n_3431;
input n_3169;
input n_3151;
input n_2078;
input n_3284;
input n_3070;
input n_4066;
input n_119;
input n_2884;
input n_4515;
input n_4351;
input n_3126;
input n_4403;
input n_1981;
input n_1663;
input n_1718;
input n_4509;
input n_4858;
input n_3700;
input n_509;
input n_147;
input n_1518;
input n_4223;
input n_1281;
input n_1889;
input n_209;
input n_1489;
input n_5025;
input n_2966;
input n_1376;
input n_2326;
input n_1569;
input n_2188;
input n_186;
input n_756;
input n_1429;
input n_4644;
input n_4456;
input n_399;
input n_2448;
input n_4346;
input n_3170;
input n_2748;
input n_3311;
input n_3272;
input n_2898;
input n_2717;
input n_1861;
input n_760;
input n_3628;
input n_3691;
input n_220;
input n_4235;
input n_1867;
input n_1945;
input n_3018;
input n_481;
input n_2573;
input n_4435;
input n_2939;
input n_3807;
input n_271;
input n_2447;
input n_4764;
input n_886;
input n_1221;
input n_167;
input n_2774;
input n_1707;
input n_853;
input n_4655;
input n_3161;
input n_377;
input n_4581;
input n_751;
input n_4827;
input n_2488;
input n_392;
input n_3477;
input n_2476;
input n_704;
input n_4399;
input n_2781;
input n_2778;
input n_771;
input n_4782;
input n_1520;
input n_4363;
input n_2887;
input n_1287;
input n_4864;
input n_1262;
input n_2691;
input n_1411;
input n_3054;
input n_4335;
input n_2526;
input n_2703;
input n_2167;
input n_3391;
input n_4259;
input n_56;
input n_2709;
input n_816;
input n_1536;
input n_4865;
input n_4056;
input n_1344;
input n_4564;
input n_1246;
input n_3840;
input n_1339;
input n_3518;
input n_2956;
input n_3733;
input n_328;
input n_2173;
input n_1842;
input n_871;
input n_3738;
input n_685;
input n_78;
input n_3464;
input n_2018;
input n_4526;
input n_1555;
input n_3245;
input n_4417;
input n_499;
input n_98;
input n_402;
input n_4899;
input n_796;
input n_2119;
input n_1502;
input n_2157;
input n_2552;
input n_1012;
input n_1;
input n_2453;
input n_4798;
input n_1525;
input n_740;
input n_3509;
input n_3352;
input n_3076;
input n_3535;
input n_2182;
input n_277;
input n_1061;
input n_3251;
input n_92;
input n_2931;
input n_1193;
input n_3118;
input n_3511;
input n_1226;
input n_3443;
input n_2146;
input n_1487;
input n_3644;
input n_3336;
input n_3935;
input n_781;
input n_542;
input n_3521;
input n_3562;
input n_3948;
input n_4750;
input n_1515;
input n_2918;
input n_3232;
input n_1673;
input n_27;
input n_2112;
input n_1739;
input n_2958;
input n_3114;
input n_3125;
input n_4981;
input n_2394;
input n_3612;
input n_2954;
input n_4835;
input n_4430;
input n_4081;
input n_1103;
input n_3132;
input n_4407;
input n_648;
input n_312;
input n_3951;
input n_4894;
input n_3238;
input n_3210;
input n_2036;
input n_3267;
input n_4995;
input n_480;
input n_425;
input n_695;
input n_37;
input n_3964;
input n_3772;
input n_229;
input n_1956;
input n_437;
input n_1642;
input n_2279;
input n_3373;
input n_4446;
input n_3884;
input n_0;
input n_3726;
input n_805;
input n_2525;
input n_2892;
input n_113;
input n_2907;
input n_3577;
input n_2820;
input n_269;
input n_2049;
input n_2273;
input n_2719;
input n_1741;
input n_1160;
input n_4057;
input n_4332;
input n_1258;
input n_4314;
input n_1074;
input n_3347;
input n_3216;
input n_1621;
input n_3809;
input n_2113;
input n_1448;
input n_4288;
input n_3567;
input n_1634;
input n_3939;
input n_4241;
input n_3321;
input n_3212;
input n_666;
input n_1433;
input n_2256;
input n_3152;
input n_319;
input n_2920;
input n_4265;
input n_1186;
input n_1018;
input n_2247;
input n_713;
input n_1622;
input n_166;
input n_1180;
input n_3705;
input n_2802;
input n_4705;
input n_3159;
input n_2268;
input n_3778;
input n_3304;
input n_1378;
input n_3912;
input n_1729;
input n_2739;
input n_469;
input n_2771;
input n_4604;
input n_549;
input n_3795;
input n_5020;
input n_4419;
input n_4477;
input n_3179;
input n_3256;
input n_667;
input n_2386;
input n_1501;
input n_3086;
input n_1007;
input n_2369;
input n_2927;
input n_4217;
input n_4395;
input n_2821;
input n_1099;
input n_2568;
input n_564;
input n_1738;
input n_3728;
input n_21;
input n_3064;
input n_3088;
input n_1021;
input n_4639;
input n_3713;
input n_3663;
input n_3246;
input n_2495;
input n_1535;
input n_1789;
input n_819;
input n_2302;
input n_951;
input n_247;
input n_1494;
input n_292;
input n_625;
input n_2069;
input n_417;
input n_3434;
input n_1806;
input n_933;
input n_1563;
input n_4227;
input n_26;
input n_4033;
input n_4289;
input n_2024;
input n_4780;
input n_755;
input n_4243;
input n_4982;
input n_530;
input n_4330;
input n_3695;
input n_556;
input n_2482;
input n_2677;
input n_3832;
input n_3987;
input n_902;
input n_4991;
input n_579;
input n_1698;
input n_2329;
input n_1098;
input n_2142;
input n_320;
input n_3332;
input n_1135;
input n_3048;
input n_3937;
input n_2203;
input n_4525;
input n_1243;
input n_101;
input n_3782;
input n_2978;
input n_2058;
input n_2458;
input n_4208;
input n_3786;
input n_371;
input n_2888;
input n_3638;
input n_1236;
input n_1633;
input n_4177;
input n_3763;
input n_2669;
input n_1778;
input n_2306;
input n_3022;
input n_4264;
input n_335;
input n_3087;
input n_3489;
input n_2566;
input n_343;
input n_308;
input n_2149;
input n_1078;
input n_3060;
input n_4276;
input n_3013;
input n_1984;
input n_2408;
input n_1877;
input n_3049;
input n_1723;
input n_339;
input n_4485;
input n_183;
input n_4626;
input n_1036;
input n_1097;
input n_347;
input n_798;
input n_2659;
input n_1414;
input n_290;
input n_4975;
input n_1852;
input n_578;
input n_344;
input n_3089;
input n_422;
input n_2470;
input n_3985;
input n_496;
input n_1391;
input n_670;
input n_4760;
input n_4652;
input n_4624;
input n_48;
input n_663;
input n_2551;
input n_1587;
input n_2682;
input n_813;
input n_1284;
input n_3440;
input n_1748;
input n_4569;
input n_2699;
input n_4897;
input n_888;
input n_2769;
input n_3542;
input n_3436;
input n_2615;
input n_3940;
input n_446;
input n_1064;
input n_858;
input n_2985;
input n_691;
input n_2753;
input n_363;
input n_1582;
input n_3637;
input n_2842;
input n_4523;
input n_1836;
input n_2868;
input n_3141;
input n_3164;
input n_3570;
input n_4919;
input n_4025;
input n_461;
input n_2712;
input n_3936;
input n_4503;
input n_3507;
input n_3821;
input n_2700;
input n_1211;
input n_3367;
input n_4464;
input n_907;
input n_3096;
input n_3496;
input n_4114;
input n_989;
input n_2544;
input n_2356;
input n_488;
input n_892;
input n_4556;
input n_2620;
input n_1581;
input n_4089;
input n_586;
input n_2919;
input n_4327;
input n_230;
input n_953;
input n_4218;
input n_2150;
input n_3146;
input n_2241;
input n_2757;
input n_963;
input n_1052;
input n_954;
input n_478;
input n_4353;
input n_2042;
input n_534;
input n_884;
input n_1754;
input n_1623;
input n_2921;
input n_2720;
input n_1854;
input n_4990;
input n_1856;
input n_143;
input n_4959;
input n_4161;
input n_237;
input n_832;
input n_1319;
input n_3992;
input n_2616;
input n_1906;
input n_4103;
input n_1387;
input n_4466;
input n_2262;
input n_2462;
input n_1532;
input n_18;
input n_3625;
input n_1156;
input n_794;
input n_2798;
input n_2945;
input n_2331;
input n_686;
input n_2837;
input n_847;
input n_4844;
input n_2979;
input n_3655;
input n_4688;
input n_4765;
input n_702;
input n_2548;
input n_822;
input n_2108;
input n_3640;
input n_4388;
input n_4206;
input n_1538;
input n_1779;
input n_4738;
input n_53;
input n_1369;
input n_3909;
input n_3207;
input n_3944;
input n_809;
input n_4434;
input n_4837;
input n_3042;
input n_1942;
input n_2510;
input n_4219;
input n_2804;
input n_3659;
input n_2120;
input n_411;
input n_414;
input n_5012;
input n_1293;
input n_1876;
input n_4620;
input n_36;
input n_1810;
input n_2813;
input n_4438;
input n_2009;
input n_2222;
input n_3510;
input n_28;
input n_3218;
input n_2667;
input n_11;
input n_3150;
input n_747;
input n_52;
input n_4325;
input n_1733;
input n_2413;
input n_615;
input n_851;
input n_843;
input n_705;
input n_3775;
input n_4133;
input n_678;
input n_4184;
input n_2518;
input n_2629;
input n_367;
input n_4481;
input n_3416;
input n_4379;
input n_2181;
input n_1829;
input n_547;
input n_4030;
input n_116;
input n_4490;
input n_3138;
input n_4397;
input n_1710;
input n_1128;
input n_2928;
input n_1734;
input n_4820;
input n_590;
input n_3770;
input n_1308;
input n_4938;
input n_4179;
input n_3469;
input n_372;
input n_677;
input n_2723;
input n_314;
input n_368;
input n_3220;
input n_4641;
input n_2539;
input n_100;
input n_3855;
input n_1008;
input n_2054;
input n_1559;
input n_4931;
input n_1765;
input n_3158;
input n_1744;
input n_2623;
input n_1617;
input n_295;
input n_133;
input n_3113;
input n_2718;
input n_3760;
input n_4078;
input n_1760;
input n_568;
input n_39;
input n_2856;
input n_1832;
input n_4146;
input n_4360;
input n_3666;
input n_3828;
input n_93;
input n_3288;
input n_4404;
input n_1509;
input n_1874;
input n_4787;
input n_2060;
input n_2613;
input n_1987;
input n_3667;
input n_878;
input n_1306;
input n_3703;
input n_4903;
input n_3558;
input n_2545;
input n_2787;
input n_906;
input n_919;
input n_4356;
input n_658;
input n_2061;
input n_4432;
input n_2378;
input n_1740;
input n_1586;
input n_4291;
input n_535;
input n_4386;
input n_9;
input n_4149;
input n_1492;
input n_592;
input n_1692;
input n_2982;
input n_2481;
input n_3545;
input n_2507;
input n_4019;
input n_2900;
input n_1095;
input n_1614;
input n_2339;
input n_457;
input n_4637;
input n_603;
input n_4935;
input n_4785;
input n_3426;
input n_3454;
input n_3820;
input n_3741;
input n_3410;
input n_2029;
input n_995;
input n_1609;
input n_396;
input n_1887;
input n_4413;
input n_1073;
input n_2346;
input n_662;
input n_3990;
input n_4493;
input n_218;
input n_3475;
input n_1215;
input n_1592;
input n_2882;
input n_1721;
input n_2338;
input n_3672;
input n_3197;
input n_3109;
input n_2721;
input n_1043;
input n_486;
input n_3002;
input n_337;
input n_3897;
input n_1159;
input n_3845;
input n_2081;
input n_299;
input n_4570;
input n_2156;
input n_4296;
input n_1820;
input n_5019;
input n_2418;
input n_2179;
input n_1416;
input n_1724;
input n_2521;
input n_3458;
input n_1420;
input n_1132;
input n_3330;
input n_4606;
input n_4774;
input n_2477;
input n_3887;
input n_4093;
input n_1486;
input n_4672;
input n_3519;
input n_4174;
input n_3374;
input n_3045;
input n_1870;
input n_309;
input n_2367;
input n_4766;
input n_84;
input n_2896;
input n_652;
input n_1365;
input n_4074;
input n_4600;
input n_1927;
input n_1349;
input n_4460;
input n_288;
input n_1031;
input n_3645;
input n_3223;
input n_3929;
input n_834;
input n_2255;
input n_2272;
input n_893;
input n_1965;
input n_1902;
input n_1941;
input n_3938;
input n_2878;
input n_504;
input n_874;
input n_3498;
input n_2015;
input n_1982;
input n_4110;
input n_3189;
input n_2066;
input n_993;
input n_3154;
input n_1551;
input n_545;
input n_450;
input n_2905;
input n_3965;
input n_3566;
input n_1217;
input n_2220;
input n_4349;
input n_628;
input n_3788;
input n_2410;
input n_4313;
input n_1084;
input n_970;
input n_1935;
input n_3366;
input n_1534;
input n_1351;
input n_2696;
input n_4863;
input n_1205;
input n_3242;
input n_495;
input n_3525;
input n_3486;
input n_2405;
input n_3995;
input n_2088;
input n_2953;
input n_4036;
input n_921;
input n_1795;
input n_2578;
input n_3483;
input n_128;
input n_1821;
input n_3894;
input n_3478;
input n_4015;
input n_3890;
input n_2740;
input n_2656;
input n_1080;
input n_1274;
input n_3524;
input n_5034;
input n_1708;
input n_426;
input n_562;
input n_1436;
input n_3549;
input n_1691;
input n_2092;
input n_2075;
input n_3658;
input n_1776;
input n_4807;
input n_2281;
input n_2131;
input n_3026;
input n_1757;
input n_890;
input n_1919;
input n_960;
input n_4230;
input n_3419;
input n_1290;
input n_1047;
input n_2053;
input n_1958;
input n_1252;
input n_348;
input n_3784;
input n_2969;
input n_3941;
input n_2864;
input n_3195;
input n_3190;
input n_1553;
input n_3678;
input n_2664;
input n_3456;
input n_444;
input n_1808;
input n_316;
input n_2266;
input n_2650;
input n_4428;
input n_146;
input n_5003;
input n_408;
input n_967;
input n_2731;
input n_3953;
input n_3166;
input n_4122;
input n_3976;
input n_1357;
input n_3979;
input n_4582;
input n_2998;
input n_4684;
input n_4840;
input n_3162;
input n_983;
input n_2760;
input n_3377;
input n_3749;
input n_3962;
input n_1826;
input n_2304;
input n_762;
input n_1283;
input n_17;
input n_2637;
input n_4384;
input n_4423;
input n_4096;
input n_2881;
input n_1203;
input n_3282;
input n_821;
input n_1763;
input n_3231;
input n_1966;
input n_321;
input n_4996;
input n_621;
input n_2475;
input n_4598;
input n_4478;
input n_507;
input n_2646;
input n_1605;
input n_1228;
input n_3920;
input n_4890;
input n_5027;
input n_3203;
input n_3866;
input n_2903;
input n_3921;
input n_828;
input n_779;
input n_4106;
input n_3717;
input n_2743;
input n_2675;
input n_1439;
input n_3052;
input n_945;
input n_3743;
input n_1932;
input n_4721;
input n_984;
input n_694;
input n_1983;
input n_4029;
input n_1594;
input n_900;
input n_3870;
input n_4496;
input n_3529;
input n_1147;
input n_1977;
input n_2153;
input n_13;
input n_4338;
input n_3094;
input n_2310;
input n_3952;
input n_2287;
input n_2860;
input n_2056;
input n_1470;
input n_1735;
input n_2318;
input n_833;
input n_2502;
input n_2504;
input n_4495;
input n_4762;
input n_2974;
input n_2901;
input n_1940;
input n_2793;
input n_3442;
input n_1201;
input n_1114;
input n_3998;
input n_2285;
input n_3147;
input n_4141;
input n_669;
input n_1176;
input n_1149;
input n_1020;
input n_211;
input n_1824;
input n_1917;
input n_3386;
input n_4107;
input n_3;
input n_4667;
input n_2325;
input n_178;
input n_2446;
input n_3488;
input n_1035;
input n_4547;
input n_2893;
input n_2588;
input n_2962;
input n_4004;
input n_661;
input n_4668;
input n_4953;
input n_3898;
input n_849;
input n_584;
input n_1786;
input n_50;
input n_430;
input n_4997;
input n_4274;
input n_2627;
input n_4759;
input n_1413;
input n_801;
input n_4467;
input n_2080;
input n_2377;
input n_2340;
input n_3552;
input n_875;
input n_357;
input n_3684;
input n_4735;
input n_3137;
input n_165;
input n_2361;
input n_1173;
input n_1603;
input n_969;
input n_1401;
input n_4113;
input n_1019;
input n_1998;
input n_4686;
input n_304;
input n_3759;
input n_4321;
input n_4342;
input n_2034;
input n_3933;
input n_3206;
input n_3966;
input n_1702;
input n_4183;
input n_778;
input n_1122;
input n_4068;
input n_4872;
input n_4233;
input n_3192;
input n_3764;
input n_4709;
input n_5038;
input n_2649;
input n_1187;
input n_1929;
input n_2807;
input n_2542;
input n_2313;
input n_489;
input n_1174;
input n_3324;
input n_3914;
input n_4625;
input n_2558;
input n_2063;
input n_3803;
input n_3742;
input n_2252;
input n_4819;
input n_1685;
input n_917;
input n_1714;
input n_1541;
input n_2576;
input n_4900;
input n_3390;
input n_1573;
input n_3746;
input n_2373;
input n_1713;
input n_3817;
input n_2745;
input n_1253;
input n_210;
input n_1737;
input n_774;
input n_2493;
input n_4930;
input n_1059;
input n_1133;
input n_4537;
input n_2885;
input n_5011;
input n_3318;
input n_4070;
input n_4282;
input n_3485;
input n_4180;
input n_665;
input n_3839;
input n_1440;
input n_3333;
input n_2845;
input n_4143;
input n_4659;
input n_2602;
input n_205;
input n_4579;
input n_4616;
input n_1496;
input n_1125;
input n_3014;
input n_2547;
input n_5023;
input n_1812;
input n_4105;
input n_232;
input n_2532;
input n_3791;
input n_2665;
input n_3905;
input n_427;
input n_3368;
input n_3530;
input n_1930;
input n_1955;
input n_2765;
input n_3329;
input n_2994;
input n_2401;
input n_3135;
input n_2003;
input n_1457;
input n_4895;
input n_3573;
input n_3148;
input n_2264;
input n_3534;
input n_1482;
input n_4275;
input n_1266;
input n_3970;
input n_3438;
input n_4098;
input n_872;
input n_594;
input n_200;
input n_1297;
input n_4789;
input n_1972;
input n_2806;
input n_1184;
input n_2184;
input n_985;
input n_3217;
input n_3404;
input n_3425;
input n_4055;
input n_2926;
input n_626;
input n_3540;
input n_3670;
input n_3973;
input n_2023;
input n_3249;
input n_2351;
input n_676;
input n_4442;
input n_4698;
input n_642;
input n_1602;
input n_194;
input n_1178;
input n_4779;
input n_2286;
input n_4966;
input n_503;
input n_2065;
input n_4017;
input n_3397;
input n_3740;
input n_620;
input n_1081;
input n_4418;
input n_2549;
input n_2705;
input n_2332;
input n_703;
input n_1318;
input n_780;
input n_2977;
input n_1454;
input n_3723;
input n_1227;
input n_3600;
input n_245;
input n_4134;
input n_1388;
input n_2836;
input n_672;
input n_581;
input n_1625;
input n_2130;
input n_898;
input n_3239;
input n_2773;
input n_3365;
input n_3476;
input n_3686;
input n_4913;
input n_1452;
input n_265;
input n_443;
input n_1791;
input n_2850;
input n_1747;
input n_4251;
input n_1817;
input n_3982;
input n_2654;
input n_4621;
input n_1326;
input n_3176;
input n_4559;
input n_2186;
input n_4368;
input n_4740;
input n_5007;
input n_3581;
input n_2562;
input n_4077;
input n_67;
input n_4642;
input n_1192;
input n_2221;
input n_1024;
input n_3576;
input n_1792;
input n_1564;
input n_1868;
input n_1613;
input n_4049;
input n_941;
input n_3862;
input n_68;
input n_3495;
input n_3879;
input n_2348;
input n_4724;
input n_1238;
input n_1772;
input n_282;
input n_752;
input n_1476;
input n_1108;
input n_2818;
input n_1100;
input n_3646;
input n_2129;
input n_3345;
input n_1395;
input n_4546;
input n_862;
input n_3584;
input n_3756;
input n_381;
input n_2889;
input n_390;
input n_5021;
input n_2772;
input n_1675;
input n_1924;
input n_4382;
input n_1554;
input n_3999;
input n_42;
input n_2844;
input n_2138;
input n_2260;
input n_1813;
input n_4833;
input n_3056;
input n_2345;
input n_1172;
input n_379;
input n_428;
input n_1341;
input n_3295;
input n_2382;
input n_4719;
input n_4178;
input n_3062;
input n_2317;
input n_3289;
input n_1973;
input n_786;
input n_1142;
input n_2579;
input n_1770;
input n_138;
input n_4228;
input n_4401;
input n_1756;
input n_1716;
input n_2788;
input n_2984;
input n_3364;
input n_1873;
input n_3201;
input n_221;
input n_622;
input n_1087;
input n_3472;
input n_2874;
input n_4605;
input n_4877;
input n_3235;
input n_4968;
input n_1272;
input n_104;
input n_5030;
input n_3949;
input n_3543;
input n_1247;
input n_591;
input n_3050;
input n_313;
input n_1478;
input n_3903;
input n_4834;
input n_1210;
input n_1364;
input n_2183;
input n_2742;
input n_3314;
input n_4158;
input n_2360;
input n_3254;
input n_369;
input n_4171;
input n_4045;
input n_598;
input n_1367;
input n_4562;
input n_3634;
input n_1460;
input n_2834;
input n_2531;
input n_517;
input n_413;
input n_5015;
input n_2702;
input n_2030;
input n_903;
input n_3115;
input n_4749;
input n_203;
input n_4390;
input n_4979;
input n_1404;
input n_1794;
input n_2234;
input n_4804;
input n_2209;
input n_4270;
input n_2797;
input n_1255;
input n_79;
input n_2321;
input n_722;
input n_3680;
input n_844;
input n_201;
input n_3497;
input n_40;
input n_1601;
input n_2940;
input n_2612;
input n_1495;
input n_4566;
input n_979;
input n_2841;
input n_3322;
input n_4576;
input n_846;
input n_2427;
input n_2505;
input n_76;
input n_4061;
input n_2070;
input n_3250;
input n_585;
input n_270;
input n_2594;
input n_1914;
input n_2335;
input n_2904;
input n_4767;
input n_4328;
input n_3004;
input n_3112;
input n_2349;
input n_1379;
input n_3874;
input n_4676;
input n_4544;
input n_2170;
input n_1091;
input n_641;
input n_3175;
input n_3522;
input n_4429;
input n_575;
input n_4591;
input n_3266;
input n_4646;
input n_1130;
input n_4563;
input n_4725;
input n_2210;
input n_4169;
input n_3247;
input n_3091;
input n_3066;
input n_246;
input n_2426;
input n_657;
input n_4320;
input n_4881;
input n_491;
input n_160;
input n_566;
input n_565;
input n_3613;
input n_3444;
input n_1181;
input n_1505;
input n_4012;
input n_651;
input n_4636;
input n_4584;
input n_807;
input n_3910;
input n_4711;
input n_835;
input n_3319;
input n_3335;
input n_99;
input n_3413;
input n_1969;
input n_4680;
input n_2044;
input n_1138;
input n_927;
input n_2689;
input n_3259;
input n_4191;
input n_4293;
input n_2010;
input n_3688;
input n_3016;
input n_1693;
input n_2599;
input n_904;
input n_3338;
input n_3414;
input n_1827;
input n_4671;
input n_4209;
input n_1271;
input n_1542;
input n_1423;
input n_1166;
input n_1751;
input n_1508;
input n_82;
input n_785;
input n_2200;
input n_3261;
input n_5026;
input n_1161;
input n_3863;
input n_3027;
input n_2746;
input n_1150;
input n_3127;
input n_226;
input n_1780;
input n_3732;
input n_4250;
input n_1055;
input n_3596;
input n_4699;
input n_111;
input n_3906;
input n_4127;
input n_880;
input n_3297;
input n_544;
input n_155;
input n_2683;
input n_1370;
input n_1360;
input n_2388;
input n_4292;
input n_3641;
input n_4577;
input n_4854;
input n_105;
input n_4202;
input n_5000;
input n_2853;
input n_1323;
input n_688;
input n_3766;
input n_1353;
input n_800;
input n_2880;
input n_1666;
input n_3350;
input n_2389;
input n_4165;
input n_4866;
input n_4038;
input n_4109;
input n_915;
input n_864;
input n_1264;
input n_447;
input n_4412;
input n_3407;
input n_3599;
input n_3621;
input n_1580;
input n_2244;
input n_3815;
input n_2257;
input n_497;
input n_1607;
input n_2538;
input n_2105;
input n_2;
input n_3163;
input n_1118;
input n_1686;
input n_947;
input n_373;
input n_3710;
input n_307;
input n_4155;
input n_1359;
input n_2031;
input n_3891;
input n_1230;
input n_4144;
input n_375;
input n_2165;
input n_929;
input n_3379;
input n_4374;
input n_3532;
input n_1124;
input n_1818;
input n_2127;
input n_1576;
input n_1104;
input n_1294;
input n_51;
input n_1257;
input n_1182;
input n_3531;
input n_2963;
input n_3834;
input n_4548;
input n_3258;
input n_24;
input n_4989;
input n_4622;
input n_1016;
input n_4315;
input n_2959;
input n_2047;
input n_1845;
input n_240;
input n_2193;
input n_2478;
input n_4816;
input n_231;
input n_1483;
input n_2983;
input n_227;
input n_3810;
input n_1289;
input n_94;
input n_2715;
input n_2085;
input n_1669;
input n_370;
input n_4483;
input n_2782;
input n_1670;
input n_2672;
input n_2651;
input n_4358;
input n_3656;
input n_2071;
input n_2561;
input n_2643;
input n_1374;
input n_4793;
input n_4168;
input n_3446;
input n_955;
input n_3028;
input n_4806;
input n_1146;
input n_4350;
input n_550;
input n_897;
input n_1428;
input n_1216;
input n_3836;
input n_3963;
input n_1872;
input n_3389;
input n_1931;
input n_4187;
input n_1070;
input n_4166;
input n_1030;
input n_3222;
input n_1071;
input n_1267;
input n_1801;
input n_1513;
input n_2970;
input n_2235;
input n_673;
input n_837;
input n_4937;
input n_3980;
input n_2791;
input n_680;
input n_1473;
input n_3755;
input n_4258;
input n_4498;
input n_1590;
input n_2174;
input n_2714;
input n_3563;
input n_2506;
input n_675;
input n_4064;
input n_4936;
input n_1556;
input n_184;
input n_1863;
input n_3841;
input n_114;
input n_2118;
input n_4770;
input n_2944;
input n_881;
input n_2407;
input n_4907;
input n_468;
input n_129;
input n_3262;
input n_1450;
input n_5018;
input n_4006;
input n_4861;
input n_1322;
input n_3690;
input n_889;
input n_2358;
input n_973;
input n_3716;
input n_1700;
input n_2833;
input n_4712;
input n_477;
input n_3191;
input n_3837;
input n_3193;
input n_1971;
input n_3252;
input n_2275;
input n_2855;
input n_3273;
input n_3544;
input n_4310;
input n_1523;
input n_1950;
input n_1447;
input n_2370;
input n_3954;
input n_3025;
input n_4674;
input n_4908;
input n_736;
input n_2750;
input n_3899;
input n_1278;
input n_4159;
input n_3714;
input n_49;
input n_3071;
input n_3739;
input n_593;
input n_4069;
input n_12;
input n_2784;
input n_3718;
input n_3092;
input n_3470;
input n_4862;
input n_2557;
input n_1248;
input n_70;
input n_289;
input n_4850;
input n_3781;
input n_4813;
input n_4912;
input n_2590;
input n_2330;
input n_2942;
input n_3106;
input n_1882;
input n_3328;
input n_944;
input n_3889;
input n_4256;
input n_4224;
input n_3508;
input n_4024;
input n_2218;
input n_2267;
input n_857;
input n_2636;
input n_1825;
input n_1951;
input n_1883;
input n_2759;
input n_4415;
input n_4702;
input n_4252;
input n_4457;
input n_971;
input n_117;
input n_404;
input n_1393;
input n_2319;
input n_596;
input n_3481;
input n_2808;
input n_2676;
input n_1709;
input n_2679;
input n_4491;
input n_266;
input n_2930;
input n_1838;
input n_3514;
input n_2777;
input n_2434;
input n_4132;
input n_2660;
input n_2611;
input n_4261;
input n_1660;
input n_4886;
input n_4090;
input n_2529;
input n_2698;
input n_1662;
input n_1481;
input n_4001;
input n_3047;
input n_868;
input n_2454;
input n_4371;
input n_914;
input n_4473;
input n_3120;
input n_4007;
input n_1743;
input n_4268;
input n_5028;
input n_1479;
input n_4480;
input n_2350;
input n_3895;
input n_4194;
input n_759;
input n_4824;
input n_1892;
input n_4120;
input n_4427;
input n_3745;
input n_806;
input n_2990;
input n_1766;
input n_324;
input n_1571;
input n_3119;
input n_4142;
input n_1189;
input n_4082;
input n_3479;
input n_4085;
input n_4073;
input n_4260;
input n_1649;
input n_4163;
input n_4439;
input n_2064;
input n_3867;
input n_4372;
input n_3500;
input n_3279;
input n_2621;
input n_5024;
input n_523;
input n_1537;
input n_4262;
input n_2671;
input n_1798;
input n_1790;
input n_4720;
input n_525;
input n_1647;
input n_4685;
input n_2563;
input n_43;
input n_2387;
input n_4334;
input n_1674;
input n_1830;
input n_2073;
input n_4511;
input n_139;
input n_4014;
input n_3144;
input n_4757;
input n_2913;
input n_2336;
input n_254;
input n_1233;
input n_1615;
input n_4175;
input n_2005;
input n_526;
input n_1916;
input n_293;
input n_244;
input n_4648;
input n_47;
input n_1333;
input n_5006;
input n_1443;
input n_946;
input n_1539;
input n_4892;
input n_3823;
input n_1866;
input n_4173;
input n_689;
input n_738;
input n_1624;
input n_4970;
input n_640;
input n_3816;
input n_1279;
input n_4108;
input n_4486;
input n_610;
input n_2960;
input n_1090;
input n_633;
input n_439;
input n_4627;
input n_758;
input n_2290;
input n_2045;
input n_3369;
input n_3783;
input n_2040;
input n_3199;
input n_3843;
input n_1049;
input n_2145;
input n_1639;
input n_1068;
input n_3030;
input n_2580;
input n_3685;
input n_4249;
input n_122;
input n_331;
input n_10;
input n_2039;
input n_4961;
input n_90;
input n_3753;
input n_2035;
input n_4718;
input n_3555;
input n_3579;
input n_2509;
input n_3236;
input n_4317;
input n_1362;
input n_4855;
input n_3969;
input n_2459;
input n_4154;
input n_152;
input n_3396;
input n_1445;
input n_4023;
input n_4420;
input n_1923;
input n_1017;
input n_2116;
input n_1434;
input n_1054;
input n_1828;
input n_2320;
input n_1045;
input n_2038;
input n_2137;
input n_4973;
input n_4640;
input n_2583;
input n_484;
input n_1033;
input n_4396;
input n_636;
input n_4367;
input n_2087;
input n_1009;
input n_109;
input n_454;
input n_1989;
input n_3818;
input n_2523;
input n_255;
input n_4387;
input n_4951;
input n_4453;
input n_4170;
input n_1578;
input n_3719;
input n_1959;
input n_3681;
input n_2737;
input n_1574;
input n_2399;
input n_4308;
input n_2812;
input n_473;
input n_2355;
input n_2133;
input n_1426;
input n_3830;
input n_2585;
input n_2725;
input n_614;
input n_3883;
input n_1355;
input n_2565;
input n_4152;
input n_773;
input n_208;
input n_142;
input n_743;
input n_4392;
input n_4660;
input n_3149;
input n_296;
input n_3268;
input n_4281;
input n_65;
input n_4661;
input n_4200;
input n_3614;
input n_2111;
input n_3301;
input n_3466;
input n_4962;
input n_1237;
input n_2595;
input n_761;
input n_3411;
input n_4958;
input n_329;
input n_4271;
input n_3586;
input n_1390;
input n_30;
input n_4071;
input n_4921;
input n_130;
input n_1980;
input n_3065;
input n_4361;
input n_1093;
input n_263;
input n_4614;
input n_1265;
input n_44;
input n_224;
input n_2681;
input n_3103;
input n_765;
input n_4945;
input n_2424;
input n_4922;
input n_4732;
input n_1015;
input n_1651;
input n_2775;
input n_4693;
input n_511;
input n_358;
input n_1101;
input n_77;
input n_1106;
input n_4326;
input n_3557;
input n_2230;
input n_4744;
input n_2851;
input n_4305;
input n_174;
input n_1455;
input n_767;
input n_2490;
input n_1407;
input n_441;
input n_4213;
input n_2849;
input n_3692;
input n_2204;
input n_365;
input n_4929;
input n_729;
input n_1961;
input n_4964;
input n_911;
input n_1430;
input n_4802;
input n_513;
input n_1354;
input n_4139;
input n_1044;
input n_3029;
input n_2508;
input n_4031;
input n_2416;
input n_623;
input n_3881;
input n_2461;
input n_490;
input n_2243;
input n_4583;
input n_233;
input n_572;
input n_4210;
input n_4666;
input n_2929;
input n_3751;
input n_2555;
input n_2662;
input n_1611;
input n_2368;
input n_2890;
input n_2554;
input n_3698;
input n_3927;
input n_1082;
input n_1840;
input n_4540;
input n_3961;
input n_716;
input n_1630;
input n_4891;
input n_391;
input n_701;
input n_1023;
input n_539;
input n_803;
input n_1092;
input n_3559;
input n_2661;
input n_2572;
input n_3993;
input n_4940;
input n_1056;
input n_3588;
input n_2308;
input n_4590;
input n_4830;
input n_4664;
input n_3860;
input n_1029;
input n_1206;
input n_3160;
input n_2191;
input n_2428;
input n_3847;
input n_4946;
input n_1346;
input n_4906;
input n_2158;
input n_3290;
input n_4663;
input n_1060;
input n_2824;
input n_3033;
input n_3298;
input n_248;
input n_2440;
input n_4883;
input n_1386;
input n_2923;
input n_1442;
input n_4162;
input n_3665;
input n_74;
input n_3264;
input n_2333;
input n_2916;
input n_483;
input n_4297;
input n_1632;
input n_1085;
input n_1066;
input n_3800;
input n_2403;
input n_4608;
input n_46;
input n_2792;
input n_2870;
input n_3991;
input n_378;
input n_1112;
input n_3134;
input n_4172;
input n_4791;
input n_4536;
input n_2463;
input n_4773;
input n_4497;
input n_2472;
input n_4611;
input n_4755;
input n_1768;
input n_2294;
input n_4960;
input n_455;
input n_2993;
input n_1719;
input n_3864;
input n_385;
input n_4658;
input n_2732;
input n_2309;
input n_2948;
input n_1560;
input n_4362;
input n_4306;
input n_2123;
input n_3209;
input n_3504;
input n_2037;
input n_2685;
input n_1953;
input n_4422;
input n_2589;
input n_1301;
input n_1363;
input n_3482;
input n_2233;
input n_1312;
input n_804;
input n_537;
input n_4555;
input n_2827;
input n_153;
input n_1504;
input n_3956;
input n_3572;
input n_250;
input n_992;
input n_4215;
input n_4280;
input n_3375;
input n_4047;
input n_260;
input n_842;
input n_2082;
input n_1643;
input n_3167;
input n_3423;
input n_2362;
input n_2609;
input n_1976;
input n_2223;
input n_3044;
input n_3854;
input n_2468;
input n_1610;
input n_1077;
input n_1422;
input n_3078;
input n_540;
input n_323;
input n_894;
input n_3253;
input n_4027;
input n_831;
input n_2280;
input n_4599;
input n_3363;
input n_4812;
input n_1511;
input n_234;
input n_3689;
input n_2020;
input n_4628;
input n_1881;
input n_988;
input n_2749;
input n_3451;
input n_4873;
input n_4657;
input n_2971;
input n_2311;
input n_3950;
input n_4458;
input n_4121;
input n_1616;
input n_4476;
input n_2298;
input n_4756;
input n_3869;
input n_4307;
input n_4860;
input n_4359;
input n_635;
input n_2303;
input n_2810;
input n_2747;
input n_1848;
input n_2126;
input n_4573;
input n_4118;
input n_4803;
input n_4079;
input n_15;
input n_4091;
input n_681;
input n_1638;
input n_2002;
input n_3712;
input n_2371;
input n_2935;
input n_830;
input n_3085;
input n_1655;
input n_749;
input n_2574;
input n_1134;
input n_1358;
input n_717;
input n_4316;
input n_939;
input n_3697;
input n_482;
input n_1232;
input n_734;
input n_2638;
input n_4044;
input n_4062;
input n_4524;
input n_4843;
input n_3971;
input n_1338;
input n_2016;
input n_1522;
input n_2949;
input n_2711;
input n_338;
input n_1653;
input n_1506;
input n_14;
input n_990;
input n_2867;
input n_1894;
input n_975;
input n_2794;
input n_567;
input n_3145;
input n_3124;
input n_4253;
input n_151;
input n_2608;
input n_2657;
input n_770;
input n_2852;
input n_2392;
input n_711;
input n_85;
input n_3517;
input n_1441;
input n_3100;
input n_2522;
input n_1834;
input n_3758;
input n_3356;
input n_2835;
input n_617;
input n_1572;
input n_1968;
input n_3269;
input n_1516;
input n_3506;
input n_1736;
input n_3605;
input n_2409;
input n_3402;
input n_217;
input n_4679;
input n_4115;
input n_726;
input n_4998;
input n_2988;
input n_1731;
input n_818;
input n_1970;
input n_2766;
input n_2201;
input n_2117;
input n_4167;
input n_1993;
input n_3835;
input n_2205;
input n_1335;
input n_1777;
input n_1957;
input n_3967;
input n_5016;
input n_1912;
input n_3401;
input n_3226;
input n_1410;
input n_707;
input n_3902;
input n_4730;
input n_937;
input n_2779;
input n_1584;
input n_487;
input n_3654;
input n_2164;
input n_2115;
input n_2232;
input n_1302;
input n_1774;
input n_4713;
input n_2811;
input n_3348;
input n_179;
input n_410;
input n_895;
input n_3358;
input n_2121;
input n_1803;
input n_4204;
input n_1543;
input n_1991;
input n_2224;
input n_732;
input n_4743;
input n_500;
input n_1067;
input n_3805;
input n_3825;
input n_148;
input n_3657;
input n_4924;
input n_3928;
input n_4859;
input n_2692;
input n_538;
input n_2008;
input n_4654;
input n_799;
input n_1213;
input n_4733;
input n_3792;
input n_4272;
input n_3974;
input n_3871;
input n_1753;
input n_2283;
input n_3278;
input n_89;
input n_1689;
input n_4269;
input n_4695;
input n_1855;
input n_869;
input n_401;
input n_3312;
input n_1352;
input n_2197;
input n_2199;
input n_3285;
input n_137;
input n_294;
input n_3968;
input n_2228;
input n_4704;
input n_4551;
input n_684;
input n_124;
input n_268;
input n_2421;
input n_2902;
input n_4957;
input n_664;
input n_2480;
input n_235;
input n_2363;
input n_643;
input n_4072;
input n_916;
input n_1115;
input n_4781;
input n_3606;
input n_5004;
input n_2550;
input n_467;
input n_4424;
input n_823;
input n_725;
input n_3055;
input n_3711;
input n_3315;
input n_3172;
input n_3292;
input n_4436;
input n_3878;
input n_4450;
input n_3553;
input n_719;
input n_4746;
input n_1683;
input n_1530;
input n_997;
input n_932;
input n_3131;
input n_1409;
input n_3850;
input n_788;
input n_4459;
input n_1268;
input n_2996;
input n_559;
input n_508;
input n_1320;
input n_4050;
input n_986;
input n_2315;
input n_3228;
input n_1317;
input n_2102;
input n_1063;
input n_4853;
input n_981;
input n_867;
input n_2422;
input n_134;
input n_2239;
input n_587;
input n_2950;
input n_3852;
input n_548;
input n_812;
input n_4520;
input n_518;
input n_2057;
input n_4008;
input n_905;
input n_782;
input n_3858;
input n_1901;
input n_4502;
input n_3032;
input n_4851;
input n_1330;
input n_31;
input n_3072;
input n_3081;
input n_3313;
input n_2710;
input n_1745;
input n_3924;
input n_769;
input n_4571;
input n_2006;
input n_934;
input n_1618;
input n_826;
input n_2343;
input n_3439;
input n_654;
input n_2535;
input n_4205;
input n_2726;
input n_570;
input n_4723;
input n_2799;
input n_4454;
input n_4229;
input n_1083;
input n_4739;
input n_2376;
input n_3017;
input n_787;
input n_2456;
input n_3904;
input n_2678;
input n_95;
input n_4838;
input n_2872;
input n_2451;
input n_522;
input n_4879;
input n_930;
input n_181;
input n_3926;
input n_1962;
input n_3996;
input n_4221;
input n_1577;
input n_2854;
input n_386;
input n_1701;
input n_4181;
input n_1550;
input n_2764;
input n_1498;
input n_4225;
input n_682;
input n_141;
input n_2567;
input n_3102;
input n_922;
input n_1648;
input n_4153;
input n_3627;
input n_4300;
input n_3551;
input n_432;
input n_1769;
input n_4783;
input n_839;
input n_2964;
input n_3769;
input n_2673;
input n_4530;
input n_4267;
input n_140;
input n_2292;
input n_3865;
input n_3859;
input n_3722;
input n_2442;
input n_928;
input n_1943;
input n_3117;
input n_3428;
input n_2961;
input n_3351;
input n_3527;
input n_236;
input n_1396;
input n_1348;
input n_2883;
input n_1752;
input n_4182;
input n_80;
input n_2912;
input n_35;
input n_1315;
input n_4825;
input n_4440;
input n_4549;
input n_1910;
input n_3955;
input n_462;
input n_4565;
input n_4039;
input n_3227;
input n_3300;
input n_4303;
input n_4574;
input n_471;
input n_4839;
input n_1028;
input n_4016;
input n_474;
input n_3435;
input n_3575;
input n_1546;
input n_595;
input n_632;
input n_4231;
input n_3165;
input n_4923;
input n_3652;
input n_4097;
input n_170;
input n_161;
input n_4083;
input n_1937;
input n_81;
input n_4461;
input n_3234;
input n_745;
input n_2381;
input n_3303;
input n_1654;
input n_3916;
input n_2569;
input n_3556;
input n_4101;
input n_2196;
input n_3591;
input n_4273;
input n_3024;
input n_3512;
input n_4939;
input n_4389;
input n_3930;
input n_4448;
input n_1325;
input n_1595;
input n_2161;
input n_2404;
input n_2083;
input n_2503;
input n_1540;
input n_1936;
input n_2027;
input n_453;
input n_403;
input n_2642;
input n_720;
input n_2500;
input n_1918;
input n_863;
input n_4831;
input n_2513;
input n_2695;
input n_3480;
input n_3057;
input n_3194;
input n_2414;
input n_1402;
input n_3662;
input n_4319;
input n_644;
input n_2229;
input n_1397;
input n_4596;
input n_2004;
input n_251;
input n_3694;
input n_2586;
input n_4726;
input n_1398;
input n_1879;
input n_4751;
input n_4222;
input n_1196;
input n_2274;
input n_2972;
input n_3225;
input n_334;
input n_811;
input n_175;
input n_4119;
input n_3799;
input n_4298;
input n_4474;
input n_1089;
input n_1004;
input n_242;
input n_2511;
input n_1681;
input n_3383;
input n_3585;
input n_2975;
input n_438;
input n_5029;
input n_2704;
input n_4214;
input n_4884;
input n_533;
input n_4366;
input n_1251;
input n_4009;
input n_278;
input n_4580;
input n_1263;
input n_611;
input n_1126;
input n_4129;
input n_4871;
input n_2617;
input n_4999;
input n_1859;
input n_1677;
input n_2955;
input n_4112;
input n_4337;
input n_4138;
input n_552;
input n_1528;
input n_1292;
input n_2520;
input n_1198;
input n_956;
input n_423;
input n_2134;
input n_4236;
input n_2185;
input n_3270;
input n_2143;
input n_5002;
input n_3595;
input n_1347;
input n_4238;
input n_1451;
input n_1022;
input n_1545;
input n_2374;
input n_173;
input n_859;
input n_1947;
input n_2114;
input n_3571;
input n_854;
input n_1799;
input n_2396;
input n_4734;
input n_674;
input n_1939;
input n_2486;
input n_516;
input n_4635;
input n_1152;
input n_3501;
input n_1869;
input n_4013;
input n_606;
input n_3039;
input n_275;
input n_2011;
input n_4242;
input n_6;
input n_4984;
input n_3851;
input n_2543;
input n_150;
input n_3036;
input n_1896;
input n_3180;
input n_191;
input n_1705;
input n_659;
input n_4561;
input n_2639;
input n_3325;
input n_3107;
input n_4021;
input n_3880;
input n_1261;
input n_938;
input n_3186;
input n_4955;
input n_1154;
input n_4501;
input n_3696;
input n_406;
input n_546;
input n_1280;
input n_3650;
input n_291;
input n_2761;
input n_257;
input n_3157;
input n_709;
input n_2537;
input n_2144;
input n_920;
input n_2515;
input n_2466;
input n_2652;
input n_2635;
input n_4197;
input n_4829;
input n_976;
input n_1949;
input n_1946;
input n_2936;
input n_775;
input n_1484;
input n_1328;
input n_4715;
input n_2141;
input n_4369;
input n_4543;
input n_2099;
input n_4941;
input n_1831;
input n_1598;
input n_4394;
input n_1850;
input n_163;
input n_243;
input n_1749;
input n_59;
input n_3101;
input n_3669;
input n_215;
input n_350;
input n_196;
input n_2663;
input n_1394;
input n_580;
input n_2693;
input n_3798;
input n_4065;
input n_4944;
input n_926;
input n_2180;
input n_2249;
input n_4135;
input n_1218;
input n_2632;
input n_475;
input n_1547;
input n_777;
input n_1755;
input n_415;
input n_485;
input n_958;
input n_2908;
input n_3744;
input n_4263;
input n_1862;
input n_1239;
input n_2915;
input n_2300;
input n_3291;
input n_4716;
input n_4942;
input n_164;
input n_2432;
input n_1521;
input n_3405;
input n_214;
input n_4745;
input n_2337;
input n_1167;
input n_1384;
input n_3907;
input n_923;
input n_4629;
input n_213;
input n_2932;
input n_2980;
input n_464;
input n_1069;
input n_3306;
input n_1784;
input n_4857;
input n_3136;
input n_4080;
input n_4226;
input n_4741;
input n_2101;
input n_1471;
input n_1986;
input n_4752;
input n_1750;
input n_1459;
input n_460;
input n_3986;
input n_4376;
input n_4753;
input n_571;
input n_4552;
input n_3885;
input n_2713;
input n_2644;
input n_1197;
input n_2951;
input n_3008;
input n_3709;
input n_1039;
input n_2214;
input n_34;
input n_2055;
input n_3427;
input n_4067;
input n_1403;
input n_4042;
input n_4176;
input n_4385;
input n_3320;
input n_5009;
input n_2688;
input n_1202;
input n_1463;
input n_3651;
input n_4333;
input n_3359;
input n_2865;
input n_349;
input n_2706;
input n_3676;
input n_4375;
input n_4788;
input n_4717;
input n_4986;
input n_3789;
input n_2152;
input n_3598;
input n_627;
input n_4815;
input n_4246;
input n_3580;
input n_2139;
input n_4609;
input n_91;
input n_2674;
input n_1565;
input n_4088;
input n_3682;
input n_4357;
input n_3371;
input n_1809;
input n_4462;
input n_4472;
input n_647;
input n_3433;
input n_1072;
input n_2305;
input n_2450;
input n_561;
input n_3447;
input n_3305;
input n_4148;
input n_4151;
input n_1712;
input n_3528;
input n_4373;
input n_4934;
input n_2322;
input n_2271;
input n_2625;
input n_4630;
input n_4643;
input n_4331;
input n_3989;
input n_4475;
input n_4846;
input n_3804;
input n_4344;
input n_1775;
input n_3296;
input n_1368;
input n_2762;
input n_4683;
input n_728;
input n_1162;
input n_272;
input n_1847;
input n_2767;
input n_2603;
input n_3116;
input n_1884;
input n_3602;
input n_2967;
input n_409;
input n_887;
input n_1905;
input n_2553;
input n_3706;
input n_2195;
input n_300;
input n_3923;
input n_931;
input n_599;
input n_4696;
input n_2626;
input n_3441;
input n_1978;
input n_1544;
input n_639;
input n_1629;
input n_2801;
input n_4011;
input n_4905;
input n_121;
input n_2763;
input n_360;
input n_2825;
input n_3643;
input n_4876;
input n_1997;
input n_3748;
input n_1477;
input n_3142;
input n_4278;
input n_1635;
input n_4623;
input n_187;
input n_4910;
input n_2690;
input n_4410;
input n_3370;
input n_2215;
input n_1259;
input n_4553;
input n_706;
input n_746;
input n_784;
input n_3978;
input n_110;
input n_4809;
input n_1244;
input n_1925;
input n_3660;
input n_1815;
input n_1788;
input n_2491;
input n_913;
input n_3833;
input n_865;
input n_61;
input n_697;
input n_1222;
input n_75;
input n_1679;
input n_4841;
input n_776;
input n_2022;
input n_3814;
input n_1415;
input n_2592;
input n_2838;
input n_4842;
input n_4911;
input n_4340;
input n_3513;
input n_3133;
input n_4645;
input n_1191;
input n_2992;
input n_3725;
input n_1833;
input n_4920;
input n_4972;
input n_2517;
input n_284;
input n_3128;
input n_744;
input n_629;
input n_2631;
input n_2178;
input n_1767;
input n_23;
input n_1529;
input n_2469;
input n_3355;
input n_604;
input n_2007;
input n_3917;
input n_3942;
input n_2736;
input n_3765;
input n_498;
input n_3000;
input n_252;
input n_624;
input n_1010;
input n_1231;
input n_739;
input n_1406;
input n_3108;
input n_3111;
input n_1837;
input n_1839;
input n_4557;
input n_4451;
input n_2875;
input n_936;
input n_1500;
input n_3844;
input n_3280;
input n_4054;
input n_3471;
input n_259;
input n_448;
input n_999;
input n_3205;
input n_2046;
input n_2848;
input n_2741;
input n_3003;
input n_3610;
input n_1933;
input n_1656;
input n_3564;
input n_1158;
input n_3988;
input n_563;
input n_3457;
input n_204;
input n_1678;
input n_4324;
input n_4821;
input n_1871;
input n_3630;
input n_3271;
input n_4771;
input n_908;
input n_4086;
input n_2412;
input n_4814;
input n_724;
input n_1781;
input n_2084;
input n_3648;
input n_3075;
input n_3173;
input n_4692;
input n_456;
input n_959;
input n_3031;
input n_3701;
input n_1773;
input n_3243;
input n_1169;
input n_45;
input n_2666;
input n_3385;
input n_2171;
input n_4708;
input n_2768;
input n_2314;
input n_4826;
input n_2420;
input n_3343;
input n_514;
input n_1079;
input n_1593;
input n_3767;
input n_442;
input n_2299;
input n_131;
input n_2540;
input n_2873;
input n_4589;
input n_4578;
input n_1640;
input n_2162;
input n_2847;
input n_1148;
input n_2051;
input n_3221;
input n_742;
input n_750;
input n_2168;
input n_2790;
input n_3629;
input n_3021;
input n_185;
input n_2359;
input n_3674;
input n_3502;
input n_3098;
input n_1383;
input n_5013;
input n_2312;
input n_3015;
input n_1171;
input n_1920;
input n_1065;
input n_4147;
input n_2048;
input n_3607;
input n_4925;
input n_1921;
input n_1309;
input n_4974;
input n_355;
input n_1800;
input n_1548;
input n_4932;
input n_1421;
input n_4510;
input n_2571;
input n_1286;
input n_1177;
input n_3276;
input n_3787;
input n_2124;
input n_613;
input n_1119;
input n_1240;
input n_3827;
input n_829;
input n_2519;
input n_3354;
input n_2724;
input n_4447;
input n_4285;
input n_4651;
input n_361;
input n_700;
input n_573;
input n_4818;
input n_4514;
input n_388;
input n_1366;
input n_4800;
input n_3960;
input n_3248;
input n_2277;
input n_1568;
input n_2110;
input n_274;
input n_582;
input n_1332;
input n_4433;
input n_2879;
input n_73;
input n_2474;
input n_19;
input n_2090;
input n_3153;
input n_512;
input n_1591;
input n_2033;
input n_4341;
input n_1682;
input n_4312;
input n_2628;
input n_3399;
input n_1249;
input n_1111;
input n_25;
input n_2132;
input n_2400;
input n_4633;
input n_609;
input n_3838;
input n_1909;
input n_4277;
input n_112;
input n_4140;
input n_3675;
input n_1140;
input n_891;
input n_3387;
input n_4662;
input n_3779;
input n_2464;
input n_2831;
input n_102;
input n_1456;
input n_4882;
input n_4993;
input n_2365;
input n_4832;
input n_4207;
input n_987;
input n_4545;
input n_3037;
input n_261;
input n_4868;
input n_1885;
input n_2452;
input n_3925;
input n_2176;
input n_1816;
input n_4059;
input n_2455;
input n_4595;
input n_1849;
input n_1131;
input n_2467;
input n_1094;
input n_2288;
input n_4063;
input n_346;
input n_1209;
input n_3592;
input n_4650;
input n_602;
input n_4888;
input n_1435;
input n_879;
input n_3394;
input n_4874;
input n_3793;
input n_16;
input n_4669;
input n_405;
input n_4339;
input n_1645;
input n_4041;
input n_2858;
input n_4060;
input n_996;
input n_2658;
input n_1717;
input n_2895;
input n_2128;
input n_3097;
input n_120;
input n_327;
input n_135;
input n_4541;
input n_3824;
input n_3388;
input n_4494;
input n_3059;
input n_3465;
input n_1316;
input n_4796;
input n_1438;
input n_3589;
input n_62;
input n_952;
input n_2534;
input n_1229;
input n_4799;
input n_3449;
input n_2694;
input n_2198;
input n_2610;
input n_2989;
input n_2789;
input n_4775;
input n_2216;
input n_531;
input n_1897;
input n_764;
input n_1424;
input n_162;
input n_2933;
input n_4381;
input n_4266;
input n_3886;
input n_4455;
input n_2328;
input n_199;
input n_4248;
input n_4754;
input n_4554;
input n_4845;
input n_3053;
input n_1299;
input n_3893;
input n_1141;
input n_2465;
input n_3548;
input n_4585;
input n_418;
input n_315;
input n_451;
input n_1699;
input n_3334;
input n_2541;
input n_4383;
input n_1139;
input n_57;
input n_397;
input n_1432;
input n_3875;
input n_4003;
input n_2402;
input n_4301;
input n_841;
input n_1050;
input n_4586;
input n_1954;
input n_4048;
input n_1844;
input n_3777;
input n_4784;
input n_2999;
input n_1644;
input n_4046;
input n_1974;
input n_2086;
input n_3537;
input n_3080;
input n_4199;
input n_2701;
input n_3362;
input n_1631;
input n_3105;
input n_1179;
input n_753;
input n_1048;
input n_4286;
input n_2556;
input n_2269;
input n_3274;
input n_3041;
input n_4470;
input n_2236;
input n_330;
input n_2816;
input n_692;
input n_820;
input n_1911;
input n_3616;
input n_2460;
input n_4058;
input n_3664;
input n_4188;
input n_1668;
input n_3913;
input n_3417;
input n_1143;
input n_1579;
input n_4034;
input n_1688;
input n_492;
input n_3327;
input n_4689;
input n_341;
input n_3067;
input n_2755;
input n_543;
input n_3237;
input n_1992;
input n_4402;
input n_4239;
input n_3400;
input n_449;
input n_4550;
input n_1214;
input n_1342;
input n_1400;
input n_3382;
input n_3574;
input n_2169;
input n_1557;
input n_4201;
input n_618;
input n_896;
input n_3316;
input n_356;
input n_3099;
input n_3704;
input n_2596;
input n_1730;
input n_3603;
input n_4123;
input n_2192;
input n_964;
input n_3633;
input n_4479;
input n_1373;
input n_2670;
input n_5;
input n_1646;
input n_1307;
input n_4416;
input n_3372;
input n_4539;
input n_814;
input n_2707;
input n_2471;
input n_1472;
input n_1671;
input n_3230;
input n_1062;
input n_3342;
input n_4682;
input n_3708;
input n_1204;
input n_3729;
input n_4978;
input n_4690;
input n_4437;
input n_3861;
input n_4736;
input n_3780;
input n_783;
input n_1928;
input n_1188;
input n_3957;
input n_3848;
input n_41;
input n_4284;
input n_2600;
input n_3919;
input n_336;
input n_3608;
input n_510;
input n_216;
input n_4513;
input n_3233;
input n_3829;
input n_3177;
input n_4053;
input n_2352;
input n_4040;
input n_2207;
input n_2619;
input n_2444;
input n_241;
input n_1110;
input n_3123;
input n_1088;
input n_3393;
input n_638;
input n_866;
input n_4887;
input n_4617;
input n_3520;
input n_2492;
input n_249;
input n_577;
input n_4005;
input n_1687;
input n_1637;
input n_4904;
input n_1419;
input n_693;
input n_4792;
input n_3578;
input n_3812;
input n_1886;
input n_1389;
input n_1256;
input n_4980;
input n_1465;
input n_4290;
input n_306;
input n_1375;
input n_3727;
input n_3774;
input n_3093;
input n_1843;
input n_3061;
input n_1597;
input n_1659;
input n_2431;
input n_1371;
input n_4956;
input n_2206;
input n_3182;
input n_2564;
input n_4947;
input n_876;
input n_4656;
input n_1190;
input n_3896;
input n_3958;
input n_3450;
input n_966;
input n_4729;
input n_4987;
input n_4971;
input n_1116;
input n_2000;
input n_1212;
input n_2074;
input n_206;
input n_3174;
input n_982;
input n_1453;
input n_2217;
input n_1183;
input n_3398;
input n_2307;
input n_3408;
input n_899;
input n_2722;
input n_2640;
input n_4823;
input n_4875;
input n_1628;
input n_3432;
input n_1514;
input n_1771;
input n_557;
input n_1005;
input n_607;
input n_679;
input n_710;
input n_3090;
input n_527;
input n_1168;
input n_2437;
input n_3762;
input n_2445;
input n_1427;
input n_108;
input n_1835;
input n_66;
input n_177;
input n_1988;
input n_1853;
input n_1356;
input n_1787;
input n_4137;
input n_2634;
input n_4529;
input n_910;
input n_4323;
input n_3034;
input n_2212;
input n_3972;
input n_125;
input n_529;
input n_126;
input n_202;
input n_3308;
input n_791;
input n_1533;
input n_5036;
input n_4772;
input n_3467;
input n_4322;
input n_1720;
input n_2830;
input n_4354;
input n_159;
input n_4653;
input n_2354;
input n_2246;
input n_4677;
input n_3901;
input n_715;
input n_1480;
input n_3757;
input n_3381;
input n_1782;
input n_2245;
input n_4909;
input n_1524;
input n_1485;
input n_115;
input n_810;
input n_2965;
input n_416;
input n_3635;
input n_5022;
input n_5005;
input n_1144;
input n_2814;
input n_1570;
input n_3882;
input n_3046;
input n_1170;
input n_305;
input n_2213;
input n_3826;
input n_3211;
input n_2211;
input n_2095;
input n_3121;
input n_4634;
input n_3337;
input n_2527;
input n_855;
input n_1461;
input n_3204;
input n_2136;
input n_1273;
input n_1822;
input n_4952;
input n_3005;
input n_1235;
input n_4380;
input n_980;
input n_698;
input n_3129;
input n_4126;
input n_1282;
input n_1783;
input n_2601;
input n_3043;
input n_998;
input n_3802;
input n_2375;
input n_4506;
input n_4880;
input n_1907;
input n_501;
input n_2686;
input n_2344;
input n_3892;
input n_4896;
input n_1417;
input n_1295;
input n_1985;
input n_2107;
input n_3219;
input n_2906;
input n_4943;
input n_382;
input n_2187;
input n_1762;
input n_1013;
input n_718;
input n_3023;
input n_4193;
input n_4075;
input n_3104;
input n_612;
input n_4737;
input n_3647;
input n_825;
input n_2819;
input n_506;
input n_737;
input n_3609;
input n_4136;
input n_1715;
input n_1952;
input n_4393;
input n_3720;
input n_4535;
input n_733;
input n_1922;
input n_2560;
input n_4522;
input n_4794;
input n_3959;
input n_63;
input n_792;
input n_3140;
input n_3724;
input n_298;
input n_2104;
input n_505;
input n_3011;
input n_4196;
input n_1425;
input n_4592;
input n_4675;
input n_3069;
input n_4370;
input n_1900;
input n_1620;
input n_3084;
input n_1727;
input n_2735;
input n_2497;
input n_3412;
input n_1995;
input n_2411;
input n_1046;
input n_3761;
input n_4889;
input n_2014;
input n_2986;
input n_1641;
input n_1361;
input n_3184;
input n_4828;
input n_4558;
input n_2172;
input n_4722;
input n_1129;
input n_158;
input n_3626;
input n_4768;
input n_4100;
input n_961;
input n_2250;
input n_276;
input n_1225;
input n_169;
input n_400;
input n_4092;
input n_3908;
input n_2423;
input n_3671;
input n_994;
input n_3344;
input n_2194;
input n_848;
input n_4465;
input n_3302;
input n_1223;
input n_2680;
input n_1567;
input n_3122;
input n_4808;
input n_3842;
input n_145;
input n_3265;
input n_1857;
input n_4482;
input n_2041;
input n_631;
input n_479;
input n_1797;
input n_2957;
input n_2357;
input n_1250;
input n_3309;
input n_608;
input n_772;
input n_3260;
input n_4926;
input n_3357;
input n_1589;
input n_4116;
input n_1086;
input n_2570;
input n_1858;
input n_1619;
input n_2815;
input n_3754;
input n_4612;
input n_1469;
input n_2744;
input n_4287;
input n_2397;
input n_384;
input n_2208;
input n_3063;
input n_3617;
input n_333;
input n_1298;
input n_1652;
input n_4516;
input n_3794;
input n_2809;
input n_2050;
input n_4505;
input n_1676;
input n_258;
input n_1113;
input n_29;
input n_1277;
input n_2591;
input n_188;
input n_3384;
input n_852;
input n_4602;
input n_4449;
input n_1864;
input n_463;
input n_502;
input n_466;
input n_420;
input n_1337;
input n_4445;
input n_699;
input n_1627;
input n_1245;
input n_4870;
input n_2438;
input n_465;
input n_2832;
input n_362;
input n_1321;
input n_1975;
input n_2296;
input n_273;
input n_3181;
input n_616;
input n_2278;
input n_4915;
input n_2135;
input n_3493;
input n_3323;
input n_2734;
input n_4914;
input n_1076;
input n_2823;
input n_1408;
input n_494;
input n_1761;
input n_730;
input n_354;
input n_795;
input n_4345;
input n_180;
input n_3281;
input n_656;
input n_3307;
input n_1606;
input n_1220;
input n_1694;
input n_4318;
input n_2485;
input n_2655;
input n_60;
input n_4185;
input n_4797;
input n_2366;
input n_1526;
input n_3997;
input n_1604;
input n_1275;
input n_4032;
input n_1764;
input n_3582;
input n_712;
input n_1583;
input n_2826;
input n_3539;
input n_1042;
input n_285;
input n_412;
input n_4343;
input n_1493;
input n_4212;
input n_4124;
input n_4492;
input n_2708;
input n_4994;
input n_4245;
input n_4364;
input n_4928;
input n_2225;
input n_1507;
input n_4378;
input n_2383;
input n_1996;
input n_597;
input n_3406;
input n_3604;
input n_3853;
input n_4216;
input n_2019;
input n_1340;
input n_1558;
input n_2166;
input n_2938;
input n_4309;
input n_3594;
input n_262;
input n_1704;
input n_3721;
input n_1254;
input n_1026;
input n_2026;
input n_1234;
input n_2109;
input n_364;
input n_2013;
input n_20;
input n_1990;
input n_1032;
input n_2614;
input n_2991;
input n_2242;
input n_2752;
input n_2894;
input n_3473;
input n_4560;
input n_2839;
input n_1588;
input n_2237;
input n_3463;
input n_3699;
input n_3360;
input n_2524;
input n_3873;
input n_3693;
input n_2728;
input n_3857;

output n_18332;

wire n_13115;
wire n_6643;
wire n_18022;
wire n_6122;
wire n_10564;
wire n_13903;
wire n_7981;
wire n_9936;
wire n_5567;
wire n_15472;
wire n_12148;
wire n_16520;
wire n_14870;
wire n_15741;
wire n_9194;
wire n_15969;
wire n_12407;
wire n_6579;
wire n_15974;
wire n_9325;
wire n_7164;
wire n_16559;
wire n_17478;
wire n_10794;
wire n_5287;
wire n_6546;
wire n_12872;
wire n_13683;
wire n_14881;
wire n_15306;
wire n_9655;
wire n_15349;
wire n_14101;
wire n_15948;
wire n_5484;
wire n_10515;
wire n_11207;
wire n_11326;
wire n_5978;
wire n_8174;
wire n_5161;
wire n_15269;
wire n_5776;
wire n_14036;
wire n_13241;
wire n_6551;
wire n_13217;
wire n_16007;
wire n_5512;
wire n_14764;
wire n_10793;
wire n_14635;
wire n_5207;
wire n_12853;
wire n_17997;
wire n_9044;
wire n_6786;
wire n_12327;
wire n_13927;
wire n_17360;
wire n_18151;
wire n_7206;
wire n_7303;
wire n_10552;
wire n_9083;
wire n_12215;
wire n_13112;
wire n_15682;
wire n_16276;
wire n_14631;
wire n_8363;
wire n_9408;
wire n_13779;
wire n_12975;
wire n_17821;
wire n_11802;
wire n_7710;
wire n_8383;
wire n_5282;
wire n_10885;
wire n_11583;
wire n_11349;
wire n_16000;
wire n_8328;
wire n_13499;
wire n_7461;
wire n_12641;
wire n_8060;
wire n_6649;
wire n_9331;
wire n_14203;
wire n_14939;
wire n_7154;
wire n_8551;
wire n_14264;
wire n_17586;
wire n_13768;
wire n_8002;
wire n_12924;
wire n_15935;
wire n_10108;
wire n_8594;
wire n_6810;
wire n_13386;
wire n_7660;
wire n_14070;
wire n_12071;
wire n_6276;
wire n_11016;
wire n_6072;
wire n_12738;
wire n_16752;
wire n_8976;
wire n_17501;
wire n_8617;
wire n_14144;
wire n_10883;
wire n_7686;
wire n_16119;
wire n_17921;
wire n_10117;
wire n_15940;
wire n_16152;
wire n_12139;
wire n_9846;
wire n_12328;
wire n_17049;
wire n_8603;
wire n_17014;
wire n_7024;
wire n_12493;
wire n_14762;
wire n_16301;
wire n_7205;
wire n_16997;
wire n_9204;
wire n_6742;
wire n_9769;
wire n_11342;
wire n_15734;
wire n_16153;
wire n_9312;
wire n_16454;
wire n_13493;
wire n_10363;
wire n_16208;
wire n_8319;
wire n_6694;
wire n_9610;
wire n_15411;
wire n_7616;
wire n_17714;
wire n_7486;
wire n_13220;
wire n_15406;
wire n_13822;
wire n_11450;
wire n_14287;
wire n_8244;
wire n_12028;
wire n_9273;
wire n_12357;
wire n_16963;
wire n_6580;
wire n_6090;
wire n_12515;
wire n_7010;
wire n_17679;
wire n_11678;
wire n_17857;
wire n_5480;
wire n_6549;
wire n_8105;
wire n_17947;
wire n_14471;
wire n_6913;
wire n_7867;
wire n_13158;
wire n_10756;
wire n_7315;
wire n_11801;
wire n_14435;
wire n_13516;
wire n_16013;
wire n_11653;
wire n_7004;
wire n_8961;
wire n_13415;
wire n_16240;
wire n_7772;
wire n_10761;
wire n_18152;
wire n_11299;
wire n_5402;
wire n_13146;
wire n_17017;
wire n_5851;
wire n_13889;
wire n_5509;
wire n_13775;
wire n_9773;
wire n_15311;
wire n_8574;
wire n_16846;
wire n_11089;
wire n_14045;
wire n_11077;
wire n_8864;
wire n_15797;
wire n_16498;
wire n_16602;
wire n_12861;
wire n_9173;
wire n_12709;
wire n_7641;
wire n_16910;
wire n_11296;
wire n_17191;
wire n_15567;
wire n_5154;
wire n_9363;
wire n_8681;
wire n_7468;
wire n_9796;
wire n_5469;
wire n_6431;
wire n_11800;
wire n_13906;
wire n_14721;
wire n_16313;
wire n_12462;
wire n_12012;
wire n_5744;
wire n_14714;
wire n_12266;
wire n_9049;
wire n_17526;
wire n_17244;
wire n_11947;
wire n_5453;
wire n_14411;
wire n_11917;
wire n_15377;
wire n_14537;
wire n_7861;
wire n_9907;
wire n_16655;
wire n_8413;
wire n_9738;
wire n_15543;
wire n_5202;
wire n_5648;
wire n_10745;
wire n_13748;
wire n_14898;
wire n_16663;
wire n_18100;
wire n_13178;
wire n_7667;
wire n_13072;
wire n_6931;
wire n_9539;
wire n_14270;
wire n_8114;
wire n_15657;
wire n_17833;
wire n_9811;
wire n_12970;
wire n_6618;
wire n_13771;
wire n_6408;
wire n_9993;
wire n_17870;
wire n_9208;
wire n_17245;
wire n_14729;
wire n_10421;
wire n_7523;
wire n_16256;
wire n_16388;
wire n_14800;
wire n_17914;
wire n_8706;
wire n_13000;
wire n_16722;
wire n_5922;
wire n_16182;
wire n_17101;
wire n_8158;
wire n_11594;
wire n_15727;
wire n_12100;
wire n_14959;
wire n_6698;
wire n_15990;
wire n_9500;
wire n_15484;
wire n_18109;
wire n_16017;
wire n_8104;
wire n_10399;
wire n_5848;
wire n_10420;
wire n_12575;
wire n_16295;
wire n_11635;
wire n_17436;
wire n_17912;
wire n_16689;
wire n_18117;
wire n_5406;
wire n_12501;
wire n_17124;
wire n_6085;
wire n_14408;
wire n_15805;
wire n_12819;
wire n_7421;
wire n_7306;
wire n_11505;
wire n_14403;
wire n_8819;
wire n_15753;
wire n_10535;
wire n_6214;
wire n_7493;
wire n_10360;
wire n_12027;
wire n_16311;
wire n_9420;
wire n_7804;
wire n_8089;
wire n_12111;
wire n_12075;
wire n_12078;
wire n_13401;
wire n_9557;
wire n_13708;
wire n_9382;
wire n_5241;
wire n_12175;
wire n_16558;
wire n_6939;
wire n_12604;
wire n_7528;
wire n_16275;
wire n_16383;
wire n_11615;
wire n_10307;
wire n_14519;
wire n_10781;
wire n_8262;
wire n_8290;
wire n_9206;
wire n_11507;
wire n_7562;
wire n_12626;
wire n_11497;
wire n_10193;
wire n_9388;
wire n_14611;
wire n_11541;
wire n_5661;
wire n_8885;
wire n_6991;
wire n_5562;
wire n_16192;
wire n_9772;
wire n_10437;
wire n_12142;
wire n_16390;
wire n_10430;
wire n_8147;
wire n_6586;
wire n_11111;
wire n_11354;
wire n_16764;
wire n_10177;
wire n_13782;
wire n_8310;
wire n_11052;
wire n_5398;
wire n_13875;
wire n_6096;
wire n_15548;
wire n_17791;
wire n_6707;
wire n_14170;
wire n_10175;
wire n_5852;
wire n_12767;
wire n_6920;
wire n_13110;
wire n_6868;
wire n_17502;
wire n_18260;
wire n_9311;
wire n_17685;
wire n_16339;
wire n_12754;
wire n_5144;
wire n_17297;
wire n_9422;
wire n_16942;
wire n_14892;
wire n_16514;
wire n_10672;
wire n_9040;
wire n_9795;
wire n_14336;
wire n_15551;
wire n_8380;
wire n_16326;
wire n_9027;
wire n_15813;
wire n_8962;
wire n_12225;
wire n_7402;
wire n_5577;
wire n_10626;
wire n_7592;
wire n_15697;
wire n_11316;
wire n_7152;
wire n_16452;
wire n_14579;
wire n_18237;
wire n_15312;
wire n_6512;
wire n_9966;
wire n_11272;
wire n_13571;
wire n_13096;
wire n_15154;
wire n_16324;
wire n_8126;
wire n_5689;
wire n_13087;
wire n_17635;
wire n_13309;
wire n_10392;
wire n_5894;
wire n_12670;
wire n_12152;
wire n_15336;
wire n_7801;
wire n_7992;
wire n_11588;
wire n_11689;
wire n_9161;
wire n_10231;
wire n_7463;
wire n_12101;
wire n_17010;
wire n_8556;
wire n_10316;
wire n_9369;
wire n_13753;
wire n_9033;
wire n_18035;
wire n_13542;
wire n_8305;
wire n_10683;
wire n_6725;
wire n_14109;
wire n_7613;
wire n_16557;
wire n_16683;
wire n_9429;
wire n_12576;
wire n_17265;
wire n_7083;
wire n_7086;
wire n_7349;
wire n_14458;
wire n_13610;
wire n_16687;
wire n_15343;
wire n_10514;
wire n_6464;
wire n_8317;
wire n_10730;
wire n_10958;
wire n_13095;
wire n_10562;
wire n_11273;
wire n_11962;
wire n_18060;
wire n_14856;
wire n_15008;
wire n_13706;
wire n_8653;
wire n_7647;
wire n_5825;
wire n_7779;
wire n_7712;
wire n_14792;
wire n_11303;
wire n_14711;
wire n_7316;
wire n_6820;
wire n_12224;
wire n_5343;
wire n_9780;
wire n_10252;
wire n_12237;
wire n_10438;
wire n_9824;
wire n_6098;
wire n_7019;
wire n_12751;
wire n_13612;
wire n_16487;
wire n_6686;
wire n_16876;
wire n_17230;
wire n_11664;
wire n_10523;
wire n_15481;
wire n_11720;
wire n_5062;
wire n_10202;
wire n_11398;
wire n_15106;
wire n_11659;
wire n_6561;
wire n_6584;
wire n_7452;
wire n_5184;
wire n_7956;
wire n_8939;
wire n_17587;
wire n_12824;
wire n_15823;
wire n_9489;
wire n_8604;
wire n_16656;
wire n_7323;
wire n_14605;
wire n_14405;
wire n_15932;
wire n_11365;
wire n_13755;
wire n_12269;
wire n_17998;
wire n_7195;
wire n_6701;
wire n_13243;
wire n_17269;
wire n_10988;
wire n_7478;
wire n_11836;
wire n_16030;
wire n_6769;
wire n_7683;
wire n_13131;
wire n_16782;
wire n_6592;
wire n_11150;
wire n_5686;
wire n_16822;
wire n_12298;
wire n_12019;
wire n_13457;
wire n_5463;
wire n_14263;
wire n_14824;
wire n_5236;
wire n_7903;
wire n_6062;
wire n_6191;
wire n_11003;
wire n_12299;
wire n_16684;
wire n_9625;
wire n_8440;
wire n_15995;
wire n_16956;
wire n_10980;
wire n_5433;
wire n_10367;
wire n_8525;
wire n_8416;
wire n_13734;
wire n_13219;
wire n_17273;
wire n_9570;
wire n_12232;
wire n_9368;
wire n_15040;
wire n_15981;
wire n_8064;
wire n_13547;
wire n_7575;
wire n_5909;
wire n_15564;
wire n_17637;
wire n_8879;
wire n_10664;
wire n_13458;
wire n_9115;
wire n_9694;
wire n_9367;
wire n_17166;
wire n_6043;
wire n_15544;
wire n_16780;
wire n_17427;
wire n_11520;
wire n_13747;
wire n_12812;
wire n_16341;
wire n_16314;
wire n_6271;
wire n_7171;
wire n_11099;
wire n_7701;
wire n_13223;
wire n_5315;
wire n_11859;
wire n_13416;
wire n_8931;
wire n_18081;
wire n_15290;
wire n_5348;
wire n_5055;
wire n_8214;
wire n_9072;
wire n_14973;
wire n_16025;
wire n_6793;
wire n_7873;
wire n_9612;
wire n_16154;
wire n_15762;
wire n_12777;
wire n_9971;
wire n_13620;
wire n_8729;
wire n_14886;
wire n_7127;
wire n_16141;
wire n_5397;
wire n_6550;
wire n_17852;
wire n_10575;
wire n_17744;
wire n_11746;
wire n_16883;
wire n_5709;
wire n_7568;
wire n_10803;
wire n_15331;
wire n_15503;
wire n_6021;
wire n_16179;
wire n_9720;
wire n_5695;
wire n_9213;
wire n_7814;
wire n_10187;
wire n_10400;
wire n_14227;
wire n_14345;
wire n_11330;
wire n_17318;
wire n_14698;
wire n_10778;
wire n_17799;
wire n_18135;
wire n_15896;
wire n_5860;
wire n_6926;
wire n_11121;
wire n_9607;
wire n_7589;
wire n_6928;
wire n_7965;
wire n_13283;
wire n_15911;
wire n_15857;
wire n_5862;
wire n_8228;
wire n_6304;
wire n_8210;
wire n_5189;
wire n_10586;
wire n_17957;
wire n_6956;
wire n_10040;
wire n_16638;
wire n_5381;
wire n_13555;
wire n_7026;
wire n_6782;
wire n_13582;
wire n_5854;
wire n_11911;
wire n_5516;
wire n_15316;
wire n_17603;
wire n_9554;
wire n_15281;
wire n_9262;
wire n_17261;
wire n_11599;
wire n_16376;
wire n_15649;
wire n_12412;
wire n_16731;
wire n_8387;
wire n_7002;
wire n_12782;
wire n_17593;
wire n_8898;
wire n_8410;
wire n_14852;
wire n_7141;
wire n_14019;
wire n_10935;
wire n_13809;
wire n_5936;
wire n_16578;
wire n_6126;
wire n_9761;
wire n_12284;
wire n_17612;
wire n_12612;
wire n_11102;
wire n_8795;
wire n_9649;
wire n_10164;
wire n_10269;
wire n_11039;
wire n_8501;
wire n_12567;
wire n_15622;
wire n_10401;
wire n_14228;
wire n_15264;
wire n_6598;
wire n_9529;
wire n_6027;
wire n_9254;
wire n_15205;
wire n_15345;
wire n_11535;
wire n_6342;
wire n_14854;
wire n_14627;
wire n_6638;
wire n_10651;
wire n_16183;
wire n_16732;
wire n_7308;
wire n_5254;
wire n_12180;
wire n_15828;
wire n_17822;
wire n_6900;
wire n_8953;
wire n_14016;
wire n_13295;
wire n_12731;
wire n_13644;
wire n_9726;
wire n_12153;
wire n_8823;
wire n_11686;
wire n_10851;
wire n_7264;
wire n_14046;
wire n_11730;
wire n_12608;
wire n_7457;
wire n_12383;
wire n_7718;
wire n_10918;
wire n_16556;
wire n_17383;
wire n_18078;
wire n_16629;
wire n_7617;
wire n_13629;
wire n_14671;
wire n_15041;
wire n_16940;
wire n_13360;
wire n_9197;
wire n_17525;
wire n_14265;
wire n_13351;
wire n_6269;
wire n_17450;
wire n_8843;
wire n_11942;
wire n_17316;
wire n_14709;
wire n_5615;
wire n_12057;
wire n_14098;
wire n_15913;
wire n_5902;
wire n_7768;
wire n_13083;
wire n_5479;
wire n_10964;
wire n_13294;
wire n_14143;
wire n_15165;
wire n_13234;
wire n_16020;
wire n_15632;
wire n_7974;
wire n_13896;
wire n_16669;
wire n_16814;
wire n_12902;
wire n_16723;
wire n_9106;
wire n_7357;
wire n_6013;
wire n_5083;
wire n_8247;
wire n_9564;
wire n_6927;
wire n_15257;
wire n_9627;
wire n_7975;
wire n_10864;
wire n_13380;
wire n_6503;
wire n_8172;
wire n_5888;
wire n_17319;
wire n_8941;
wire n_8940;
wire n_9739;
wire n_7310;
wire n_10598;
wire n_12070;
wire n_11835;
wire n_13021;
wire n_15687;
wire n_16031;
wire n_14797;
wire n_16555;
wire n_11444;
wire n_17464;
wire n_17642;
wire n_5698;
wire n_5592;
wire n_7521;
wire n_12430;
wire n_17406;
wire n_7593;
wire n_7716;
wire n_6256;
wire n_13971;
wire n_15798;
wire n_7406;
wire n_7600;
wire n_11353;
wire n_10223;
wire n_17938;
wire n_5870;
wire n_13884;
wire n_9812;
wire n_14905;
wire n_14415;
wire n_16778;
wire n_11823;
wire n_9646;
wire n_5303;
wire n_15594;
wire n_17978;
wire n_13686;
wire n_18328;
wire n_10451;
wire n_10553;
wire n_12718;
wire n_12393;
wire n_10201;
wire n_12249;
wire n_7076;
wire n_16914;
wire n_11814;
wire n_12719;
wire n_8780;
wire n_10215;
wire n_11205;
wire n_9465;
wire n_12932;
wire n_17489;
wire n_14093;
wire n_9928;
wire n_14150;
wire n_8456;
wire n_17410;
wire n_9970;
wire n_13719;
wire n_11138;
wire n_14238;
wire n_5081;
wire n_9894;
wire n_10100;
wire n_10278;
wire n_5124;
wire n_17161;
wire n_10436;
wire n_15425;
wire n_5807;
wire n_5863;
wire n_17500;
wire n_5943;
wire n_17810;
wire n_16553;
wire n_11048;
wire n_15341;
wire n_16203;
wire n_9129;
wire n_14641;
wire n_6982;
wire n_14616;
wire n_14842;
wire n_7286;
wire n_7137;
wire n_12625;
wire n_9957;
wire n_10915;
wire n_13172;
wire n_9558;
wire n_11292;
wire n_14713;
wire n_15642;
wire n_16766;
wire n_18019;
wire n_13167;
wire n_15185;
wire n_11487;
wire n_11753;
wire n_16935;
wire n_7848;
wire n_6727;
wire n_11782;
wire n_8218;
wire n_10689;
wire n_9267;
wire n_12371;
wire n_7539;
wire n_16231;
wire n_8769;
wire n_7229;
wire n_17119;
wire n_10538;
wire n_8514;
wire n_14628;
wire n_14117;
wire n_13487;
wire n_16232;
wire n_5954;
wire n_11865;
wire n_18154;
wire n_8368;
wire n_12258;
wire n_8334;
wire n_12163;
wire n_15605;
wire n_15743;
wire n_9918;
wire n_16500;
wire n_8159;
wire n_6097;
wire n_10773;
wire n_11397;
wire n_8639;
wire n_10621;
wire n_5047;
wire n_11600;
wire n_15506;
wire n_14116;
wire n_12516;
wire n_14342;
wire n_16143;
wire n_18045;
wire n_5346;
wire n_14916;
wire n_5517;
wire n_7125;
wire n_6677;
wire n_7797;
wire n_8216;
wire n_14979;
wire n_13887;
wire n_14740;
wire n_5109;
wire n_6624;
wire n_7121;
wire n_10924;
wire n_15186;
wire n_11844;
wire n_10874;
wire n_7869;
wire n_6466;
wire n_12871;
wire n_18215;
wire n_10942;
wire n_18034;
wire n_12602;
wire n_12295;
wire n_14171;
wire n_13912;
wire n_15307;
wire n_16501;
wire n_15285;
wire n_14830;
wire n_17546;
wire n_9956;
wire n_15134;
wire n_9095;
wire n_9715;
wire n_14975;
wire n_16363;
wire n_6008;
wire n_15048;
wire n_15338;
wire n_15679;
wire n_12198;
wire n_8337;
wire n_11201;
wire n_14141;
wire n_8257;
wire n_11781;
wire n_10292;
wire n_7983;
wire n_11550;
wire n_12077;
wire n_15404;
wire n_7781;
wire n_8125;
wire n_12166;
wire n_12786;
wire n_13467;
wire n_14677;
wire n_5624;
wire n_14860;
wire n_17962;
wire n_16718;
wire n_5714;
wire n_16069;
wire n_17455;
wire n_5806;
wire n_9246;
wire n_13675;
wire n_16304;
wire n_7624;
wire n_10653;
wire n_9683;
wire n_11945;
wire n_12117;
wire n_12110;
wire n_14716;
wire n_12216;
wire n_6221;
wire n_16741;
wire n_18250;
wire n_7160;
wire n_8063;
wire n_9931;
wire n_6805;
wire n_12098;
wire n_15229;
wire n_6185;
wire n_7762;
wire n_13097;
wire n_13749;
wire n_15064;
wire n_8731;
wire n_14334;
wire n_14683;
wire n_15744;
wire n_18044;
wire n_12102;
wire n_13009;
wire n_14373;
wire n_17718;
wire n_18284;
wire n_14325;
wire n_8950;
wire n_16682;
wire n_16075;
wire n_13535;
wire n_14955;
wire n_17481;
wire n_10624;
wire n_15776;
wire n_12802;
wire n_16254;
wire n_13982;
wire n_6568;
wire n_9011;
wire n_9899;
wire n_5358;
wire n_8295;
wire n_16697;
wire n_13668;
wire n_12570;
wire n_15124;
wire n_13577;
wire n_14836;
wire n_13034;
wire n_6004;
wire n_6351;
wire n_7552;
wire n_8059;
wire n_14292;
wire n_8995;
wire n_17521;
wire n_8146;
wire n_11502;
wire n_14583;
wire n_6901;
wire n_8082;
wire n_11965;
wire n_13046;
wire n_11997;
wire n_16661;
wire n_9094;
wire n_5580;
wire n_5937;
wire n_14589;
wire n_7183;
wire n_13300;
wire n_16693;
wire n_18006;
wire n_12456;
wire n_11424;
wire n_6411;
wire n_15617;
wire n_18082;
wire n_8339;
wire n_15898;
wire n_13405;
wire n_11816;
wire n_9195;
wire n_7746;
wire n_13641;
wire n_5435;
wire n_12768;
wire n_10867;
wire n_11361;
wire n_10701;
wire n_14735;
wire n_14233;
wire n_15848;
wire n_11062;
wire n_14068;
wire n_18131;
wire n_6873;
wire n_14610;
wire n_15253;
wire n_14584;
wire n_17321;
wire n_10741;
wire n_5373;
wire n_5745;
wire n_15223;
wire n_8032;
wire n_16607;
wire n_14505;
wire n_7139;
wire n_14655;
wire n_12710;
wire n_12483;
wire n_8640;
wire n_9332;
wire n_16947;
wire n_10016;
wire n_16019;
wire n_10070;
wire n_5279;
wire n_14121;
wire n_17246;
wire n_8351;
wire n_10190;
wire n_17432;
wire n_14673;
wire n_11499;
wire n_8196;
wire n_11580;
wire n_16753;
wire n_15084;
wire n_12128;
wire n_6594;
wire n_5493;
wire n_17604;
wire n_7857;
wire n_9054;
wire n_10812;
wire n_10150;
wire n_15132;
wire n_9460;
wire n_17011;
wire n_17328;
wire n_17184;
wire n_9638;
wire n_17600;
wire n_12682;
wire n_13028;
wire n_14896;
wire n_6387;
wire n_13613;
wire n_12389;
wire n_16531;
wire n_7223;
wire n_7890;
wire n_16902;
wire n_12464;
wire n_6179;
wire n_9281;
wire n_7338;
wire n_5321;
wire n_10134;
wire n_11379;
wire n_13700;
wire n_7964;
wire n_13135;
wire n_5096;
wire n_9740;
wire n_16024;
wire n_9475;
wire n_8865;
wire n_9661;
wire n_13721;
wire n_13056;
wire n_10861;
wire n_6019;
wire n_12313;
wire n_15672;
wire n_17575;
wire n_17469;
wire n_12147;
wire n_11070;
wire n_9190;
wire n_7165;
wire n_8110;
wire n_6222;
wire n_11245;
wire n_17290;
wire n_10635;
wire n_12874;
wire n_14749;
wire n_8475;
wire n_8838;
wire n_6223;
wire n_6435;
wire n_12909;
wire n_9143;
wire n_14871;
wire n_12990;
wire n_17813;
wire n_7235;
wire n_5210;
wire n_16805;
wire n_6976;
wire n_6486;
wire n_8488;
wire n_15547;
wire n_11286;
wire n_16095;
wire n_5657;
wire n_16685;
wire n_6889;
wire n_8766;
wire n_6083;
wire n_15785;
wire n_17363;
wire n_6844;
wire n_13628;
wire n_7795;
wire n_8969;
wire n_12240;
wire n_11631;
wire n_7404;
wire n_13326;
wire n_9891;
wire n_10555;
wire n_6295;
wire n_11147;
wire n_10897;
wire n_9087;
wire n_11700;
wire n_15894;
wire n_15151;
wire n_9804;
wire n_16392;
wire n_10287;
wire n_8087;
wire n_8119;
wire n_15793;
wire n_15227;
wire n_10135;
wire n_9321;
wire n_7885;
wire n_12468;
wire n_18130;
wire n_5857;
wire n_10983;
wire n_15243;
wire n_16204;
wire n_8173;
wire n_11833;
wire n_9800;
wire n_7437;
wire n_15242;
wire n_17055;
wire n_11053;
wire n_8420;
wire n_6241;
wire n_15283;
wire n_6087;
wire n_14035;
wire n_17675;
wire n_8019;
wire n_9186;
wire n_15266;
wire n_15327;
wire n_13307;
wire n_9951;
wire n_6846;
wire n_11335;
wire n_9243;
wire n_14346;
wire n_14921;
wire n_13509;
wire n_14902;
wire n_17036;
wire n_16349;
wire n_15416;
wire n_5756;
wire n_12294;
wire n_11336;
wire n_11247;
wire n_11057;
wire n_7822;
wire n_6041;
wire n_12186;
wire n_15943;
wire n_8851;
wire n_14949;
wire n_6994;
wire n_15069;
wire n_10987;
wire n_15523;
wire n_17931;
wire n_7449;
wire n_11262;
wire n_7329;
wire n_9359;
wire n_5708;
wire n_10402;
wire n_15083;
wire n_15599;
wire n_13238;
wire n_8687;
wire n_6790;
wire n_14813;
wire n_15280;
wire n_12860;
wire n_15357;
wire n_10001;
wire n_13598;
wire n_15801;
wire n_10666;
wire n_17054;
wire n_7194;
wire n_11363;
wire n_6273;
wire n_14482;
wire n_17825;
wire n_11783;
wire n_16451;
wire n_8740;
wire n_11661;
wire n_14450;
wire n_15664;
wire n_11026;
wire n_11889;
wire n_6807;
wire n_15066;
wire n_14990;
wire n_14806;
wire n_5927;
wire n_15433;
wire n_16581;
wire n_10189;
wire n_17091;
wire n_12939;
wire n_16795;
wire n_9879;
wire n_17206;
wire n_18132;
wire n_17114;
wire n_8221;
wire n_8468;
wire n_7708;
wire n_7696;
wire n_14708;
wire n_11756;
wire n_18137;
wire n_13153;
wire n_11419;
wire n_11232;
wire n_13211;
wire n_15570;
wire n_17630;
wire n_5638;
wire n_9975;
wire n_10997;
wire n_7115;
wire n_16494;
wire n_9335;
wire n_13763;
wire n_18251;
wire n_5670;
wire n_9171;
wire n_12778;
wire n_17004;
wire n_8815;
wire n_18102;
wire n_14994;
wire n_17034;
wire n_18244;
wire n_9942;
wire n_11081;
wire n_13304;
wire n_12813;
wire n_13711;
wire n_13391;
wire n_11407;
wire n_17381;
wire n_5584;
wire n_8952;
wire n_14102;
wire n_11654;
wire n_9247;
wire n_9933;
wire n_5965;
wire n_12907;
wire n_16863;
wire n_7958;
wire n_10209;
wire n_18174;
wire n_17750;
wire n_8128;
wire n_11519;
wire n_17770;
wire n_18148;
wire n_16368;
wire n_17327;
wire n_5751;
wire n_13475;
wire n_17071;
wire n_10434;
wire n_5664;
wire n_12011;
wire n_9441;
wire n_11668;
wire n_11913;
wire n_11978;
wire n_15013;
wire n_15718;
wire n_15014;
wire n_10829;
wire n_5641;
wire n_8667;
wire n_6218;
wire n_8863;
wire n_7281;
wire n_10233;
wire n_11810;
wire n_8106;
wire n_9362;
wire n_16323;
wire n_15710;
wire n_10690;
wire n_15723;
wire n_14212;
wire n_10311;
wire n_15639;
wire n_16286;
wire n_14001;
wire n_6824;
wire n_11198;
wire n_11767;
wire n_8717;
wire n_14712;
wire n_6189;
wire n_11595;
wire n_18188;
wire n_16201;
wire n_16857;
wire n_13305;
wire n_9216;
wire n_11168;
wire n_8299;
wire n_5262;
wire n_9200;
wire n_16483;
wire n_6993;
wire n_6037;
wire n_7245;
wire n_11872;
wire n_13787;
wire n_16187;
wire n_18204;
wire n_5963;
wire n_5980;
wire n_8892;
wire n_15303;
wire n_11235;
wire n_12007;
wire n_18070;
wire n_18257;
wire n_10146;
wire n_14445;
wire n_14550;
wire n_9067;
wire n_16776;
wire n_18120;
wire n_12712;
wire n_5310;
wire n_9152;
wire n_12846;
wire n_8287;
wire n_11906;
wire n_13837;
wire n_18166;
wire n_16374;
wire n_17974;
wire n_15139;
wire n_14604;
wire n_16827;
wire n_6153;
wire n_16769;
wire n_15604;
wire n_9074;
wire n_13550;
wire n_7989;
wire n_14528;
wire n_13908;
wire n_15019;
wire n_10790;
wire n_16241;
wire n_5970;
wire n_6418;
wire n_12908;
wire n_6564;
wire n_13461;
wire n_13955;
wire n_15997;
wire n_8657;
wire n_12505;
wire n_12747;
wire n_15150;
wire n_12577;
wire n_12426;
wire n_17069;
wire n_16175;
wire n_5146;
wire n_11122;
wire n_9287;
wire n_18055;
wire n_8197;
wire n_16892;
wire n_9511;
wire n_17279;
wire n_14500;
wire n_13733;
wire n_15621;
wire n_10052;
wire n_16600;
wire n_13067;
wire n_8081;
wire n_7192;
wire n_12309;
wire n_13974;
wire n_15158;
wire n_6671;
wire n_10407;
wire n_10449;
wire n_11324;
wire n_12164;
wire n_15803;
wire n_6591;
wire n_6266;
wire n_10950;
wire n_14235;
wire n_14425;
wire n_7161;
wire n_11566;
wire n_17403;
wire n_14352;
wire n_7580;
wire n_7153;
wire n_9880;
wire n_17944;
wire n_10072;
wire n_14929;
wire n_9843;
wire n_5213;
wire n_8609;
wire n_17568;
wire n_16913;
wire n_11869;
wire n_14609;
wire n_15640;
wire n_5441;
wire n_6517;
wire n_14326;
wire n_11579;
wire n_17248;
wire n_14196;
wire n_8559;
wire n_7350;
wire n_15938;
wire n_10838;
wire n_5690;
wire n_12140;
wire n_13312;
wire n_10369;
wire n_14075;
wire n_16366;
wire n_6967;
wire n_5885;
wire n_10920;
wire n_9248;
wire n_17237;
wire n_6433;
wire n_10321;
wire n_12178;
wire n_7535;
wire n_6893;
wire n_9128;
wire n_13003;
wire n_16626;
wire n_8452;
wire n_14261;
wire n_17368;
wire n_10506;
wire n_5461;
wire n_11082;
wire n_7178;
wire n_13192;
wire n_7480;
wire n_10224;
wire n_16333;
wire n_7632;
wire n_12554;
wire n_16608;
wire n_10671;
wire n_8771;
wire n_15212;
wire n_8140;
wire n_9528;
wire n_8476;
wire n_17693;
wire n_18028;
wire n_13213;
wire n_12912;
wire n_6501;
wire n_8981;
wire n_10157;
wire n_12200;
wire n_16803;
wire n_11529;
wire n_9507;
wire n_6028;
wire n_17301;
wire n_14603;
wire n_16389;
wire n_13557;
wire n_16001;
wire n_14332;
wire n_5629;
wire n_9533;
wire n_5634;
wire n_5430;
wire n_13890;
wire n_12611;
wire n_13767;
wire n_5362;
wire n_8137;
wire n_6709;
wire n_15630;
wire n_14285;
wire n_17275;
wire n_15924;
wire n_14443;
wire n_12322;
wire n_8469;
wire n_13270;
wire n_10808;
wire n_6798;
wire n_12303;
wire n_16901;
wire n_12507;
wire n_5702;
wire n_5050;
wire n_16023;
wire n_5063;
wire n_15941;
wire n_17801;
wire n_5229;
wire n_7844;
wire n_5199;
wire n_11430;
wire n_11882;
wire n_12023;
wire n_14379;
wire n_13802;
wire n_14128;
wire n_14991;
wire n_16754;
wire n_9665;
wire n_12171;
wire n_8423;
wire n_13476;
wire n_12395;
wire n_12472;
wire n_12815;
wire n_5527;
wire n_6986;
wire n_11146;
wire n_8090;
wire n_5609;
wire n_12239;
wire n_5416;
wire n_10504;
wire n_11279;
wire n_15715;
wire n_10975;
wire n_13176;
wire n_5266;
wire n_7471;
wire n_13443;
wire n_17024;
wire n_18268;
wire n_13418;
wire n_9436;
wire n_16434;
wire n_17540;
wire n_5355;
wire n_18068;
wire n_17913;
wire n_9562;
wire n_6745;
wire n_18163;
wire n_11516;
wire n_11005;
wire n_16659;
wire n_8260;
wire n_8481;
wire n_13961;
wire n_15342;
wire n_5977;
wire n_15261;
wire n_6811;
wire n_15867;
wire n_14811;
wire n_6209;
wire n_6875;
wire n_13799;
wire n_10566;
wire n_15369;
wire n_17755;
wire n_15745;
wire n_15491;
wire n_14685;
wire n_16215;
wire n_11451;
wire n_16969;
wire n_14146;
wire n_17891;
wire n_15870;
wire n_15763;
wire n_11980;
wire n_11076;
wire n_17105;
wire n_7905;
wire n_14877;
wire n_6853;
wire n_12121;
wire n_15020;
wire n_5551;
wire n_7766;
wire n_7594;
wire n_7803;
wire n_7340;
wire n_10837;
wire n_6699;
wire n_7747;
wire n_15648;
wire n_6073;
wire n_17409;
wire n_8205;
wire n_5767;
wire n_8401;
wire n_6324;
wire n_12116;
wire n_8651;
wire n_18124;
wire n_14260;
wire n_5640;
wire n_10199;
wire n_13020;
wire n_13621;
wire n_8284;
wire n_10688;
wire n_14999;
wire n_12261;
wire n_9255;
wire n_16189;
wire n_15873;
wire n_18003;
wire n_10039;
wire n_15625;
wire n_8828;
wire n_5655;
wire n_5475;
wire n_11239;
wire n_12338;
wire n_12259;
wire n_14310;
wire n_17080;
wire n_17995;
wire n_14608;
wire n_7603;
wire n_6138;
wire n_8510;
wire n_8810;
wire n_13163;
wire n_16825;
wire n_9034;
wire n_15611;
wire n_15778;
wire n_17437;
wire n_9203;
wire n_9601;
wire n_13173;
wire n_5692;
wire n_10443;
wire n_7726;
wire n_11623;
wire n_12825;
wire n_16923;
wire n_17532;
wire n_18091;
wire n_7494;
wire n_5921;
wire n_12222;
wire n_8024;
wire n_9946;
wire n_14383;
wire n_5168;
wire n_10887;
wire n_13253;
wire n_13119;
wire n_9967;
wire n_6477;
wire n_16492;
wire n_10735;
wire n_10274;
wire n_16621;
wire n_8739;
wire n_8373;
wire n_8133;
wire n_8919;
wire n_14469;
wire n_11740;
wire n_17697;
wire n_13525;
wire n_17624;
wire n_10482;
wire n_15478;
wire n_6159;
wire n_11012;
wire n_17154;
wire n_9647;
wire n_16197;
wire n_6283;
wire n_7396;
wire n_9912;
wire n_14237;
wire n_16617;
wire n_16649;
wire n_17103;
wire n_17694;
wire n_17397;
wire n_16292;
wire n_16775;
wire n_5322;
wire n_14774;
wire n_16884;
wire n_11698;
wire n_7116;
wire n_12779;
wire n_14782;
wire n_16018;
wire n_14694;
wire n_7519;
wire n_10485;
wire n_16879;
wire n_17365;
wire n_6943;
wire n_9329;
wire n_17549;
wire n_6827;
wire n_10652;
wire n_12465;
wire n_8318;
wire n_6173;
wire n_13042;
wire n_16170;
wire n_8542;
wire n_17007;
wire n_11059;
wire n_17652;
wire n_14592;
wire n_8543;
wire n_8846;
wire n_10791;
wire n_17293;
wire n_6312;
wire n_14803;
wire n_14895;
wire n_11236;
wire n_13514;
wire n_14183;
wire n_12852;
wire n_13994;
wire n_5371;
wire n_17068;
wire n_12334;
wire n_15502;
wire n_13162;
wire n_17553;
wire n_6997;
wire n_15044;
wire n_5418;
wire n_15095;
wire n_15910;
wire n_11196;
wire n_11629;
wire n_10411;
wire n_12847;
wire n_7770;
wire n_16037;
wire n_10286;
wire n_12511;
wire n_11643;
wire n_17751;
wire n_18000;
wire n_16868;
wire n_16939;
wire n_7664;
wire n_10913;
wire n_13199;
wire n_15068;
wire n_5316;
wire n_9890;
wire n_13969;
wire n_14736;
wire n_10273;
wire n_15005;
wire n_6300;
wire n_9609;
wire n_9883;
wire n_10172;
wire n_16642;
wire n_7815;
wire n_16011;
wire n_13209;
wire n_12014;
wire n_9046;
wire n_13407;
wire n_9361;
wire n_8163;
wire n_13980;
wire n_11609;
wire n_17534;
wire n_6131;
wire n_17053;
wire n_16853;
wire n_15554;
wire n_10806;
wire n_6537;
wire n_13712;
wire n_5933;
wire n_13059;
wire n_15759;
wire n_12305;
wire n_17152;
wire n_14864;
wire n_13681;
wire n_9864;
wire n_13521;
wire n_18101;
wire n_12485;
wire n_12408;
wire n_7023;
wire n_8972;
wire n_9300;
wire n_15749;
wire n_13263;
wire n_17153;
wire n_17555;
wire n_12238;
wire n_16271;
wire n_16373;
wire n_7428;
wire n_5112;
wire n_10694;
wire n_5386;
wire n_11509;
wire n_6783;
wire n_11351;
wire n_17797;
wire n_9353;
wire n_9766;
wire n_7465;
wire n_13720;
wire n_16673;
wire n_11271;
wire n_8293;
wire n_9832;
wire n_14421;
wire n_16213;
wire n_10754;
wire n_14480;
wire n_14663;
wire n_12409;
wire n_13565;
wire n_17542;
wire n_11307;
wire n_13685;
wire n_5123;
wire n_9954;
wire n_8737;
wire n_13129;
wire n_14091;
wire n_7961;
wire n_10953;
wire n_15477;
wire n_11761;
wire n_7847;
wire n_9997;
wire n_10703;
wire n_16048;
wire n_17606;
wire n_11973;
wire n_15144;
wire n_9334;
wire n_7149;
wire n_8252;
wire n_15052;
wire n_6459;
wire n_9622;
wire n_10847;
wire n_11565;
wire n_14088;
wire n_13446;
wire n_17169;
wire n_16387;
wire n_11252;
wire n_16569;
wire n_15786;
wire n_8450;
wire n_7700;
wire n_9284;
wire n_16964;
wire n_16257;
wire n_16394;
wire n_5644;
wire n_14318;
wire n_13865;
wire n_16432;
wire n_9147;
wire n_16720;
wire n_8367;
wire n_12454;
wire n_10103;
wire n_8834;
wire n_6869;
wire n_8078;
wire n_10922;
wire n_16713;
wire n_10413;
wire n_11571;
wire n_16647;
wire n_16793;
wire n_10738;
wire n_13197;
wire n_12587;
wire n_17861;
wire n_5424;
wire n_15222;
wire n_7914;
wire n_17052;
wire n_17922;
wire n_13916;
wire n_10995;
wire n_17443;
wire n_7967;
wire n_9794;
wire n_11858;
wire n_14812;
wire n_13963;
wire n_17847;
wire n_7117;
wire n_14845;
wire n_9354;
wire n_8471;
wire n_11904;
wire n_15890;
wire n_12324;
wire n_13925;
wire n_17189;
wire n_12130;
wire n_17262;
wire n_18179;
wire n_6977;
wire n_8474;
wire n_12643;
wire n_7984;
wire n_16397;
wire n_16789;
wire n_13448;
wire n_15931;
wire n_10185;
wire n_11131;
wire n_17226;
wire n_17820;
wire n_11478;
wire n_10591;
wire n_11656;
wire n_14426;
wire n_16228;
wire n_12955;
wire n_16565;
wire n_11673;
wire n_11821;
wire n_8361;
wire n_15412;
wire n_17285;
wire n_18266;
wire n_6313;
wire n_16378;
wire n_14348;
wire n_11701;
wire n_10856;
wire n_16337;
wire n_15757;
wire n_13626;
wire n_18276;
wire n_6569;
wire n_18216;
wire n_17792;
wire n_15356;
wire n_16916;
wire n_17629;
wire n_9494;
wire n_16132;
wire n_6555;
wire n_9614;
wire n_11283;
wire n_13616;
wire n_16745;
wire n_16729;
wire n_17551;
wire n_12948;
wire n_16589;
wire n_14329;
wire n_9551;
wire n_13653;
wire n_6639;
wire n_7516;
wire n_15552;
wire n_5496;
wire n_13694;
wire n_9154;
wire n_13233;
wire n_10677;
wire n_7596;
wire n_13189;
wire n_16089;
wire n_13640;
wire n_5864;
wire n_6536;
wire n_14211;
wire n_8553;
wire n_6490;
wire n_8301;
wire n_15003;
wire n_10610;
wire n_6961;
wire n_13392;
wire n_12574;
wire n_12697;
wire n_9437;
wire n_16871;
wire n_18150;
wire n_5460;
wire n_7628;
wire n_9276;
wire n_6761;
wire n_15760;
wire n_14572;
wire n_9346;
wire n_11229;
wire n_15626;
wire n_5333;
wire n_15724;
wire n_6294;
wire n_14851;
wire n_11636;
wire n_6767;
wire n_8518;
wire n_7427;
wire n_6802;
wire n_7527;
wire n_13962;
wire n_17486;
wire n_12162;
wire n_5570;
wire n_9514;
wire n_6326;
wire n_18206;
wire n_11919;
wire n_9402;
wire n_14118;
wire n_10456;
wire n_12634;
wire n_11675;
wire n_10343;
wire n_17236;
wire n_7838;
wire n_8364;
wire n_7786;
wire n_5983;
wire n_9580;
wire n_14134;
wire n_9005;
wire n_5804;
wire n_12236;
wire n_7979;
wire n_6376;
wire n_8621;
wire n_6167;
wire n_15231;
wire n_8993;
wire n_7926;
wire n_7411;
wire n_5910;
wire n_12632;
wire n_7101;
wire n_12398;
wire n_14545;
wire n_17779;
wire n_5040;
wire n_6730;
wire n_6948;
wire n_15415;
wire n_10979;
wire n_13591;
wire n_10487;
wire n_10332;
wire n_16491;
wire n_9162;
wire n_16861;
wire n_18265;
wire n_9921;
wire n_9443;
wire n_6582;
wire n_13479;
wire n_8910;
wire n_7752;
wire n_13631;
wire n_15453;
wire n_9897;
wire n_11570;
wire n_15364;
wire n_10807;
wire n_6996;
wire n_11855;
wire n_9817;
wire n_14930;
wire n_15389;
wire n_11667;
wire n_15166;
wire n_9301;
wire n_17573;
wire n_6974;
wire n_7731;
wire n_8753;
wire n_15265;
wire n_6765;
wire n_7577;
wire n_8388;
wire n_9401;
wire n_16171;
wire n_16701;
wire n_8321;
wire n_6921;
wire n_11290;
wire n_13738;
wire n_15739;
wire n_8044;
wire n_15937;
wire n_8091;
wire n_14137;
wire n_16502;
wire n_8486;
wire n_7845;
wire n_13122;
wire n_10750;
wire n_17259;
wire n_12292;
wire n_7709;
wire n_9689;
wire n_15628;
wire n_11592;
wire n_11466;
wire n_5194;
wire n_15536;
wire n_13346;
wire n_9982;
wire n_6898;
wire n_12056;
wire n_6710;
wire n_13149;
wire n_5717;
wire n_7162;
wire n_6565;
wire n_5464;
wire n_8508;
wire n_12679;
wire n_8261;
wire n_14179;
wire n_15262;
wire n_12811;
wire n_18230;
wire n_18059;
wire n_13100;
wire n_14821;
wire n_5886;
wire n_7080;
wire n_16096;
wire n_9886;
wire n_7744;
wire n_13232;
wire n_17340;
wire n_12897;
wire n_8034;
wire n_8841;
wire n_17179;
wire n_17447;
wire n_10970;
wire n_14401;
wire n_7302;
wire n_6533;
wire n_12837;
wire n_18286;
wire n_17193;
wire n_10264;
wire n_6960;
wire n_8201;
wire n_6426;
wire n_6634;
wire n_7180;
wire n_6836;
wire n_5239;
wire n_5610;
wire n_11983;
wire n_13840;
wire n_15735;
wire n_12605;
wire n_11043;
wire n_8947;
wire n_5197;
wire n_15792;
wire n_16233;
wire n_9671;
wire n_6972;
wire n_9297;
wire n_8788;
wire n_10472;
wire n_13460;
wire n_13389;
wire n_7111;
wire n_7549;
wire n_14180;
wire n_16978;
wire n_5785;
wire n_11415;
wire n_15849;
wire n_17928;
wire n_13578;
wire n_6344;
wire n_14773;
wire n_5305;
wire n_5994;
wire n_6093;
wire n_10499;
wire n_8093;
wire n_11680;
wire n_13870;
wire n_15096;
wire n_6010;
wire n_14958;
wire n_15791;
wire n_15696;
wire n_7247;
wire n_13088;
wire n_11446;
wire n_9225;
wire n_8061;
wire n_6833;
wire n_11972;
wire n_14247;
wire n_5376;
wire n_13862;
wire n_16674;
wire n_13600;
wire n_17556;
wire n_11103;
wire n_7481;
wire n_10435;
wire n_12220;
wire n_13843;
wire n_10066;
wire n_13605;
wire n_14707;
wire n_5204;
wire n_17177;
wire n_7292;
wire n_10341;
wire n_12230;
wire n_15987;
wire n_14511;
wire n_8811;
wire n_12995;
wire n_7150;
wire n_13486;
wire n_14176;
wire n_17574;
wire n_7687;
wire n_10184;
wire n_10498;
wire n_13599;
wire n_16936;
wire n_12867;
wire n_18229;
wire n_8507;
wire n_9662;
wire n_10508;
wire n_9057;
wire n_12497;
wire n_14173;
wire n_14323;
wire n_16610;
wire n_14667;
wire n_12406;
wire n_6265;
wire n_8861;
wire n_14544;
wire n_18026;
wire n_11749;
wire n_14875;
wire n_6821;
wire n_8661;
wire n_15740;
wire n_11417;
wire n_18312;
wire n_8545;
wire n_12725;
wire n_6373;
wire n_6988;
wire n_8755;
wire n_5788;
wire n_11490;
wire n_12401;
wire n_13404;
wire n_8573;
wire n_8191;
wire n_11704;
wire n_16534;
wire n_7692;
wire n_5897;
wire n_6887;
wire n_11343;
wire n_10865;
wire n_14777;
wire n_16984;
wire n_15065;
wire n_9809;
wire n_13277;
wire n_12185;
wire n_16041;
wire n_13518;
wire n_14157;
wire n_17782;
wire n_8683;
wire n_17983;
wire n_15293;
wire n_10081;
wire n_8836;
wire n_6676;
wire n_7016;
wire n_6347;
wire n_6492;
wire n_13540;
wire n_14366;
wire n_12161;
wire n_15756;
wire n_15676;
wire n_16750;
wire n_9448;
wire n_16220;
wire n_17919;
wire n_8446;
wire n_8136;
wire n_9799;
wire n_7742;
wire n_10577;
wire n_9313;
wire n_15085;
wire n_8916;
wire n_14650;
wire n_14657;
wire n_7955;
wire n_5795;
wire n_17566;
wire n_7072;
wire n_5508;
wire n_10037;
wire n_17743;
wire n_13370;
wire n_12424;
wire n_5582;
wire n_16385;
wire n_15844;
wire n_10234;
wire n_14801;
wire n_7374;
wire n_7440;
wire n_9989;
wire n_11766;
wire n_7758;
wire n_11639;
wire n_17491;
wire n_7547;
wire n_14802;
wire n_12114;
wire n_13171;
wire n_11967;
wire n_9438;
wire n_13528;
wire n_7201;
wire n_13419;
wire n_17621;
wire n_14087;
wire n_16277;
wire n_11457;
wire n_10832;
wire n_12490;
wire n_10036;
wire n_12571;
wire n_11932;
wire n_15053;
wire n_5746;
wire n_15559;
wire n_17561;
wire n_5292;
wire n_14656;
wire n_10853;
wire n_12508;
wire n_12582;
wire n_6648;
wire n_7880;
wire n_12052;
wire n_14757;
wire n_8075;
wire n_13937;
wire n_14298;
wire n_14623;
wire n_8857;
wire n_11275;
wire n_14253;
wire n_8587;
wire n_12337;
wire n_9675;
wire n_10030;
wire n_17215;
wire n_5630;
wire n_9667;
wire n_10676;
wire n_11819;
wire n_8071;
wire n_13159;
wire n_17929;
wire n_15766;
wire n_10815;
wire n_12928;
wire n_16064;
wire n_17266;
wire n_17221;
wire n_11589;
wire n_11309;
wire n_17496;
wire n_12927;
wire n_15161;
wire n_15401;
wire n_13347;
wire n_11803;
wire n_16690;
wire n_7513;
wire n_11067;
wire n_12321;
wire n_17227;
wire n_11274;
wire n_5264;
wire n_9537;
wire n_10833;
wire n_7413;
wire n_11174;
wire n_11770;
wire n_11795;
wire n_7540;
wire n_8646;
wire n_15381;
wire n_15829;
wire n_9866;
wire n_5504;
wire n_8630;
wire n_7622;
wire n_9602;
wire n_14392;
wire n_15373;
wire n_7005;
wire n_11266;
wire n_11151;
wire n_7353;
wire n_6219;
wire n_10071;
wire n_9885;
wire n_15216;
wire n_14115;
wire n_12592;
wire n_15654;
wire n_14992;
wire n_15811;
wire n_12698;
wire n_13343;
wire n_17980;
wire n_8315;
wire n_14282;
wire n_6965;
wire n_9260;
wire n_13938;
wire n_16063;
wire n_8314;
wire n_12048;
wire n_6720;
wire n_14615;
wire n_8149;
wire n_16279;
wire n_16169;
wire n_6032;
wire n_11413;
wire n_8581;
wire n_16654;
wire n_15729;
wire n_13932;
wire n_13094;
wire n_7174;
wire n_8565;
wire n_6205;
wire n_6362;
wire n_6402;
wire n_14668;
wire n_14509;
wire n_7166;
wire n_5060;
wire n_15495;
wire n_17250;
wire n_7607;
wire n_8209;
wire n_9159;
wire n_5334;
wire n_15973;
wire n_16784;
wire n_16309;
wire n_15317;
wire n_7816;
wire n_13290;
wire n_9654;
wire n_8560;
wire n_7591;
wire n_15500;
wire n_17039;
wire n_8141;
wire n_5775;
wire n_14139;
wire n_7830;
wire n_7282;
wire n_6491;
wire n_13198;
wire n_8302;
wire n_10015;
wire n_17892;
wire n_17900;
wire n_9306;
wire n_7151;
wire n_11652;
wire n_11682;
wire n_16453;
wire n_12801;
wire n_6229;
wire n_17986;
wire n_11091;
wire n_15325;
wire n_11929;
wire n_9978;
wire n_17863;
wire n_16116;
wire n_5731;
wire n_8612;
wire n_5581;
wire n_17954;
wire n_18308;
wire n_7446;
wire n_16139;
wire n_6668;
wire n_10362;
wire n_16921;
wire n_15952;
wire n_7053;
wire n_8724;
wire n_11331;
wire n_11640;
wire n_14702;
wire n_16288;
wire n_5831;
wire n_10171;
wire n_12552;
wire n_7473;
wire n_10183;
wire n_10471;
wire n_14674;
wire n_8070;
wire n_6835;
wire n_13039;
wire n_6419;
wire n_18224;
wire n_6039;
wire n_12704;
wire n_11237;
wire n_15304;
wire n_11601;
wire n_11741;
wire n_14130;
wire n_14402;
wire n_15839;
wire n_14305;
wire n_5884;
wire n_14400;
wire n_17924;
wire n_17492;
wire n_9279;
wire n_8457;
wire n_8922;
wire n_5653;
wire n_10095;
wire n_8248;
wire n_7966;
wire n_9509;
wire n_6258;
wire n_10549;
wire n_7070;
wire n_5394;
wire n_15775;
wire n_17382;
wire n_11721;
wire n_17828;
wire n_6755;
wire n_16601;
wire n_9563;
wire n_7276;
wire n_7351;
wire n_12256;
wire n_7942;
wire n_10057;
wire n_12477;
wire n_12245;
wire n_11093;
wire n_12184;
wire n_6084;
wire n_10301;
wire n_15888;
wire n_16777;
wire n_9496;
wire n_13156;
wire n_15531;
wire n_8411;
wire n_12657;
wire n_12740;
wire n_9644;
wire n_7412;
wire n_7157;
wire n_6436;
wire n_7666;
wire n_12089;
wire n_13957;
wire n_6472;
wire n_14051;
wire n_5421;
wire n_8527;
wire n_11097;
wire n_7211;
wire n_10394;
wire n_10154;
wire n_11681;
wire n_6531;
wire n_5309;
wire n_7901;
wire n_8689;
wire n_11522;
wire n_14724;
wire n_17158;
wire n_9750;
wire n_18201;
wire n_9980;
wire n_13164;
wire n_16476;
wire n_10818;
wire n_12145;
wire n_17271;
wire n_16888;
wire n_8988;
wire n_11105;
wire n_12647;
wire n_12377;
wire n_12721;
wire n_9251;
wire n_10141;
wire n_15906;
wire n_7368;
wire n_16398;
wire n_16681;
wire n_16839;
wire n_17691;
wire n_15420;
wire n_13624;
wire n_8549;
wire n_12541;
wire n_12316;
wire n_6567;
wire n_5889;
wire n_11849;
wire n_6771;
wire n_11578;
wire n_13484;
wire n_10916;
wire n_10208;
wire n_13714;
wire n_6389;
wire n_10182;
wire n_13655;
wire n_9616;
wire n_15142;
wire n_15037;
wire n_12399;
wire n_15189;
wire n_8004;
wire n_10929;
wire n_8658;
wire n_16609;
wire n_16785;
wire n_9959;
wire n_8375;
wire n_10403;
wire n_17495;
wire n_5764;
wire n_10260;
wire n_6910;
wire n_5428;
wire n_9291;
wire n_9092;
wire n_10261;
wire n_6442;
wire n_12285;
wire n_16725;
wire n_16180;
wire n_16870;
wire n_17737;
wire n_13606;
wire n_6102;
wire n_18311;
wire n_16473;
wire n_8908;
wire n_5541;
wire n_15067;
wire n_13438;
wire n_16003;
wire n_10384;
wire n_6441;
wire n_15868;
wire n_5543;
wire n_10372;
wire n_9818;
wire n_10237;
wire n_9283;
wire n_5678;
wire n_5935;
wire n_11219;
wire n_13498;
wire n_14453;
wire n_16842;
wire n_17048;
wire n_17960;
wire n_7677;
wire n_5085;
wire n_8569;
wire n_16886;
wire n_13661;
wire n_17925;
wire n_10118;
wire n_8676;
wire n_5950;
wire n_16593;
wire n_17029;
wire n_15260;
wire n_12379;
wire n_15413;
wire n_17819;
wire n_13496;
wire n_7929;
wire n_10028;
wire n_12257;
wire n_10691;
wire n_17089;
wire n_8399;
wire n_5995;
wire n_12246;
wire n_16060;
wire n_18285;
wire n_16864;
wire n_15363;
wire n_11069;
wire n_6162;
wire n_5116;
wire n_6331;
wire n_13674;
wire n_14099;
wire n_6006;
wire n_16582;
wire n_8421;
wire n_6109;
wire n_17746;
wire n_11268;
wire n_6278;
wire n_9304;
wire n_12655;
wire n_13818;
wire n_14855;
wire n_6787;
wire n_10777;
wire n_11066;
wire n_6872;
wire n_6208;
wire n_14642;
wire n_15858;
wire n_6632;
wire n_13133;
wire n_9310;
wire n_18200;
wire n_7754;
wire n_5411;
wire n_14246;
wire n_9830;
wire n_17332;
wire n_9913;
wire n_11728;
wire n_7027;
wire n_8001;
wire n_5671;
wire n_8322;
wire n_12272;
wire n_6990;
wire n_12862;
wire n_16563;
wire n_8403;
wire n_6349;
wire n_14885;
wire n_13140;
wire n_17008;
wire n_11796;
wire n_18092;
wire n_13573;
wire n_7631;
wire n_16625;
wire n_17444;
wire n_6830;
wire n_8999;
wire n_12662;
wire n_8754;
wire n_5185;
wire n_7939;
wire n_17676;
wire n_8675;
wire n_7898;
wire n_10715;
wire n_12136;
wire n_14889;
wire n_16770;
wire n_9375;
wire n_6359;
wire n_15111;
wire n_16068;
wire n_8596;
wire n_10665;
wire n_10073;
wire n_10291;
wire n_13251;
wire n_14890;
wire n_8858;
wire n_8666;
wire n_11873;
wire n_17963;
wire n_15579;
wire n_8313;
wire n_7763;
wire n_10296;
wire n_13154;
wire n_7498;
wire n_17831;
wire n_5076;
wire n_7377;
wire n_17739;
wire n_11228;
wire n_8555;
wire n_5379;
wire n_15149;
wire n_16458;
wire n_15769;
wire n_17771;
wire n_12517;
wire n_13796;
wire n_16308;
wire n_18168;
wire n_16173;
wire n_16875;
wire n_6301;
wire n_17688;
wire n_12031;
wire n_11743;
wire n_14274;
wire n_10512;
wire n_8610;
wire n_13195;
wire n_13314;
wire n_14456;
wire n_13679;
wire n_16648;
wire n_17419;
wire n_12993;
wire n_10324;
wire n_16402;
wire n_13658;
wire n_12663;
wire n_7945;
wire n_5945;
wire n_14850;
wire n_11261;
wire n_13667;
wire n_9323;
wire n_17623;
wire n_6744;
wire n_10765;
wire n_9985;
wire n_12039;
wire n_17344;
wire n_11023;
wire n_17473;
wire n_8615;
wire n_11382;
wire n_5811;
wire n_6439;
wire n_14278;
wire n_10026;
wire n_8677;
wire n_9355;
wire n_17286;
wire n_8602;
wire n_9714;
wire n_12938;
wire n_7381;
wire n_13772;
wire n_16348;
wire n_10041;
wire n_5565;
wire n_7948;
wire n_16210;
wire n_7291;
wire n_8102;
wire n_16449;
wire n_9540;
wire n_14840;
wire n_15859;
wire n_17939;
wire n_13033;
wire n_9753;
wire n_5780;
wire n_8460;
wire n_9105;
wire n_13746;
wire n_5643;
wire n_11305;
wire n_10149;
wire n_16088;
wire n_12680;
wire n_13017;
wire n_14530;
wire n_11137;
wire n_11607;
wire n_5846;
wire n_17202;
wire n_7430;
wire n_9700;
wire n_14234;
wire n_15511;
wire n_12930;
wire n_13914;
wire n_13752;
wire n_15093;
wire n_8871;
wire n_10649;
wire n_14360;
wire n_9476;
wire n_12722;
wire n_7870;
wire n_17910;
wire n_13529;
wire n_17390;
wire n_9875;
wire n_11265;
wire n_10593;
wire n_12042;
wire n_5524;
wire n_8824;
wire n_14827;
wire n_16671;
wire n_10597;
wire n_9963;
wire n_6104;
wire n_6475;
wire n_12469;
wire n_8470;
wire n_9582;
wire n_16058;
wire n_16641;
wire n_12172;
wire n_15533;
wire n_18029;
wire n_11739;
wire n_10817;
wire n_16919;
wire n_6465;
wire n_10060;
wire n_16810;
wire n_9574;
wire n_17690;
wire n_16459;
wire n_12049;
wire n_6496;
wire n_13229;
wire n_13973;
wire n_11687;
wire n_14160;
wire n_9732;
wire n_11050;
wire n_13070;
wire n_15576;
wire n_14440;
wire n_12666;
wire n_17769;
wire n_8238;
wire n_9882;
wire n_12205;
wire n_6998;
wire n_10779;
wire n_13177;
wire n_15230;
wire n_6145;
wire n_11789;
wire n_16239;
wire n_17051;
wire n_8699;
wire n_14946;
wire n_7305;
wire n_13878;
wire n_10242;
wire n_10086;
wire n_16135;
wire n_9992;
wire n_12885;
wire n_14899;
wire n_15204;
wire n_11347;
wire n_17641;
wire n_15899;
wire n_14166;
wire n_16488;
wire n_17067;
wire n_7980;
wire n_14363;
wire n_11617;
wire n_14952;
wire n_7075;
wire n_7545;
wire n_11581;
wire n_17078;
wire n_7846;
wire n_10981;
wire n_6076;
wire n_14626;
wire n_8438;
wire n_14831;
wire n_6194;
wire n_10673;
wire n_10869;
wire n_7695;
wire n_16549;
wire n_5066;
wire n_13850;
wire n_12917;
wire n_6092;
wire n_7275;
wire n_15254;
wire n_5401;
wire n_6357;
wire n_17564;
wire n_5843;
wire n_8095;
wire n_12616;
wire n_7537;
wire n_13690;
wire n_18176;
wire n_14356;
wire n_14429;
wire n_14705;
wire n_10128;
wire n_10746;
wire n_12287;
wire n_12217;
wire n_12950;
wire n_15845;
wire n_16644;
wire n_7489;
wire n_5106;
wire n_10339;
wire n_15572;
wire n_18016;
wire n_11559;
wire n_14629;
wire n_18121;
wire n_18005;
wire n_5468;
wire n_11867;
wire n_15197;
wire n_17903;
wire n_6335;
wire n_8112;
wire n_12835;
wire n_14727;
wire n_14343;
wire n_5883;
wire n_6985;
wire n_8642;
wire n_5319;
wire n_16516;
wire n_14996;
wire n_15072;
wire n_13552;
wire n_13432;
wire n_15800;
wire n_7451;
wire n_8624;
wire n_16161;
wire n_17856;
wire n_6238;
wire n_17474;
wire n_9090;
wire n_17647;
wire n_14066;
wire n_15780;
wire n_11989;
wire n_12800;
wire n_13495;
wire n_10684;
wire n_16677;
wire n_15030;
wire n_10441;
wire n_12036;
wire n_12177;
wire n_9149;
wire n_10590;
wire n_9174;
wire n_12850;
wire n_17762;
wire n_11175;
wire n_12962;
wire n_17378;
wire n_17243;
wire n_6548;
wire n_17866;
wire n_14755;
wire n_17210;
wire n_5455;
wire n_8894;
wire n_17440;
wire n_9226;
wire n_5706;
wire n_6366;
wire n_5337;
wire n_9018;
wire n_12336;
wire n_10949;
wire n_17317;
wire n_18066;
wire n_7236;
wire n_9835;
wire n_12044;
wire n_15135;
wire n_11727;
wire n_12905;
wire n_7269;
wire n_8878;
wire n_17625;
wire n_15663;
wire n_15706;
wire n_5223;
wire n_10934;
wire n_5962;
wire n_6602;
wire n_14018;
wire n_6620;
wire n_6502;
wire n_15856;
wire n_9702;
wire n_13409;
wire n_17633;
wire n_7560;
wire n_15348;
wire n_11725;
wire n_15565;
wire n_10279;
wire n_11291;
wire n_15138;
wire n_7326;
wire n_13548;
wire n_7060;
wire n_15643;
wire n_16618;
wire n_7572;
wire n_15301;
wire n_17062;
wire n_17351;
wire n_6885;
wire n_12495;
wire n_13139;
wire n_17407;
wire n_8807;
wire n_14207;
wire n_12565;
wire n_17083;
wire n_18147;
wire n_9968;
wire n_5074;
wire n_16328;
wire n_16957;
wire n_5364;
wire n_9924;
wire n_16848;
wire n_6529;
wire n_8732;
wire n_8169;
wire n_15174;
wire n_11958;
wire n_15954;
wire n_16950;
wire n_17257;
wire n_16207;
wire n_8803;
wire n_9515;
wire n_17835;
wire n_8017;
wire n_10527;
wire n_13506;
wire n_5895;
wire n_14756;
wire n_6951;
wire n_17294;
wire n_8801;
wire n_17140;
wire n_12584;
wire n_14258;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_7169;
wire n_12654;
wire n_13255;
wire n_6423;
wire n_9252;
wire n_15017;
wire n_14938;
wire n_15779;
wire n_10785;
wire n_7140;
wire n_7233;
wire n_10228;
wire n_11311;
wire n_12999;
wire n_14084;
wire n_13120;
wire n_5088;
wire n_6558;
wire n_8522;
wire n_5457;
wire n_16596;
wire n_15123;
wire n_7352;
wire n_15863;
wire n_7986;
wire n_15869;
wire n_9948;
wire n_7134;
wire n_5532;
wire n_12823;
wire n_11528;
wire n_12422;
wire n_6950;
wire n_7246;
wire n_18198;
wire n_12234;
wire n_6525;
wire n_7650;
wire n_9871;
wire n_11807;
wire n_16657;
wire n_14907;
wire n_6631;
wire n_6892;
wire n_11705;
wire n_8203;
wire n_15162;
wire n_15678;
wire n_14587;
wire n_15653;
wire n_16988;
wire n_17267;
wire n_7663;
wire n_13125;
wire n_15566;
wire n_9423;
wire n_11378;
wire n_11521;
wire n_11998;
wire n_17780;
wire n_9660;
wire n_14513;
wire n_9108;
wire n_14472;
wire n_11222;
wire n_15562;
wire n_16917;
wire n_15015;
wire n_14910;
wire n_8680;
wire n_9631;
wire n_10643;
wire n_7056;
wire n_14590;
wire n_12293;
wire n_16130;
wire n_10427;
wire n_6683;
wire n_8727;
wire n_15333;
wire n_17178;
wire n_17136;
wire n_10389;
wire n_13069;
wire n_13254;
wire n_16211;
wire n_15658;
wire n_10423;
wire n_6292;
wire n_5544;
wire n_15094;
wire n_16573;
wire n_9900;
wire n_14042;
wire n_15305;
wire n_11080;
wire n_7729;
wire n_7339;
wire n_7740;
wire n_5987;
wire n_6180;
wire n_17157;
wire n_5352;
wire n_16258;
wire n_5824;
wire n_16767;
wire n_14409;
wire n_11533;
wire n_12572;
wire n_5538;
wire n_8138;
wire n_17258;
wire n_6658;
wire n_10863;
wire n_6264;
wire n_9608;
wire n_9137;
wire n_15344;
wire n_6925;
wire n_8990;
wire n_15616;
wire n_16529;
wire n_5919;
wire n_10077;
wire n_12988;
wire n_16698;
wire n_17539;
wire n_8206;
wire n_9144;
wire n_17973;
wire n_12512;
wire n_7767;
wire n_11940;
wire n_13736;
wire n_8190;
wire n_6176;
wire n_13727;
wire n_9778;
wire n_16009;
wire n_8622;
wire n_13352;
wire n_15247;
wire n_5410;
wire n_11808;
wire n_13986;
wire n_15035;
wire n_7146;
wire n_18253;
wire n_8092;
wire n_13953;
wire n_15520;
wire n_10250;
wire n_15819;
wire n_7672;
wire n_6124;
wire n_14251;
wire n_8242;
wire n_17920;
wire n_12118;
wire n_12609;
wire n_14053;
wire n_14494;
wire n_7482;
wire n_12176;
wire n_14503;
wire n_9850;
wire n_14940;
wire n_6864;
wire n_9531;
wire n_13453;
wire n_7893;
wire n_8331;
wire n_15921;
wire n_17144;
wire n_7090;
wire n_17826;
wire n_15105;
wire n_16887;
wire n_11549;
wire n_16123;
wire n_7158;
wire n_17849;
wire n_14174;
wire n_15644;
wire n_7156;
wire n_5742;
wire n_5992;
wire n_8649;
wire n_15438;
wire n_16244;
wire n_8684;
wire n_6494;
wire n_17416;
wire n_5503;
wire n_18093;
wire n_8323;
wire n_10828;
wire n_12353;
wire n_6199;
wire n_17745;
wire n_11139;
wire n_8296;
wire n_13846;
wire n_9139;
wire n_11584;
wire n_17615;
wire n_9430;
wire n_10417;
wire n_5958;
wire n_6614;
wire n_7749;
wire n_15059;
wire n_11695;
wire n_16148;
wire n_17413;
wire n_7839;
wire n_8882;
wire n_10310;
wire n_12053;
wire n_7504;
wire n_10333;
wire n_10996;
wire n_13583;
wire n_12795;
wire n_16628;
wire n_9272;
wire n_10880;
wire n_8708;
wire n_17850;
wire n_12045;
wire n_7360;
wire n_10810;
wire n_12274;
wire n_7681;
wire n_10636;
wire n_12348;
wire n_8448;
wire n_8076;
wire n_7301;
wire n_9041;
wire n_11360;
wire n_16715;
wire n_5129;
wire n_11886;
wire n_9643;
wire n_8904;
wire n_7375;
wire n_7102;
wire n_5500;
wire n_8277;
wire n_11920;
wire n_15215;
wire n_7794;
wire n_11479;
wire n_13388;
wire n_12006;
wire n_7366;
wire n_16196;
wire n_8184;
wire n_13344;
wire n_5219;
wire n_13336;
wire n_14516;
wire n_15851;
wire n_5605;
wire n_9944;
wire n_14103;
wire n_16245;
wire n_5170;
wire n_16664;
wire n_5654;
wire n_7025;
wire n_8304;
wire n_5320;
wire n_13915;
wire n_18318;
wire n_14935;
wire n_10258;
wire n_11534;
wire n_6947;
wire n_16315;
wire n_8586;
wire n_5107;
wire n_9648;
wire n_5999;
wire n_9376;
wire n_8557;
wire n_10507;
wire n_16184;
wire n_8636;
wire n_7309;
wire n_13885;
wire n_6863;
wire n_9288;
wire n_10835;
wire n_6637;
wire n_15240;
wire n_15507;
wire n_6100;
wire n_13259;
wire n_7860;
wire n_6735;
wire n_14815;
wire n_9521;
wire n_9541;
wire n_13477;
wire n_8212;
wire n_17151;
wire n_6358;
wire n_9759;
wire n_14737;
wire n_12500;
wire n_13204;
wire n_12781;
wire n_16038;
wire n_16675;
wire n_7911;
wire n_15469;
wire n_13085;
wire n_15455;
wire n_11848;
wire n_8530;
wire n_9278;
wire n_16497;
wire n_9378;
wire n_11227;
wire n_8665;
wire n_5602;
wire n_9456;
wire n_13778;
wire n_9086;
wire n_7876;
wire n_15532;
wire n_6050;
wire n_11401;
wire n_15329;
wire n_15164;
wire n_14925;
wire n_9711;
wire n_8933;
wire n_14805;
wire n_13206;
wire n_16321;
wire n_15309;
wire n_7244;
wire n_15709;
wire n_16869;
wire n_7960;
wire n_5405;
wire n_13462;
wire n_12922;
wire n_14123;
wire n_5253;
wire n_17812;
wire n_17837;
wire n_9485;
wire n_11375;
wire n_9555;
wire n_10959;
wire n_7610;
wire n_12842;
wire n_9999;
wire n_11813;
wire n_14353;
wire n_9994;
wire n_10814;
wire n_5903;
wire n_6371;
wire n_16973;
wire n_17950;
wire n_8690;
wire n_17663;
wire n_8538;
wire n_7043;
wire n_16933;
wire n_12753;
wire n_16248;
wire n_16945;
wire n_15214;
wire n_10859;
wire n_6171;
wire n_7751;
wire n_8643;
wire n_15366;
wire n_6510;
wire n_15430;
wire n_17200;
wire n_6468;
wire n_9142;
wire n_9613;
wire n_11134;
wire n_9440;
wire n_11716;
wire n_5491;
wire n_8825;
wire n_12366;
wire n_7788;
wire n_14548;
wire n_5842;
wire n_6352;
wire n_8300;
wire n_13954;
wire n_10531;
wire n_14419;
wire n_5722;
wire n_7534;
wire n_9462;
wire n_7719;
wire n_5636;
wire n_11357;
wire n_9202;
wire n_16652;
wire n_18169;
wire n_5065;
wire n_7287;
wire n_10699;
wire n_12208;
wire n_7032;
wire n_17873;
wire n_8451;
wire n_11386;
wire n_13383;
wire n_14161;
wire n_5492;
wire n_9237;
wire n_10941;
wire n_11448;
wire n_5084;
wire n_10567;
wire n_6850;
wire n_8435;
wire n_17232;
wire n_5667;
wire n_18012;
wire n_16120;
wire n_12122;
wire n_14600;
wire n_10770;
wire n_5260;
wire n_16612;
wire n_11693;
wire n_7119;
wire n_8835;
wire n_13728;
wire n_15038;
wire n_10714;
wire n_9788;
wire n_13584;
wire n_15358;
wire n_13722;
wire n_5328;
wire n_14060;
wire n_14936;
wire n_16145;
wire n_6354;
wire n_7634;
wire n_5918;
wire n_14634;
wire n_16527;
wire n_11755;
wire n_17401;
wire n_6959;
wire n_6909;
wire n_16329;
wire n_17975;
wire n_16859;
wire n_11221;
wire n_7851;
wire n_6332;
wire n_9807;
wire n_14613;
wire n_13567;
wire n_13642;
wire n_7006;
wire n_15473;
wire n_15912;
wire n_17180;
wire n_9573;
wire n_17644;
wire n_5877;
wire n_8963;
wire n_12351;
wire n_6306;
wire n_7682;
wire n_15659;
wire n_14297;
wire n_13618;
wire n_18254;
wire n_17885;
wire n_6434;
wire n_12040;
wire n_12443;
wire n_16958;
wire n_8713;
wire n_17107;
wire n_6751;
wire n_7068;
wire n_9392;
wire n_12133;
wire n_11084;
wire n_13371;
wire n_14573;
wire n_16474;
wire n_6322;
wire n_14048;
wire n_8353;
wire n_8668;
wire n_13301;
wire n_5454;
wire n_9390;
wire n_16327;
wire n_17577;
wire n_13492;
wire n_14376;
wire n_7704;
wire n_16924;
wire n_10326;
wire n_7773;
wire n_17735;
wire n_9416;
wire n_14728;
wire n_6667;
wire n_7526;
wire n_13333;
wire n_8817;
wire n_6530;
wire n_9518;
wire n_15578;
wire n_13329;
wire n_12491;
wire n_7376;
wire n_13826;
wire n_6156;
wire n_13966;
wire n_14498;
wire n_5913;
wire n_7268;
wire n_16198;
wire n_7044;
wire n_12452;
wire n_5621;
wire n_13788;
wire n_13437;
wire n_16082;
wire n_8213;
wire n_12233;
wire n_18323;
wire n_8591;
wire n_7973;
wire n_11885;
wire n_16357;
wire n_6429;
wire n_16335;
wire n_18304;
wire n_13423;
wire n_10966;
wire n_5165;
wire n_15914;
wire n_7239;
wire n_17139;
wire n_10047;
wire n_16319;
wire n_12633;
wire n_5573;
wire n_11253;
wire n_6405;
wire n_11551;
wire n_14761;
wire n_8532;
wire n_11380;
wire n_12936;
wire n_15199;
wire n_12035;
wire n_17805;
wire n_13928;
wire n_6613;
wire n_8043;
wire n_9196;
wire n_11172;
wire n_13947;
wire n_14420;
wire n_17594;
wire n_15584;
wire n_7969;
wire n_6248;
wire n_17858;
wire n_18018;
wire n_17104;
wire n_14059;
wire n_15462;
wire n_12915;
wire n_7821;
wire n_15854;
wire n_6088;
wire n_17582;
wire n_12275;
wire n_10784;
wire n_5529;
wire n_10248;
wire n_6894;
wire n_12947;
wire n_14678;
wire n_7267;
wire n_9589;
wire n_5800;
wire n_11539;
wire n_9898;
wire n_14520;
wire n_15224;
wire n_16344;
wire n_13257;
wire n_17599;
wire n_17061;
wire n_9373;
wire n_11976;
wire n_17896;
wire n_12308;
wire n_13063;
wire n_8606;
wire n_17079;
wire n_14669;
wire n_15702;
wire n_6204;
wire n_10351;
wire n_13834;
wire n_17827;
wire n_13951;
wire n_15236;
wire n_17329;
wire n_16110;
wire n_7915;
wire n_8121;
wire n_8868;
wire n_10408;
wire n_10921;
wire n_13340;
wire n_7387;
wire n_7431;
wire n_11731;
wire n_7654;
wire n_10551;
wire n_12760;
wire n_16783;
wire n_10656;
wire n_16330;
wire n_16622;
wire n_6296;
wire n_11531;
wire n_12318;
wire n_13379;
wire n_15624;
wire n_10313;
wire n_10639;
wire n_15557;
wire n_5257;
wire n_16012;
wire n_9983;
wire n_6290;
wire n_14983;
wire n_6288;
wire n_12700;
wire n_14517;
wire n_8276;
wire n_8718;
wire n_12364;
wire n_8182;
wire n_14512;
wire n_5645;
wire n_15540;
wire n_11392;
wire n_17252;
wire n_5180;
wire n_13490;
wire n_13025;
wire n_11204;
wire n_13672;
wire n_13754;
wire n_14785;
wire n_15923;
wire n_12985;
wire n_5779;
wire n_11627;
wire n_13697;
wire n_12340;
wire n_12478;
wire n_6140;
wire n_16911;
wire n_9039;
wire n_13744;
wire n_8359;
wire n_7441;
wire n_9849;
wire n_16345;
wire n_8597;
wire n_6211;
wire n_12788;
wire n_8562;
wire n_13470;
wire n_11485;
wire n_16597;
wire n_8211;
wire n_13998;
wire n_13943;
wire n_16838;
wire n_9962;
wire n_14814;
wire n_17795;
wire n_16261;
wire n_12826;
wire n_8430;
wire n_17559;
wire n_6307;
wire n_8007;
wire n_10871;
wire n_6164;
wire n_12752;
wire n_15434;
wire n_7394;
wire n_8600;
wire n_8311;
wire n_8943;
wire n_8441;
wire n_12194;
wire n_16262;
wire n_10747;
wire n_7022;
wire n_15395;
wire n_16306;
wire n_9829;
wire n_14772;
wire n_13637;
wire n_15322;
wire n_6860;
wire n_10459;
wire n_16384;
wire n_8978;
wire n_10121;
wire n_15558;
wire n_11387;
wire n_8198;
wire n_9988;
wire n_14417;
wire n_5697;
wire n_14652;
wire n_17611;
wire n_14002;
wire n_15596;
wire n_15945;
wire n_16566;
wire n_7188;
wire n_8526;
wire n_10705;
wire n_13099;
wire n_7573;
wire n_17631;
wire n_7879;
wire n_16242;
wire n_9848;
wire n_7087;
wire n_18185;
wire n_6147;
wire n_14911;
wire n_17969;
wire n_16619;
wire n_10334;
wire n_7985;
wire n_16221;
wire n_17338;
wire n_12689;
wire n_11691;
wire n_11358;
wire n_18180;
wire n_9045;
wire n_9466;
wire n_6515;
wire n_15021;
wire n_9348;
wire n_6011;
wire n_8278;
wire n_16650;
wire n_7722;
wire n_7935;
wire n_8592;
wire n_15783;
wire n_6645;
wire n_11128;
wire n_12271;
wire n_13595;
wire n_17045;
wire n_14358;
wire n_14006;
wire n_8226;
wire n_15140;
wire n_16841;
wire n_6984;
wire n_12843;
wire n_16343;
wire n_13780;
wire n_10716;
wire n_12273;
wire n_17289;
wire n_10235;
wire n_13212;
wire n_15167;
wire n_13701;
wire n_10090;
wire n_13247;
wire n_10153;
wire n_16138;
wire n_14271;
wire n_15681;
wire n_11649;
wire n_10937;
wire n_13922;
wire n_7193;
wire n_10018;
wire n_13278;
wire n_8987;
wire n_16583;
wire n_16707;
wire n_17185;
wire n_13836;
wire n_11489;
wire n_6897;
wire n_7256;
wire n_12391;
wire n_5203;
wire n_12420;
wire n_17147;
wire n_14181;
wire n_9071;
wire n_17658;
wire n_10568;
wire n_9356;
wire n_9464;
wire n_12314;
wire n_6460;
wire n_7595;
wire n_7128;
wire n_9239;
wire n_10053;
wire n_6183;
wire n_10051;
wire n_11373;
wire n_7522;
wire n_5882;
wire n_13341;
wire n_15388;
wire n_16034;
wire n_9606;
wire n_13856;
wire n_17738;
wire n_10359;
wire n_7881;
wire n_14416;
wire n_14796;
wire n_14961;
wire n_15619;
wire n_16906;
wire n_18156;
wire n_7436;
wire n_15726;
wire n_7380;
wire n_7012;
wire n_11216;
wire n_12356;
wire n_10998;
wire n_15272;
wire n_7502;
wire n_9492;
wire n_13271;
wire n_17330;
wire n_8960;
wire n_7335;
wire n_7103;
wire n_13553;
wire n_10648;
wire n_10151;
wire n_6246;
wire n_14602;
wire n_14133;
wire n_11194;
wire n_11804;
wire n_18195;
wire n_17712;
wire n_8025;
wire n_5094;
wire n_6383;
wire n_9031;
wire n_15612;
wire n_15976;
wire n_16828;
wire n_17904;
wire n_11107;
wire n_9717;
wire n_11434;
wire n_9516;
wire n_11645;
wire n_12073;
wire n_15732;
wire n_16505;
wire n_18127;
wire n_7020;
wire n_8434;
wire n_11244;
wire n_17256;
wire n_12848;
wire n_8175;
wire n_9693;
wire n_9991;
wire n_5336;
wire n_15378;
wire n_12155;
wire n_13356;
wire n_14286;
wire n_17927;
wire n_9103;
wire n_8850;
wire n_11254;
wire n_14865;
wire n_13693;
wire n_16801;
wire n_9477;
wire n_15761;
wire n_16413;
wire n_14277;
wire n_17798;
wire n_5672;
wire n_13673;
wire n_5548;
wire n_10253;
wire n_10822;
wire n_7248;
wire n_7662;
wire n_5601;
wire n_14793;
wire n_8895;
wire n_10589;
wire n_12390;
wire n_12160;
wire n_13501;
wire n_15927;
wire n_11297;
wire n_10349;
wire n_11991;
wire n_5339;
wire n_13376;
wire n_6099;
wire n_10946;
wire n_12150;
wire n_5693;
wire n_8046;
wire n_11183;
wire n_11173;
wire n_6904;
wire n_17350;
wire n_11922;
wire n_16115;
wire n_13897;
wire n_18187;
wire n_8867;
wire n_15480;
wire n_17497;
wire n_15651;
wire n_16542;
wire n_10473;
wire n_8239;
wire n_9599;
wire n_13104;
wire n_7825;
wire n_8183;
wire n_8924;
wire n_9001;
wire n_12840;
wire n_10893;
wire n_15339;
wire n_16382;
wire n_13215;
wire n_17213;
wire n_10218;
wire n_13482;
wire n_16026;
wire n_17874;
wire n_12964;
wire n_5514;
wire n_13075;
wire n_5091;
wire n_7533;
wire n_8578;
wire n_11548;
wire n_9777;
wire n_8848;
wire n_13445;
wire n_10903;
wire n_10458;
wire n_11868;
wire n_13562;
wire n_9222;
wire n_16513;
wire n_18245;
wire n_10148;
wire n_15198;
wire n_6626;
wire n_6563;
wire n_5486;
wire n_9366;
wire n_6611;
wire n_10775;
wire n_11248;
wire n_10543;
wire n_17441;
wire n_9449;
wire n_15098;
wire n_15669;
wire n_11114;
wire n_17536;
wire n_16637;
wire n_18234;
wire n_11260;
wire n_11901;
wire n_12994;
wire n_5599;
wire n_14771;
wire n_6116;
wire n_16081;
wire n_15834;
wire n_18170;
wire n_7186;
wire n_10337;
wire n_16912;
wire n_8230;
wire n_9869;
wire n_10478;
wire n_12252;
wire n_11981;
wire n_16265;
wire n_15831;
wire n_6819;
wire n_8725;
wire n_13929;
wire n_5251;
wire n_7936;
wire n_13680;
wire n_13534;
wire n_6473;
wire n_16561;
wire n_12951;
wire n_13750;
wire n_9741;
wire n_13275;
wire n_11956;
wire n_10956;
wire n_10637;
wire n_13331;
wire n_16425;
wire n_13536;
wire n_15996;
wire n_11805;
wire n_15043;
wire n_5403;
wire n_12131;
wire n_12280;
wire n_8391;
wire n_7840;
wire n_6310;
wire n_10698;
wire n_15728;
wire n_16834;
wire n_17796;
wire n_11381;
wire n_16835;
wire n_14607;
wire n_9397;
wire n_8202;
wire n_12453;
wire n_11797;
wire n_11775;
wire n_17887;
wire n_10834;
wire n_7429;
wire n_18063;
wire n_17305;
wire n_6688;
wire n_12557;
wire n_16852;
wire n_7906;
wire n_8948;
wire n_8678;
wire n_9754;
wire n_18306;
wire n_16898;
wire n_15295;
wire n_10783;
wire n_9179;
wire n_17888;
wire n_7148;
wire n_15582;
wire n_5782;
wire n_8340;
wire n_6714;
wire n_7017;
wire n_7462;
wire n_7250;
wire n_7658;
wire n_7828;
wire n_8905;
wire n_12020;
wire n_13439;
wire n_8691;
wire n_13249;
wire n_12051;
wire n_6365;
wire n_16044;
wire n_16285;
wire n_16710;
wire n_10619;
wire n_14225;
wire n_13502;
wire n_16808;
wire n_13801;
wire n_5608;
wire n_13468;
wire n_11322;
wire n_12455;
wire n_18048;
wire n_10136;
wire n_7401;
wire n_13789;
wire n_8812;
wire n_12920;
wire n_14759;
wire n_13403;
wire n_9169;
wire n_6828;
wire n_12785;
wire n_16603;
wire n_14200;
wire n_11758;
wire n_17355;
wire n_5298;
wire n_16660;
wire n_17654;
wire n_8704;
wire n_6355;
wire n_5596;
wire n_7887;
wire n_11162;
wire n_13996;
wire n_8058;
wire n_12559;
wire n_16787;
wire n_16889;
wire n_9177;
wire n_10078;
wire n_6777;
wire n_5728;
wire n_11987;
wire n_16162;
wire n_16798;
wire n_8394;
wire n_10719;
wire n_9269;
wire n_7835;
wire n_12614;
wire n_13201;
wire n_14638;
wire n_15326;
wire n_11106;
wire n_9289;
wire n_8181;
wire n_10463;
wire n_12797;
wire n_13737;
wire n_13441;
wire n_14396;
wire n_17967;
wire n_14687;
wire n_8722;
wire n_10827;
wire n_12429;
wire n_6420;
wire n_6945;
wire n_11218;
wire n_9350;
wire n_7356;
wire n_5726;
wire n_7288;
wire n_7637;
wire n_7124;
wire n_10454;
wire n_11467;
wire n_12384;
wire n_7294;
wire n_12629;
wire n_12668;
wire n_13291;
wire n_16862;
wire n_16995;
wire n_12123;
wire n_5290;
wire n_12972;
wire n_14969;
wire n_7018;
wire n_13105;
wire n_10312;
wire n_11374;
wire n_17515;
wire n_11167;
wire n_13440;
wire n_12146;
wire n_7321;
wire n_9166;
wire n_10663;
wire n_10501;
wire n_5095;
wire n_10265;
wire n_10452;
wire n_15796;
wire n_8707;
wire n_6754;
wire n_10766;
wire n_12435;
wire n_13533;
wire n_11999;
wire n_6583;
wire n_13367;
wire n_17307;
wire n_6622;
wire n_6936;
wire n_13123;
wire n_8747;
wire n_16742;
wire n_5324;
wire n_7691;
wire n_15459;
wire n_5928;
wire n_8742;
wire n_10470;
wire n_10563;
wire n_12921;
wire n_16006;
wire n_7108;
wire n_6882;
wire n_15693;
wire n_11455;
wire n_16893;
wire n_7585;
wire n_13930;
wire n_9125;
wire n_7386;
wire n_10288;
wire n_8552;
wire n_18316;
wire n_5101;
wire n_12581;
wire n_5911;
wire n_7362;
wire n_7888;
wire n_7417;
wire n_12029;
wire n_12548;
wire n_17272;
wire n_9641;
wire n_14460;
wire n_9960;
wire n_7187;
wire n_13111;
wire n_11884;
wire n_5589;
wire n_5841;
wire n_13060;
wire n_12727;
wire n_10776;
wire n_11611;
wire n_9785;
wire n_9923;
wire n_8224;
wire n_17765;
wire n_16818;
wire n_17700;
wire n_10771;
wire n_7544;
wire n_11087;
wire n_14556;
wire n_5712;
wire n_11960;
wire n_6166;
wire n_8628;
wire n_13108;
wire n_11422;
wire n_13948;
wire n_18076;
wire n_6966;
wire n_13563;
wire n_17335;
wire n_7542;
wire n_6781;
wire n_9228;
wire n_14828;
wire n_7255;
wire n_15131;
wire n_12227;
wire n_8037;
wire n_8084;
wire n_17723;
wire n_7120;
wire n_7218;
wire n_12597;
wire n_16056;
wire n_16992;
wire n_7147;
wire n_14653;
wire n_7221;
wire n_15016;
wire n_15601;
wire n_16440;
wire n_10967;
wire n_8289;
wire n_9801;
wire n_14189;
wire n_16021;
wire n_10249;
wire n_11029;
wire n_15057;
wire n_17767;
wire n_9645;
wire n_16786;
wire n_8045;
wire n_11199;
wire n_17019;
wire n_15721;
wire n_5633;
wire n_8697;
wire n_13568;
wire n_13396;
wire n_13029;
wire n_13647;
wire n_8077;
wire n_17181;
wire n_17729;
wire n_15977;
wire n_6980;
wire n_12674;
wire n_5583;
wire n_17686;
wire n_11826;
wire n_9457;
wire n_15071;
wire n_8026;
wire n_11317;
wire n_13652;
wire n_7889;
wire n_6064;
wire n_6110;
wire n_10742;
wire n_6237;
wire n_16083;
wire n_14538;
wire n_7196;
wire n_12913;
wire n_10390;
wire n_9330;
wire n_6341;
wire n_10012;
wire n_9365;
wire n_14861;
wire n_15781;
wire n_17512;
wire n_6590;
wire n_5501;
wire n_8444;
wire n_9178;
wire n_8654;
wire n_14021;
wire n_16646;
wire n_17031;
wire n_10035;
wire n_10753;
wire n_9181;
wire n_12112;
wire n_7923;
wire n_13965;
wire n_16579;
wire n_14465;
wire n_5377;
wire n_11033;
wire n_18207;
wire n_6697;
wire n_13168;
wire n_6453;
wire n_5652;
wire n_6135;
wire n_13574;
wire n_14037;
wire n_7559;
wire n_11798;
wire n_15577;
wire n_12346;
wire n_17470;
wire n_11853;
wire n_7081;
wire n_9307;
wire n_15476;
wire n_10795;
wire n_10300;
wire n_10257;
wire n_15752;
wire n_6449;
wire n_7832;
wire n_7968;
wire n_17405;
wire n_17461;
wire n_9238;
wire n_12714;
wire n_11166;
wire n_11079;
wire n_13581;
wire n_6141;
wire n_10099;
wire n_18090;
wire n_8449;
wire n_17589;
wire n_11217;
wire n_12732;
wire n_13138;
wire n_14481;
wire n_10985;
wire n_18307;
wire n_15650;
wire n_14931;
wire n_8493;
wire n_7584;
wire n_9224;
wire n_10244;
wire n_12400;
wire n_17989;
wire n_6983;
wire n_12671;
wire n_7843;
wire n_17902;
wire n_13774;
wire n_10377;
wire n_6036;
wire n_11469;
wire n_10984;
wire n_12863;
wire n_18303;
wire n_12347;
wire n_15188;
wire n_8958;
wire n_10801;
wire n_11898;
wire n_8443;
wire n_17149;
wire n_12041;
wire n_17288;
wire n_9756;
wire n_7222;
wire n_9624;
wire n_6071;
wire n_8161;
wire n_13435;
wire n_17880;
wire n_16403;
wire n_11710;
wire n_6808;
wire n_8734;
wire n_9547;
wire n_11341;
wire n_8271;
wire n_9594;
wire n_9901;
wire n_11619;
wire n_16854;
wire n_11238;
wire n_9895;
wire n_10878;
wire n_13378;
wire n_6724;
wire n_15460;
wire n_9277;
wire n_11608;
wire n_14169;
wire n_18199;
wire n_16407;
wire n_14086;
wire n_12756;
wire n_6571;
wire n_16511;
wire n_17926;
wire n_15074;
wire n_5100;
wire n_7470;
wire n_9189;
wire n_15470;
wire n_16059;
wire n_5849;
wire n_8495;
wire n_6251;
wire n_7400;
wire n_14255;
wire n_9548;
wire n_16290;
wire n_14309;
wire n_12088;
wire n_16688;
wire n_12218;
wire n_14204;
wire n_17308;
wire n_6635;
wire n_10000;
wire n_9472;
wire n_16670;
wire n_17757;
wire n_13202;
wire n_14738;
wire n_13410;
wire n_11553;
wire n_14432;
wire n_16998;
wire n_5367;
wire n_13816;
wire n_8994;
wire n_15930;
wire n_16802;
wire n_8901;
wire n_8056;
wire n_10725;
wire n_12323;
wire n_14767;
wire n_17800;
wire n_17788;
wire n_9538;
wire n_7623;
wire n_12387;
wire n_14984;
wire n_10627;
wire n_8954;
wire n_13590;
wire n_15846;
wire n_17823;
wire n_5616;
wire n_13230;
wire n_7597;
wire n_11996;
wire n_6733;
wire n_7071;
wire n_17552;
wire n_16761;
wire n_15029;
wire n_8840;
wire n_6467;
wire n_5988;
wire n_7859;
wire n_6035;
wire n_8900;
wire n_13456;
wire n_17832;
wire n_15194;
wire n_10477;
wire n_14651;
wire n_13321;
wire n_15967;
wire n_12798;
wire n_17987;
wire n_14306;
wire n_16067;
wire n_11032;
wire n_6522;
wire n_7109;
wire n_11834;
wire n_14057;
wire n_9434;
wire n_10604;
wire n_11110;
wire n_5959;
wire n_9052;
wire n_7645;
wire n_17020;
wire n_6732;
wire n_18240;
wire n_13806;
wire n_6562;
wire n_16149;
wire n_12780;
wire n_9176;
wire n_6150;
wire n_10461;
wire n_12772;
wire n_10559;
wire n_18275;
wire n_15314;
wire n_17889;
wire n_17659;
wire n_11141;
wire n_8157;
wire n_12539;
wire n_13007;
wire n_8346;
wire n_9697;
wire n_16260;
wire n_15656;
wire n_13651;
wire n_7882;
wire n_13830;
wire n_8827;
wire n_13113;
wire n_16307;
wire n_8309;
wire n_13196;
wire n_14998;
wire n_8344;
wire n_5917;
wire n_12589;
wire n_9060;
wire n_5754;
wire n_6016;
wire n_12775;
wire n_8096;
wire n_8822;
wire n_8100;
wire n_15670;
wire n_12043;
wire n_9758;
wire n_7212;
wire n_7908;
wire n_15160;
wire n_8222;
wire n_17074;
wire n_14430;
wire n_16362;
wire n_10479;
wire n_17721;
wire n_16676;
wire n_18111;
wire n_9876;
wire n_5628;
wire n_10572;
wire n_11971;
wire n_6726;
wire n_8406;
wire n_10277;
wire n_11320;
wire n_14697;
wire n_16091;
wire n_11028;
wire n_5252;
wire n_7009;
wire n_6554;
wire n_10139;
wire n_10230;
wire n_15847;
wire n_14294;
wire n_17263;
wire n_18007;
wire n_6689;
wire n_15708;
wire n_16594;
wire n_17120;
wire n_14245;
wire n_12476;
wire n_14858;
wire n_8866;
wire n_13724;
wire n_6143;
wire n_5614;
wire n_8693;
wire n_5134;
wire n_17362;
wire n_10207;
wire n_12536;
wire n_15597;
wire n_16755;
wire n_11368;
wire n_11144;
wire n_16791;
wire n_7355;
wire n_16962;
wire n_7365;
wire n_15286;
wire n_8794;
wire n_7777;
wire n_9653;
wire n_6277;
wire n_14993;
wire n_7395;
wire n_5981;
wire n_11404;
wire n_15593;
wire n_12896;
wire n_13373;
wire n_16222;
wire n_6095;
wire n_16079;
wire n_7671;
wire n_10429;
wire n_17302;
wire n_15951;
wire n_8020;
wire n_17807;
wire n_14241;
wire n_12957;
wire n_13866;
wire n_16966;
wire n_6247;
wire n_10255;
wire n_9257;
wire n_13014;
wire n_17917;
wire n_15141;
wire n_15235;
wire n_9270;
wire n_6880;
wire n_10901;
wire n_15881;
wire n_10101;
wire n_5720;
wire n_15129;
wire n_14000;
wire n_13022;
wire n_17460;
wire n_13422;
wire n_5325;
wire n_13633;
wire n_15380;
wire n_5696;
wire n_12549;
wire n_5375;
wire n_8736;
wire n_6499;
wire n_12362;
wire n_6837;
wire n_17664;
wire n_17958;
wire n_17830;
wire n_13442;
wire n_17585;
wire n_14741;
wire n_14972;
wire n_15073;
wire n_17990;
wire n_10063;
wire n_13390;
wire n_12030;
wire n_7393;
wire n_14679;
wire n_8400;
wire n_6616;
wire n_9686;
wire n_13136;
wire n_13334;
wire n_13408;
wire n_14690;
wire n_13989;
wire n_15288;
wire n_16481;
wire n_7871;
wire n_14532;
wire n_14859;
wire n_12018;
wire n_10846;
wire n_6946;
wire n_10195;
wire n_8055;
wire n_8333;
wire n_11593;
wire n_11847;
wire n_15904;
wire n_9718;
wire n_11773;
wire n_14074;
wire n_14944;
wire n_5064;
wire n_9215;
wire n_5759;
wire n_12060;
wire n_5753;
wire n_10628;
wire n_8909;
wire n_16033;
wire n_17337;
wire n_5536;
wire n_15056;
wire n_7484;
wire n_5173;
wire n_11968;
wire n_6305;
wire n_13630;
wire n_14071;
wire n_16053;
wire n_14127;
wire n_17376;
wire n_6317;
wire n_9762;
wire n_9407;
wire n_10819;
wire n_12315;
wire n_12903;
wire n_13269;
wire n_14570;
wire n_5691;
wire n_13103;
wire n_15771;
wire n_15865;
wire n_5794;
wire n_13098;
wire n_16708;
wire n_11896;
wire n_17661;
wire n_16523;
wire n_5647;
wire n_7231;
wire n_11897;
wire n_14447;
wire n_13707;
wire n_10368;
wire n_12484;
wire n_14971;
wire n_7272;
wire n_9964;
wire n_13031;
wire n_13646;
wire n_5738;
wire n_7649;
wire n_9953;
wire n_17524;
wire n_10356;
wire n_17523;
wire n_14154;
wire n_17429;
wire n_16332;
wire n_5215;
wire n_7324;
wire n_9153;
wire n_6693;
wire n_8786;
wire n_10931;
wire n_8541;
wire n_11711;
wire n_12673;
wire n_6734;
wire n_12000;
wire n_16604;
wire n_16463;
wire n_18104;
wire n_10173;
wire n_15107;
wire n_9571;
wire n_7135;
wire n_11554;
wire n_7014;
wire n_8263;
wire n_10644;
wire n_11159;
wire n_8884;
wire n_13062;
wire n_5597;
wire n_5635;
wire n_13424;
wire n_17445;
wire n_10323;
wire n_11350;
wire n_17731;
wire n_9019;
wire n_6382;
wire n_11310;
wire n_17204;
wire n_13001;
wire n_7328;
wire n_7635;
wire n_6404;
wire n_12063;
wire n_15023;
wire n_10229;
wire n_10693;
wire n_5975;
wire n_9737;
wire n_11688;
wire n_13842;
wire n_16568;
wire n_10493;
wire n_11125;
wire n_8494;
wire n_10554;
wire n_6379;
wire n_10382;
wire n_11083;
wire n_7703;
wire n_7066;
wire n_9468;
wire n_7358;
wire n_12449;
wire n_10622;
wire n_13664;
wire n_11939;
wire n_6235;
wire n_16176;
wire n_16968;
wire n_13144;
wire n_9870;
wire n_7277;
wire n_6504;
wire n_18049;
wire n_9026;
wire n_13900;
wire n_9710;
wire n_15799;
wire n_17281;
wire n_7265;
wire n_8638;
wire n_11126;
wire n_15665;
wire n_15958;
wire n_8710;
wire n_10019;
wire n_13512;
wire n_16837;
wire n_15591;
wire n_6789;
wire n_15719;
wire n_7184;
wire n_11090;
wire n_6440;
wire n_17617;
wire n_9725;
wire n_11953;
wire n_6417;
wire n_14557;
wire n_12845;
wire n_16503;
wire n_16526;
wire n_18136;
wire n_8177;
wire n_14013;
wire n_15385;
wire n_18094;
wire n_12062;
wire n_12636;
wire n_14784;
wire n_7491;
wire n_5942;
wire n_14436;
wire n_15866;
wire n_16522;
wire n_16954;
wire n_14524;
wire n_9084;
wire n_7728;
wire n_17148;
wire n_10488;
wire n_17638;
wire n_10767;
wire n_7690;
wire n_15360;
wire n_13084;
wire n_15110;
wire n_7219;
wire n_13375;
wire n_7479;
wire n_11040;
wire n_13852;
wire n_11751;
wire n_9419;
wire n_12793;
wire n_13203;
wire n_11158;
wire n_14378;
wire n_7270;
wire n_5940;
wire n_8170;
wire n_12367;
wire n_10579;
wire n_14488;
wire n_8893;
wire n_13473;
wire n_14923;
wire n_12317;
wire n_7390;
wire n_17789;
wire n_15296;
wire n_15586;
wire n_16379;
wire n_17696;
wire n_7805;
wire n_10474;
wire n_7807;
wire n_5121;
wire n_9973;
wire n_9479;
wire n_8589;
wire n_9820;
wire n_13316;
wire n_12954;
wire n_12724;
wire n_17348;
wire n_11094;
wire n_16303;
wire n_16310;
wire n_8320;
wire n_5555;
wire n_6914;
wire n_7978;
wire n_15458;
wire n_15155;
wire n_12157;
wire n_16716;
wire n_15379;
wire n_17452;
wire n_14891;
wire n_18027;
wire n_11161;
wire n_11182;
wire n_10587;
wire n_15441;
wire n_7182;
wire n_12195;
wire n_11839;
wire n_15115;
wire n_11815;
wire n_5784;
wire n_10843;
wire n_12773;
wire n_8153;
wire n_6272;
wire n_7699;
wire n_6484;
wire n_7674;
wire n_12556;
wire n_17695;
wire n_6236;
wire n_8620;
wire n_10755;
wire n_5576;
wire n_8298;
wire n_11614;
wire n_6958;
wire n_5466;
wire n_6840;
wire n_13645;
wire n_17439;
wire n_6871;
wire n_12789;
wire n_10270;
wire n_11590;
wire n_12649;
wire n_8235;
wire n_17618;
wire n_15201;
wire n_11845;
wire n_5284;
wire n_9294;
wire n_9126;
wire n_8370;
wire n_13773;
wire n_11263;
wire n_16807;
wire n_11908;
wire n_13066;
wire n_15109;
wire n_17196;
wire n_5308;
wire n_17543;
wire n_13469;
wire n_10573;
wire n_13101;
wire n_6768;
wire n_13494;
wire n_13893;
wire n_7951;
wire n_15190;
wire n_16749;
wire n_10992;
wire n_14490;
wire n_17218;
wire n_7506;
wire n_14210;
wire n_16507;
wire n_17882;
wire n_14717;
wire n_18051;
wire n_12696;
wire n_6717;
wire n_13505;
wire n_11257;
wire n_17893;
wire n_18046;
wire n_7048;
wire n_11136;
wire n_11142;
wire n_15368;
wire n_10428;
wire n_13569;
wire n_15908;
wire n_16844;
wire n_16843;
wire n_18162;
wire n_18247;
wire n_16904;
wire n_16572;
wire n_12664;
wire n_15885;
wire n_5578;
wire n_8395;
wire n_10989;
wire n_13450;
wire n_11145;
wire n_12206;
wire n_11745;
wire n_13010;
wire n_15081;
wire n_15812;
wire n_14375;
wire n_13181;
wire n_11017;
wire n_16517;
wire n_10805;
wire n_15623;
wire n_8906;
wire n_10682;
wire n_5530;
wire n_11414;
wire n_8097;
wire n_10327;
wire n_12940;
wire n_14322;
wire n_7416;
wire n_6196;
wire n_18223;
wire n_15608;
wire n_10528;
wire n_5741;
wire n_8570;
wire n_8902;
wire n_12404;
wire n_5991;
wire n_13815;
wire n_10365;
wire n_7330;
wire n_15435;
wire n_15950;
wire n_7928;
wire n_12201;
wire n_5506;
wire n_17894;
wire n_5243;
wire n_15061;
wire n_9819;
wire n_18269;
wire n_8477;
wire n_5449;
wire n_16704;
wire n_10236;
wire n_16415;
wire n_5221;
wire n_6992;
wire n_10433;
wire n_13725;
wire n_13924;
wire n_12312;
wire n_15191;
wire n_10625;
wire n_6000;
wire n_16005;
wire n_10303;
wire n_9545;
wire n_7283;
wire n_7099;
wire n_11452;
wire n_15270;
wire n_10557;
wire n_5311;
wire n_6448;
wire n_11323;
wire n_16125;
wire n_13002;
wire n_6655;
wire n_12982;
wire n_7892;
wire n_9165;
wire n_11558;
wire n_17670;
wire n_14732;
wire n_15256;
wire n_7304;
wire n_10143;
wire n_13018;
wire n_5792;
wire n_13185;
wire n_14872;
wire n_15705;
wire n_14681;
wire n_12002;
wire n_15171;
wire n_6657;
wire n_7756;
wire n_18133;
wire n_8129;
wire n_13150;
wire n_5575;
wire n_8580;
wire n_11543;
wire n_7990;
wire n_15521;
wire n_8122;
wire n_17953;
wire n_11883;
wire n_17479;
wire n_10796;
wire n_8259;
wire n_8536;
wire n_18235;
wire n_7626;
wire n_7474;
wire n_17581;
wire n_10855;
wire n_8748;
wire n_7612;
wire n_17088;
wire n_6113;
wire n_16155;
wire n_7789;
wire n_9056;
wire n_15826;
wire n_8094;
wire n_18074;
wire n_9341;
wire n_14164;
wire n_11429;
wire n_14165;
wire n_6242;
wire n_7902;
wire n_7088;
wire n_15027;
wire n_6519;
wire n_10357;
wire n_16369;
wire n_8572;
wire n_16412;
wire n_10681;
wire n_8120;
wire n_12598;
wire n_6842;
wire n_12942;
wire n_12750;
wire n_13575;
wire n_12729;
wire n_17435;
wire n_7588;
wire n_12033;
wire n_6206;
wire n_6414;
wire n_17578;
wire n_16738;
wire n_11241;
wire n_17033;
wire n_9172;
wire n_17296;
wire n_14239;
wire n_12441;
wire n_9145;
wire n_13805;
wire n_6801;
wire n_8099;
wire n_17719;
wire n_9996;
wire n_11348;
wire n_10059;
wire n_10284;
wire n_7680;
wire n_8770;
wire n_5276;
wire n_6308;
wire n_14790;
wire n_7398;
wire n_6906;
wire n_14029;
wire n_5078;
wire n_11169;
wire n_11041;
wire n_17707;
wire n_16039;
wire n_7230;
wire n_8700;
wire n_11160;
wire n_16015;
wire n_9906;
wire n_6629;
wire n_10957;
wire n_14250;
wire n_12827;
wire n_16393;
wire n_17909;
wire n_11124;
wire n_16028;
wire n_6968;
wire n_9920;
wire n_9504;
wire n_16799;
wire n_16632;
wire n_6615;
wire n_7378;
wire n_15689;
wire n_16206;
wire n_12734;
wire n_12181;
wire n_9482;
wire n_15145;
wire n_5205;
wire n_14032;
wire n_16763;
wire n_14760;
wire n_16107;
wire n_9138;
wire n_11152;
wire n_9384;
wire n_8637;
wire n_5651;
wire n_6144;
wire n_8757;
wire n_17059;
wire n_6188;
wire n_17727;
wire n_14794;
wire n_5819;
wire n_10147;
wire n_14197;
wire n_13765;
wire n_8903;
wire n_13709;
wire n_9193;
wire n_15962;
wire n_5998;
wire n_18288;
wire n_6398;
wire n_11586;
wire n_14660;
wire n_17133;
wire n_12069;
wire n_11990;
wire n_17570;
wire n_5721;
wire n_5673;
wire n_9527;
wire n_14554;
wire n_17899;
wire n_17387;
wire n_5351;
wire n_10889;
wire n_12363;
wire n_11019;
wire n_14028;
wire n_15788;
wire n_13170;
wire n_14368;
wire n_14699;
wire n_8585;
wire n_9064;
wire n_18326;
wire n_14056;
wire n_8982;
wire n_6415;
wire n_10816;
wire n_16428;
wire n_14374;
wire n_10032;
wire n_13385;
wire n_18155;
wire n_6857;
wire n_17756;
wire n_10489;
wire n_15114;
wire n_5476;
wire n_10200;
wire n_12442;
wire n_7842;
wire n_10898;
wire n_12499;
wire n_5856;
wire n_14588;
wire n_8709;
wire n_5446;
wire n_9383;
wire n_10825;
wire n_17937;
wire n_6722;
wire n_9735;
wire n_9943;
wire n_16714;
wire n_10290;
wire n_6428;
wire n_17717;
wire n_18075;
wire n_15853;
wire n_5944;
wire n_7618;
wire n_15569;
wire n_15862;
wire n_12818;
wire n_15078;
wire n_16267;
wire n_16358;
wire n_17764;
wire n_6413;
wire n_7679;
wire n_11132;
wire n_13684;
wire n_6361;
wire n_11677;
wire n_9357;
wire n_16468;
wire n_13608;
wire n_10680;
wire n_12531;
wire n_7783;
wire n_6231;
wire n_11036;
wire n_15394;
wire n_14826;
wire n_5684;
wire n_16897;
wire n_5861;
wire n_11927;
wire n_8108;
wire n_10306;
wire n_5976;
wire n_17681;
wire n_15445;
wire n_11827;
wire n_7862;
wire n_16896;
wire n_5312;
wire n_10675;
wire n_5850;
wire n_10014;
wire n_16150;
wire n_13454;
wire n_17933;
wire n_5111;
wire n_16117;
wire n_13829;
wire n_17070;
wire n_5890;
wire n_15968;
wire n_9986;
wire n_10355;
wire n_13758;
wire n_16409;
wire n_10830;
wire n_16905;
wire n_7820;
wire n_7167;
wire n_8692;
wire n_14967;
wire n_17025;
wire n_7833;
wire n_11118;
wire n_8820;
wire n_12496;
wire n_14750;
wire n_15454;
wire n_7643;
wire n_12460;
wire n_17347;
wire n_17127;
wire n_13586;
wire n_8490;
wire n_10380;
wire n_5113;
wire n_9491;
wire n_16829;
wire n_12821;
wire n_15028;
wire n_15736;
wire n_14809;
wire n_9922;
wire n_6712;
wire n_17583;
wire n_5687;
wire n_12479;
wire n_10530;
wire n_13703;
wire n_8062;
wire n_16299;
wire n_8781;
wire n_10999;
wire n_16826;
wire n_10203;
wire n_8000;
wire n_10061;
wire n_13860;
wire n_10899;
wire n_18282;
wire n_10961;
wire n_8808;
wire n_13359;
wire n_8233;
wire n_15573;
wire n_5839;
wire n_9747;
wire n_11811;
wire n_16620;
wire n_6953;
wire n_8685;
wire n_13877;
wire n_15097;
wire n_9061;
wire n_9168;
wire n_12361;
wire n_11561;
wire n_12345;
wire n_18220;
wire n_8575;
wire n_8701;
wire n_11690;
wire n_17369;
wire n_15126;
wire n_11212;
wire n_6303;
wire n_12593;
wire n_6474;
wire n_6182;
wire n_16114;
wire n_11155;
wire n_15118;
wire n_5674;
wire n_8670;
wire n_6573;
wire n_13151;
wire n_6053;
wire n_14380;
wire n_7234;
wire n_10425;
wire n_15060;
wire n_8352;
wire n_7993;
wire n_7930;
wire n_5682;
wire n_12984;
wire n_15170;
wire n_16194;
wire n_16094;
wire n_8385;
wire n_14330;
wire n_8875;
wire n_6392;
wire n_8166;
wire n_11433;
wire n_18069;
wire n_5167;
wire n_16496;
wire n_9073;
wire n_8934;
wire n_5117;
wire n_17843;
wire n_17090;
wire n_11312;
wire n_15928;
wire n_11477;
wire n_7999;
wire n_5612;
wire n_14347;
wire n_11988;
wire n_7963;
wire n_6125;
wire n_6599;
wire n_14978;
wire n_15485;
wire n_6685;
wire n_12311;
wire n_12914;
wire n_15213;
wire n_18079;
wire n_11964;
wire n_12086;
wire n_8389;
wire n_9068;
wire n_15289;
wire n_10537;
wire n_17203;
wire n_10158;
wire n_14823;
wire n_6560;
wire n_12787;
wire n_14686;
wire n_17747;
wire n_10711;
wire n_11933;
wire n_8659;
wire n_8804;
wire n_18105;
wire n_10043;
wire n_18001;
wire n_16460;
wire n_12703;
wire n_12411;
wire n_6253;
wire n_7382;
wire n_17417;
wire n_8439;
wire n_13337;
wire n_9544;
wire n_14108;
wire n_8814;
wire n_8369;
wire n_17753;
wire n_13867;
wire n_5301;
wire n_11574;
wire n_7800;
wire n_15575;
wire n_10930;
wire n_7615;
wire n_9286;
wire n_5898;
wire n_11313;
wire n_16937;
wire n_14700;
wire n_16408;
wire n_17853;
wire n_15633;
wire n_11206;
wire n_12263;
wire n_7298;
wire n_16406;
wire n_12959;
wire n_10131;
wire n_7581;
wire n_15238;
wire n_18160;
wire n_6641;
wire n_5214;
wire n_13057;
wire n_13551;
wire n_5563;
wire n_5487;
wire n_6593;
wire n_12461;
wire n_6673;
wire n_10696;
wire n_12893;
wire n_13990;
wire n_17131;
wire n_8789;
wire n_7172;
wire n_17876;
wire n_7074;
wire n_10685;
wire n_5497;
wire n_8790;
wire n_11223;
wire n_8234;
wire n_16486;
wire n_16872;
wire n_17358;
wire n_11624;
wire n_18010;
wire n_5832;
wire n_16325;
wire n_13876;
wire n_18041;
wire n_13791;
wire n_14438;
wire n_16614;
wire n_7190;
wire n_11515;
wire n_7112;
wire n_14382;
wire n_13128;
wire n_16217;
wire n_13807;
wire n_13142;
wire n_16747;
wire n_7678;
wire n_10082;
wire n_15299;
wire n_9265;
wire n_17197;
wire n_11560;
wire n_15390;
wire n_13678;
wire n_17683;
wire n_9080;
wire n_13433;
wire n_5526;
wire n_8989;
wire n_10152;
wire n_15063;
wire n_13589;
wire n_12645;
wire n_6367;
wire n_6195;
wire n_6356;
wire n_8927;
wire n_14192;
wire n_11055;
wire n_17238;
wire n_18309;
wire n_18256;
wire n_16703;
wire n_17649;
wire n_11616;
wire n_9770;
wire n_15824;
wire n_14746;
wire n_9463;
wire n_7001;
wire n_12090;
wire n_13481;
wire n_13743;
wire n_5593;
wire n_6514;
wire n_7369;
wire n_17759;
wire n_5444;
wire n_10580;
wire n_16759;
wire n_14365;
wire n_7829;
wire n_14131;
wire n_9939;
wire n_10159;
wire n_11390;
wire n_8534;
wire n_9911;
wire n_9210;
wire n_6559;
wire n_5211;
wire n_5230;
wire n_10122;
wire n_10302;
wire n_14457;
wire n_7359;
wire n_14398;
wire n_5389;
wire n_15443;
wire n_7144;
wire n_10462;
wire n_14244;
wire n_13357;
wire n_17106;
wire n_8756;
wire n_6841;
wire n_16351;
wire n_14320;
wire n_11597;
wire n_14918;
wire n_16252;
wire n_11002;
wire n_13716;
wire n_17915;
wire n_16631;
wire n_9691;
wire n_5110;
wire n_16223;
wire n_6653;
wire n_16045;
wire n_12165;
wire n_17208;
wire n_15970;
wire n_16552;
wire n_7450;
wire n_5425;
wire n_13803;
wire n_16316;
wire n_14455;
wire n_17518;
wire n_10532;
wire n_8832;
wire n_17015;
wire n_15583;
wire n_15614;
wire n_5737;
wire n_16544;
wire n_15178;
wire n_16151;
wire n_9340;
wire n_10350;
wire n_16431;
wire n_9351;
wire n_8461;
wire n_8042;
wire n_11179;
wire n_10977;
wire n_15128;
wire n_6825;
wire n_6923;
wire n_11708;
wire n_15108;
wire n_17027;
wire n_9950;
wire n_10418;
wire n_11474;
wire n_15889;
wire n_10336;
wire n_18008;
wire n_8021;
wire n_8839;
wire n_12092;
wire n_11369;
wire n_17205;
wire n_6112;
wire n_11738;
wire n_6547;
wire n_14113;
wire n_11240;
wire n_6198;
wire n_13155;
wire n_7439;
wire n_5560;
wire n_15483;
wire n_18243;
wire n_12074;
wire n_9155;
wire n_17353;
wire n_14565;
wire n_11931;
wire n_14231;
wire n_15841;
wire n_10925;
wire n_6399;
wire n_8623;
wire n_15277;
wire n_16824;
wire n_12109;
wire n_11438;
wire n_8758;
wire n_14508;
wire n_6275;
wire n_6575;
wire n_5666;
wire n_17379;
wire n_10609;
wire n_13508;
wire n_17785;
wire n_7924;
wire n_16338;
wire n_7732;
wire n_6151;
wire n_13058;
wire n_18036;
wire n_17242;
wire n_17588;
wire n_5179;
wire n_7227;
wire n_7040;
wire n_15042;
wire n_8511;
wire n_7325;
wire n_6469;
wire n_6756;
wire n_8595;
wire n_12900;
wire n_8873;
wire n_11376;
wire n_17155;
wire n_9201;
wire n_5961;
wire n_7459;
wire n_7191;
wire n_9823;
wire n_11051;
wire n_14304;
wire n_15530;
wire n_11812;
wire n_9688;
wire n_12330;
wire n_7096;
wire n_12519;
wire n_13872;
wire n_17280;
wire n_13597;
wire n_8455;
wire n_17918;
wire n_11838;
wire n_17057;
wire n_12717;
wire n_17150;
wire n_8280;
wire n_10102;
wire n_11333;
wire n_10908;
wire n_9595;
wire n_5272;
wire n_15119;
wire n_9530;
wire n_6826;
wire n_9227;
wire n_6015;
wire n_8372;
wire n_5361;
wire n_8598;
wire n_5683;
wire n_10939;
wire n_13503;
wire n_11178;
wire n_18322;
wire n_12595;
wire n_5847;
wire n_7551;
wire n_18246;
wire n_9400;
wire n_6678;
wire n_11188;
wire n_5068;
wire n_16540;
wire n_9025;
wire n_16543;
wire n_5740;
wire n_16528;
wire n_18039;
wire n_17705;
wire n_16456;
wire n_13086;
wire n_17001;
wire n_8282;
wire n_7750;
wire n_10936;
wire n_17934;
wire n_11840;
wire n_18226;
wire n_12525;
wire n_17400;
wire n_7697;
wire n_5729;
wire n_7485;
wire n_11685;
wire n_17982;
wire n_10955;
wire n_13093;
wire n_10824;
wire n_6748;
wire n_15673;
wire n_12084;
wire n_8616;
wire n_10440;
wire n_10630;
wire n_8336;
wire n_16493;
wire n_17854;
wire n_5302;
wire n_17228;
wire n_11472;
wire n_16948;
wire n_6752;
wire n_9749;
wire n_14404;
wire n_5545;
wire n_17651;
wire n_6553;
wire n_9285;
wire n_12997;
wire n_11295;
wire n_9972;
wire n_10058;
wire n_7652;
wire n_14533;
wire n_8847;
wire n_7808;
wire n_11171;
wire n_6500;
wire n_8135;
wire n_9214;
wire n_13299;
wire n_7051;
wire n_9859;
wire n_11030;
wire n_13394;
wire n_10295;
wire n_5152;
wire n_9003;
wire n_16508;
wire n_11443;
wire n_9271;
wire n_9258;
wire n_6628;
wire n_13849;
wire n_12661;
wire n_12693;
wire n_6297;
wire n_5905;
wire n_12203;
wire n_6975;
wire n_5409;
wire n_8979;
wire n_6329;
wire n_7536;
wire n_12080;
wire n_8529;
wire n_15514;
wire n_10658;
wire n_5688;
wire n_9763;
wire n_16908;
wire n_17087;
wire n_5128;
wire n_10894;
wire n_9597;
wire n_6293;
wire n_8417;
wire n_9965;
wire n_9076;
wire n_10912;
wire n_7952;
wire n_9393;
wire n_8498;
wire n_7991;
wire n_7676;
wire n_11769;
wire n_16052;
wire n_12486;
wire n_7553;
wire n_6905;
wire n_12623;
wire n_7425;
wire n_13698;
wire n_5798;
wire n_6381;
wire n_6521;
wire n_14701;
wire n_5307;
wire n_12933;
wire n_12489;
wire n_8967;
wire n_8355;
wire n_9736;
wire n_13691;
wire n_7998;
wire n_17125;
wire n_14122;
wire n_5986;
wire n_8719;
wire n_16098;
wire n_6581;
wire n_10160;
wire n_10678;
wire n_14372;
wire n_6215;
wire n_7095;
wire n_11794;
wire n_14645;
wire n_15901;
wire n_5415;
wire n_10241;
wire n_5770;
wire n_11495;
wire n_14259;
wire n_7064;
wire n_8762;
wire n_5892;
wire n_12480;
wire n_13273;
wire n_13265;
wire n_17013;
wire n_10180;
wire n_16477;
wire n_8516;
wire n_8880;
wire n_6577;
wire n_6899;
wire n_8784;
wire n_14666;
wire n_12335;
wire n_5676;
wire n_18189;
wire n_7307;
wire n_6545;
wire n_10631;
wire n_8237;
wire n_16974;
wire n_5802;
wire n_13372;
wire n_15897;
wire n_10852;
wire n_14546;
wire n_13669;
wire n_18024;
wire n_18262;
wire n_16469;
wire n_16800;
wire n_18236;
wire n_9803;
wire n_8977;
wire n_13079;
wire n_14371;
wire n_11406;
wire n_8171;
wire n_13121;
wire n_17732;
wire n_10978;
wire n_10500;
wire n_6370;
wire n_9755;
wire n_9805;
wire n_13731;
wire n_15634;
wire n_7210;
wire n_14997;
wire n_7899;
wire n_10370;
wire n_15263;
wire n_15836;
wire n_9728;
wire n_5769;
wire n_6065;
wire n_13845;
wire n_15475;
wire n_16051;
wire n_7039;
wire n_9659;
wire n_6987;
wire n_12624;
wire n_17306;
wire n_14328;
wire n_18134;
wire n_9107;
wire n_18298;
wire n_11428;
wire n_14361;
wire n_6859;
wire n_5331;
wire n_6190;
wire n_16461;
wire n_14311;
wire n_13447;
wire n_12410;
wire n_17846;
wire n_9917;
wire n_14574;
wire n_14847;
wire n_6309;
wire n_11149;
wire n_9520;
wire n_17146;
wire n_6623;
wire n_12055;
wire n_12925;
wire n_7723;
wire n_15922;
wire n_12771;
wire n_6527;
wire n_7443;
wire n_16014;
wire n_13262;
wire n_11707;
wire n_10550;
wire n_18004;
wire n_9583;
wire n_7811;
wire n_12413;
wire n_11086;
wire n_5341;
wire n_12182;
wire n_14096;
wire n_15315;
wire n_14943;
wire n_5930;
wire n_13622;
wire n_5814;
wire n_12803;
wire n_16792;
wire n_9036;
wire n_14007;
wire n_15026;
wire n_9522;
wire n_16709;
wire n_13145;
wire n_16134;
wire n_5979;
wire n_16580;
wire n_14034;
wire n_5271;
wire n_10571;
wire n_5089;
wire n_7015;
wire n_17418;
wire n_5263;
wire n_13276;
wire n_14394;
wire n_11772;
wire n_13338;
wire n_17935;
wire n_14618;
wire n_15806;
wire n_16008;
wire n_12547;
wire n_6929;
wire n_11225;
wire n_11764;
wire n_13904;
wire n_14256;
wire n_16538;
wire n_12544;
wire n_11339;
wire n_5518;
wire n_10125;
wire n_17102;
wire n_5637;
wire n_12370;
wire n_12931;
wire n_14810;
wire n_8279;
wire n_5622;
wire n_13940;
wire n_14054;
wire n_13648;
wire n_14844;
wire n_11112;
wire n_9723;
wire n_12986;
wire n_13570;
wire n_17446;
wire n_7348;
wire n_10254;
wire n_5240;
wire n_5813;
wire n_13543;
wire n_15589;
wire n_5495;
wire n_5546;
wire n_8912;
wire n_13873;
wire n_14491;
wire n_9488;
wire n_7143;
wire n_5482;
wire n_7312;
wire n_5224;
wire n_16548;
wire n_14267;
wire n_7155;
wire n_8227;
wire n_9231;
wire n_8938;
wire n_15116;
wire n_6865;
wire n_16635;
wire n_8787;
wire n_16238;
wire n_16595;
wire n_5393;
wire n_10017;
wire n_6535;
wire n_7213;
wire n_15774;
wire n_14987;
wire n_10866;
wire n_9047;
wire n_10348;
wire n_14846;
wire n_12991;
wire n_8270;
wire n_16724;
wire n_17877;
wire n_5966;
wire n_11072;
wire n_16665;
wire n_17996;
wire n_7456;
wire n_8335;
wire n_11359;
wire n_13449;
wire n_13781;
wire n_13459;
wire n_14974;
wire n_16318;
wire n_10657;
wire n_17656;
wire n_13899;
wire n_7420;
wire n_5041;
wire n_14223;
wire n_11605;
wire n_15871;
wire n_13395;
wire n_9798;
wire n_14463;
wire n_17115;
wire n_9681;
wire n_8054;
wire n_9414;
wire n_16251;
wire n_12419;
wire n_8607;
wire n_5431;
wire n_13760;
wire n_9979;
wire n_9093;
wire n_15677;
wire n_16255;
wire n_14151;
wire n_11959;
wire n_6482;
wire n_15487;
wire n_15609;
wire n_11318;
wire n_11830;
wire n_15428;
wire n_10842;
wire n_15883;
wire n_13012;
wire n_17123;
wire n_15148;
wire n_18042;
wire n_12865;
wire n_8150;
wire n_9379;
wire n_5059;
wire n_5505;
wire n_12009;
wire n_7715;
wire n_9486;
wire n_11881;
wire n_6605;
wire n_9134;
wire n_5329;
wire n_17879;
wire n_15210;
wire n_18209;
wire n_12481;
wire n_7007;
wire n_8358;
wire n_9410;
wire n_16983;
wire n_10045;
wire n_18009;
wire n_14672;
wire n_13594;
wire n_13991;
wire n_15408;
wire n_17576;
wire n_7909;
wire n_14751;
wire n_15133;
wire n_14307;
wire n_9151;
wire n_12278;
wire n_13102;
wire n_14407;
wire n_11863;
wire n_14715;
wire n_15595;
wire n_14563;
wire n_13558;
wire n_18228;
wire n_14428;
wire n_8281;
wire n_12562;
wire n_17028;
wire n_11494;
wire n_9182;
wire n_5908;
wire n_6018;
wire n_16651;
wire n_12744;
wire n_7168;
wire n_11850;
wire n_5212;
wire n_9976;
wire n_7736;
wire n_14107;
wire n_8396;
wire n_9591;
wire n_10322;
wire n_13952;
wire n_9838;
wire n_5939;
wire n_7177;
wire n_10033;
wire n_13027;
wire n_12615;
wire n_14478;
wire n_16429;
wire n_11258;
wire n_10886;
wire n_9568;
wire n_7780;
wire n_17454;
wire n_15956;
wire n_9701;
wire n_9261;
wire n_7379;
wire n_17936;
wire n_7444;
wire n_8223;
wire n_5931;
wire n_11468;
wire n_7435;
wire n_5297;
wire n_7813;
wire n_16278;
wire n_7030;
wire n_8459;
wire n_5420;
wire n_16027;
wire n_17634;
wire n_6311;
wire n_11192;
wire n_12580;
wire n_11569;
wire n_16996;
wire n_6654;
wire n_6424;
wire n_6816;
wire n_6220;
wire n_9752;
wire n_12769;
wire n_5234;
wire n_16744;
wire n_6740;
wire n_7122;
wire n_12540;
wire n_5835;
wire n_7049;
wire n_7567;
wire n_17787;
wire n_16533;
wire n_6029;
wire n_13607;
wire n_18175;
wire n_17626;
wire n_15807;
wire n_13080;
wire n_8379;
wire n_11563;
wire n_15089;
wire n_16340;
wire n_6879;
wire n_13292;
wire n_18128;
wire n_5259;
wire n_16484;
wire n_5440;
wire n_17653;
wire n_5679;
wire n_17448;
wire n_5938;
wire n_9079;
wire n_6702;
wire n_11846;
wire n_16512;
wire n_5891;
wire n_14682;
wire n_10383;
wire n_13377;
wire n_18153;
wire n_5724;
wire n_10064;
wire n_10876;
wire n_5774;
wire n_8793;
wire n_11852;
wire n_6452;
wire n_15637;
wire n_12619;
wire n_14527;
wire n_8975;
wire n_16790;
wire n_14020;
wire n_6791;
wire n_11679;
wire n_9170;
wire n_8792;
wire n_16953;
wire n_5131;
wire n_7280;
wire n_8489;
wire n_8671;
wire n_6915;
wire n_7110;
wire n_7511;
wire n_10831;
wire n_6856;
wire n_7941;
wire n_18232;
wire n_18252;
wire n_7791;
wire n_9385;
wire n_11186;
wire n_11870;
wire n_12960;
wire n_17122;
wire n_13519;
wire n_18040;
wire n_8484;
wire n_8454;
wire n_11492;
wire n_17720;
wire n_13984;
wire n_10536;
wire n_10238;
wire n_7232;
wire n_16519;
wire n_17032;
wire n_8759;
wire n_12268;
wire n_11544;
wire n_7345;
wire n_18182;
wire n_5923;
wire n_8703;
wire n_11233;
wire n_12656;
wire n_15193;
wire n_5790;
wire n_18293;
wire n_16264;
wire n_18233;
wire n_12678;
wire n_14521;
wire n_10206;
wire n_14726;
wire n_16615;
wire n_14924;
wire n_12880;
wire n_9670;
wire n_12876;
wire n_13107;
wire n_6451;
wire n_6364;
wire n_13511;
wire n_12711;
wire n_6552;
wire n_14205;
wire n_15667;
wire n_15168;
wire n_10786;
wire n_8325;
wire n_13523;
wire n_5140;
wire n_6328;
wire n_9598;
wire n_8382;
wire n_7827;
wire n_8971;
wire n_15815;
wire n_6363;
wire n_16281;
wire n_11646;
wire n_10602;
wire n_10620;
wire n_13699;
wire n_14049;
wire n_17657;
wire n_18211;
wire n_16049;
wire n_13420;
wire n_7159;
wire n_8127;
wire n_11878;
wire n_10079;
wire n_10188;
wire n_8721;
wire n_9391;
wire n_15751;
wire n_17510;
wire n_12458;
wire n_6132;
wire n_6578;
wire n_17132;
wire n_8889;
wire n_6406;
wire n_10319;
wire n_17619;
wire n_5598;
wire n_13643;
wire n_13603;
wire n_11900;
wire n_9470;
wire n_18227;
wire n_17860;
wire n_12132;
wire n_14434;
wire n_15429;
wire n_5306;
wire n_16831;
wire n_6978;
wire n_12104;
wire n_16611;
wire n_12467;
wire n_9328;
wire n_12037;
wire n_12870;
wire n_5342;
wire n_9245;
wire n_16156;
wire n_10739;
wire n_12911;
wire n_8232;
wire n_18037;
wire n_7477;
wire n_5147;
wire n_6918;
wire n_12386;
wire n_7363;
wire n_9833;
wire n_11837;
wire n_10213;
wire n_16296;
wire n_18089;
wire n_6612;
wire n_15588;
wire n_10107;
wire n_8664;
wire n_5677;
wire n_10872;
wire n_5997;
wire n_9455;
wire n_12651;
wire n_7863;
wire n_5511;
wire n_9719;
wire n_5680;
wire n_7295;
wire n_8633;
wire n_9744;
wire n_8842;
wire n_15900;
wire n_17531;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_11871;
wire n_8956;
wire n_5280;
wire n_10969;
wire n_6375;
wire n_6479;
wire n_14507;
wire n_17311;
wire n_6866;
wire n_16482;
wire n_16680;
wire n_12563;
wire n_7831;
wire n_13825;
wire n_11674;
wire n_12621;
wire n_5235;
wire n_15234;
wire n_16845;
wire n_13798;
wire n_17620;
wire n_14564;
wire n_12331;
wire n_17648;
wire n_12304;
wire n_9698;
wire n_12339;
wire n_6170;
wire n_12270;
wire n_14599;
wire n_15049;
wire n_9124;
wire n_10718;
wire n_10669;
wire n_9695;
wire n_6447;
wire n_6263;
wire n_7093;
wire n_9497;
wire n_5206;
wire n_10895;
wire n_8641;
wire n_15903;
wire n_8479;
wire n_11610;
wire n_15983;
wire n_17871;
wire n_17949;
wire n_11187;
wire n_12210;
wire n_7466;
wire n_17442;
wire n_14525;
wire n_16735;
wire n_16246;
wire n_14058;
wire n_15249;
wire n_15255;
wire n_5419;
wire n_6130;
wire n_12858;
wire n_14153;
wire n_15101;
wire n_12382;
wire n_11280;
wire n_10757;
wire n_7651;
wire n_13324;
wire n_10513;
wire n_15018;
wire n_5103;
wire n_18301;
wire n_11148;
wire n_8179;
wire n_15825;
wire n_5803;
wire n_13286;
wire n_14272;
wire n_16399;
wire n_6014;
wire n_11396;
wire n_8973;
wire n_16396;
wire n_6935;
wire n_14953;
wire n_10194;
wire n_9775;
wire n_17216;
wire n_7530;
wire n_17636;
wire n_5285;
wire n_11426;
wire n_14980;
wire n_17901;
wire n_9038;
wire n_8308;
wire n_15537;
wire n_18178;
wire n_17394;
wire n_13406;
wire n_5387;
wire n_9630;
wire n_13071;
wire n_16300;
wire n_10692;
wire n_16164;
wire n_8378;
wire n_8733;
wire n_12107;
wire n_14337;
wire n_8809;
wire n_14427;
wire n_5985;
wire n_14439;
wire n_17943;
wire n_11723;
wire n_11009;
wire n_9652;
wire n_10021;
wire n_5058;
wire n_12381;
wire n_6907;
wire n_11706;
wire n_17942;
wire n_13284;
wire n_8500;
wire n_17809;
wire n_12653;
wire n_16820;
wire n_7661;
wire n_6158;
wire n_10782;
wire n_17384;
wire n_9709;
wire n_6541;
wire n_6119;
wire n_8447;
wire n_14202;
wire n_11949;
wire n_5896;
wire n_13303;
wire n_15004;
wire n_10457;
wire n_9324;
wire n_17490;
wire n_13311;
wire n_9934;
wire n_16762;
wire n_13364;
wire n_13813;
wire n_11957;
wire n_5192;
wire n_8548;
wire n_11538;
wire n_5141;
wire n_14743;
wire n_17923;
wire n_5133;
wire n_8412;
wire n_6226;
wire n_11264;
wire n_12774;
wire n_11211;
wire n_17060;
wire n_11880;
wire n_9668;
wire n_14340;
wire n_7145;
wire n_10385;
wire n_15526;
wire n_11377;
wire n_17613;
wire n_12064;
wire n_9877;
wire n_17077;
wire n_12503;
wire n_9657;
wire n_10111;
wire n_11302;
wire n_6338;
wire n_12425;
wire n_14319;
wire n_14922;
wire n_15181;
wire n_11921;
wire n_13358;
wire n_5159;
wire n_15248;
wire n_9352;
wire n_15917;
wire n_9395;
wire n_12807;
wire n_14621;
wire n_15211;
wire n_16367;
wire n_8425;
wire n_10809;
wire n_9349;
wire n_17163;
wire n_18096;
wire n_14734;
wire n_8241;
wire n_7823;
wire n_15268;
wire n_9209;
wire n_7467;
wire n_5097;
wire n_14555;
wire n_10113;
wire n_15010;
wire n_16851;
wire n_18085;
wire n_16485;
wire n_11267;
wire n_10990;
wire n_7932;
wire n_11626;
wire n_14957;
wire n_15308;
wire n_7550;
wire n_5730;
wire n_11694;
wire n_13811;
wire n_14014;
wire n_16109;
wire n_11618;
wire n_9969;
wire n_9937;
wire n_15754;
wire n_5816;
wire n_16359;
wire n_17391;
wire n_7541;
wire n_10545;
wire n_12715;
wire n_17628;
wire n_7241;
wire n_7717;
wire n_18116;
wire n_14945;
wire n_5300;
wire n_10595;
wire n_10973;
wire n_13883;
wire n_11011;
wire n_13814;
wire n_12015;
wire n_12968;
wire n_17956;
wire n_18183;
wire n_9618;
wire n_10732;
wire n_14257;
wire n_10009;
wire n_11776;
wire n_6625;
wire n_17741;
wire n_11165;
wire n_12135;
wire n_7464;
wire n_9082;
wire n_11366;
wire n_17284;
wire n_6302;
wire n_14279;
wire n_17508;
wire n_9424;
wire n_8274;
wire n_9453;
wire n_15239;
wire n_5748;
wire n_13757;
wire n_6759;
wire n_16199;
wire n_5525;
wire n_16699;
wire n_9637;
wire n_8152;
wire n_6706;
wire n_10526;
wire n_8550;
wire n_14190;
wire n_6139;
wire n_14185;
wire n_8264;
wire n_7434;
wire n_7636;
wire n_17086;
wire n_7054;
wire n_6999;
wire n_12817;
wire n_13832;
wire n_6403;
wire n_6483;
wire n_8829;
wire n_9183;
wire n_9205;
wire n_14630;
wire n_13935;
wire n_17698;
wire n_13325;
wire n_9009;
wire n_12869;
wire n_15764;
wire n_17268;
wire n_13841;
wire n_6228;
wire n_11315;
wire n_17234;
wire n_18110;
wire n_5650;
wire n_14104;
wire n_14344;
wire n_10044;
wire n_16181;
wire n_13207;
wire n_12059;
wire n_14188;
wire n_15482;
wire n_16219;
wire n_12586;
wire n_11098;
wire n_5400;
wire n_13043;
wire n_5552;
wire n_7299;
wire n_10221;
wire n_13281;
wire n_6888;
wire n_8266;
wire n_13960;
wire n_15086;
wire n_14069;
wire n_17364;
wire n_8515;
wire n_10109;
wire n_10169;
wire n_17005;
wire n_13556;
wire n_8648;
wire n_17781;
wire n_15707;
wire n_6063;
wire n_10329;
wire n_10928;
wire n_9024;
wire n_9030;
wire n_9523;
wire n_15875;
wire n_9377;
wire n_10891;
wire n_8946;
wire n_15099;
wire n_16074;
wire n_16395;
wire n_10839;
wire n_11875;
wire n_6800;
wire n_5139;
wire n_13260;
wire n_9716;
wire n_6922;
wire n_9380;
wire n_14543;
wire n_6890;
wire n_5481;
wire n_14474;
wire n_8744;
wire n_9000;
wire n_9679;
wire n_9116;
wire n_9742;
wire n_9016;
wire n_7503;
wire n_6070;
wire n_13979;
wire n_13308;
wire n_9006;
wire n_12514;
wire n_13381;
wire n_11524;
wire n_17112;
wire n_10091;
wire n_6651;
wire n_5821;
wire n_7296;
wire n_7091;
wire n_7273;
wire n_6647;
wire n_5733;
wire n_14704;
wire n_10029;
wire n_9690;
wire n_8765;
wire n_15183;
wire n_13483;
wire n_14675;
wire n_5871;
wire n_9852;
wire n_17138;
wire n_16951;
wire n_7543;
wire n_13400;
wire n_10600;
wire n_15424;
wire n_9914;
wire n_17533;
wire n_11056;
wire n_11514;
wire n_12438;
wire n_6184;
wire n_18011;
wire n_14268;
wire n_16157;
wire n_17726;
wire n_11774;
wire n_8627;
wire n_7507;
wire n_9451;
wire n_10849;
wire n_15456;
wire n_15466;
wire n_5043;
wire n_11108;
wire n_9760;
wire n_7555;
wire n_18043;
wire n_15509;
wire n_13910;
wire n_15874;
wire n_5707;
wire n_13907;
wire n_10947;
wire n_17945;
wire n_13369;
wire n_10272;
wire n_12099;
wire n_9035;
wire n_15077;
wire n_12806;
wire n_9211;
wire n_5836;
wire n_18165;
wire n_5281;
wire n_14873;
wire n_6716;
wire n_16043;
wire n_6422;
wire n_12887;
wire n_12776;
wire n_12898;
wire n_17484;
wire n_9677;
wire n_13464;
wire n_5048;
wire n_11954;
wire n_14965;
wire n_5521;
wire n_12191;
wire n_7578;
wire n_13611;
wire n_17632;
wire n_17836;
wire n_7475;
wire n_8195;
wire n_9070;
wire n_5585;
wire n_6397;
wire n_12578;
wire n_17993;
wire n_14012;
wire n_11864;
wire n_14232;
wire n_14221;
wire n_7033;
wire n_9881;
wire n_6121;
wire n_16010;
wire n_9669;
wire n_7531;
wire n_9958;
wire n_9858;
wire n_8462;
wire n_5561;
wire n_9981;
wire n_10391;
wire n_16457;
wire n_8377;
wire n_11157;
wire n_14390;
wire n_17981;
wire n_12509;
wire n_13345;
wire n_12235;
wire n_6981;
wire n_15647;
wire n_18058;
wire n_14932;
wire n_15666;
wire n_9588;
wire n_6954;
wire n_11733;
wire n_5799;
wire n_5073;
wire n_12471;
wire n_13756;
wire n_13632;
wire n_15208;
wire n_17867;
wire n_12365;
wire n_5875;
wire n_8428;
wire n_16734;
wire n_8103;
wire n_13417;
wire n_14350;
wire n_9021;
wire n_17137;
wire n_13130;
wire n_6646;
wire n_8936;
wire n_8414;
wire n_8362;
wire n_15529;
wire n_12083;
wire n_15251;
wire n_9682;
wire n_10137;
wire n_10344;
wire n_7131;
wire n_7769;
wire n_11540;
wire n_10882;
wire n_11861;
wire n_15397;
wire n_17141;
wire n_17388;
wire n_6903;
wire n_9050;
wire n_11724;
wire n_9303;
wire n_14775;
wire n_12065;
wire n_9495;
wire n_13970;
wire n_15156;
wire n_15971;
wire n_12167;
wire n_11220;
wire n_14220;
wire n_6101;
wire n_9415;
wire n_5968;
wire n_14451;
wire n_16426;
wire n_10196;
wire n_8491;
wire n_9058;
wire n_6941;
wire n_9845;
wire n_17778;
wire n_17212;
wire n_8831;
wire n_16506;
wire n_18086;
wire n_18184;
wire n_5812;
wire n_14100;
wire n_6148;
wire n_15704;
wire n_5515;
wire n_8324;
wire n_11459;
wire n_11355;
wire n_6106;
wire n_9822;
wire n_17499;
wire n_12087;
wire n_6604;
wire n_14510;
wire n_17703;
wire n_12243;
wire n_17506;
wire n_7418;
wire n_12267;
wire n_5250;
wire n_12569;
wire n_7688;
wire n_16903;
wire n_17111;
wire n_17965;
wire n_10518;
wire n_11101;
wire n_9640;
wire n_11899;
wire n_8348;
wire n_5607;
wire n_14313;
wire n_15842;
wire n_17777;
wire n_8288;
wire n_10613;
wire n_15688;
wire n_10583;
wire n_14719;
wire n_16420;
wire n_14452;
wire n_15447;
wire n_11481;
wire n_14308;
wire n_16046;
wire n_11712;
wire n_11612;
wire n_8269;
wire n_14288;
wire n_7806;
wire n_10335;
wire n_10085;
wire n_10840;
wire n_6566;
wire n_14833;
wire n_13152;
wire n_18103;
wire n_12599;
wire n_8625;
wire n_5734;
wire n_6081;
wire n_8458;
wire n_16975;
wire n_8806;
wire n_16274;
wire n_13857;
wire n_7204;
wire n_16071;
wire n_10560;
wire n_8180;
wire n_16160;
wire n_8499;
wire n_8601;
wire n_9062;
wire n_13315;
wire n_14606;
wire n_13180;
wire n_14097;
wire n_16666;
wire n_8306;
wire n_5404;
wire n_15510;
wire n_16929;
wire n_12375;
wire n_12091;
wire n_9722;
wire n_12513;
wire n_6047;
wire n_14788;
wire n_8167;
wire n_5438;
wire n_10486;
wire n_9791;
wire n_12307;
wire n_16086;
wire n_18017;
wire n_9229;
wire n_11603;
wire n_11890;
wire n_8613;
wire n_9603;
wire n_11790;
wire n_16967;
wire n_8913;
wire n_11060;
wire n_17345;
wire n_7354;
wire n_7448;
wire n_15550;
wire n_18061;
wire n_8800;
wire n_16047;
wire n_6244;
wire n_17012;
wire n_13474;
wire n_13224;
wire n_16212;
wire n_12684;
wire n_8768;
wire n_6861;
wire n_13702;
wire n_9099;
wire n_10919;
wire n_13797;
wire n_17456;
wire n_14388;
wire n_12288;
wire n_9309;
wire n_12418;
wire n_13853;
wire n_7852;
wire n_13762;
wire n_15957;
wire n_10952;
wire n_5725;
wire n_12566;
wire n_7925;
wire n_12415;
wire n_13037;
wire n_9432;
wire n_16054;
wire n_16849;
wire n_9454;
wire n_7571;
wire n_15351;
wire n_11744;
wire n_13919;
wire n_14466;
wire n_9065;
wire n_11650;
wire n_16547;
wire n_5163;
wire n_11518;
wire n_17881;
wire n_7748;
wire n_5768;
wire n_12949;
wire n_16982;
wire n_7556;
wire n_14061;
wire n_7640;
wire n_8187;
wire n_10352;
wire n_14962;
wire n_15365;
wire n_8881;
wire n_9704;
wire n_15615;
wire n_11663;
wire n_5190;
wire n_7422;
wire n_7920;
wire n_8433;
wire n_9837;
wire n_10991;
wire n_9431;
wire n_10167;
wire n_12681;
wire n_12859;
wire n_14413;
wire n_9160;
wire n_10911;
wire n_17118;
wire n_17979;
wire n_9433;
wire n_14050;
wire n_15587;
wire n_6588;
wire n_17671;
wire n_9256;
wire n_10442;
wire n_12829;
wire n_15179;
wire n_13593;
wire n_11282;
wire n_14912;
wire n_9706;
wire n_12448;
wire n_13044;
wire n_7900;
wire n_7050;
wire n_16976;
wire n_9808;
wire n_13723;
wire n_9915;
wire n_17026;
wire n_10534;
wire n_18242;
wire n_14156;
wire n_5685;
wire n_11726;
wire n_13188;
wire n_5773;
wire n_7136;
wire n_10465;
wire n_10406;
wire n_12188;
wire n_12943;
wire n_8316;
wire n_7318;
wire n_13923;
wire n_16297;
wire n_12149;
wire n_6055;
wire n_5138;
wire n_12783;
wire n_8397;
wire n_9184;
wire n_15136;
wire n_5374;
wire n_17373;
wire n_10373;
wire n_13472;
wire n_9133;
wire n_6108;
wire n_8115;
wire n_12129;
wire n_16353;
wire n_16813;
wire n_12631;
wire n_6165;
wire n_14387;
wire n_10965;
wire n_16694;
wire n_17475;
wire n_6621;
wire n_13148;
wire n_7175;
wire n_5349;
wire n_18099;
wire n_15645;
wire n_7810;
wire n_9109;
wire n_16748;
wire n_13964;
wire n_6323;
wire n_10517;
wire n_17183;
wire n_12588;
wire n_12652;
wire n_8523;
wire n_9207;
wire n_11458;
wire n_13485;
wire n_16855;
wire n_5127;
wire n_17468;
wire n_16727;
wire n_6587;
wire n_16214;
wire n_18330;
wire n_18057;
wire n_6480;
wire n_13531;
wire n_16416;
wire n_13355;
wire n_13368;
wire n_7733;
wire n_6731;
wire n_5485;
wire n_13160;
wire n_16850;
wire n_10484;
wire n_5766;
wire n_11255;
wire n_5216;
wire n_6597;
wire n_13676;
wire n_16004;
wire n_10561;
wire n_13183;
wire n_9673;
wire n_13601;
wire n_15282;
wire n_18097;
wire n_17610;
wire n_8891;
wire n_12523;
wire n_7817;
wire n_11856;
wire n_8294;
wire n_14312;
wire n_16774;
wire n_17838;
wire n_6933;
wire n_7878;
wire n_8338;
wire n_15176;
wire n_15972;
wire n_16411;
wire n_12579;
wire n_16250;
wire n_17952;
wire n_18141;
wire n_9010;
wire n_14904;
wire n_16881;
wire n_8915;
wire n_17466;
wire n_6881;
wire n_11442;
wire n_13052;
wire n_7289;
wire n_14754;
wire n_5805;
wire n_7665;
wire n_17002;
wire n_8131;
wire n_11747;
wire n_9552;
wire n_11008;
wire n_7855;
wire n_13006;
wire n_10371;
wire n_11243;
wire n_12675;
wire n_9841;
wire n_17235;
wire n_12174;
wire n_9230;
wire n_14947;
wire n_14659;
wire n_7764;
wire n_17560;
wire n_15747;
wire n_12113;
wire n_17650;
wire n_12831;
wire n_16960;
wire n_15516;
wire n_10198;
wire n_8027;
wire n_6216;
wire n_10096;
wire n_10582;
wire n_11425;
wire n_10638;
wire n_8162;
wire n_6817;
wire n_7170;
wire n_7314;
wire n_9132;
wire n_11992;
wire n_6949;
wire n_6509;
wire n_14198;
wire n_15882;
wire n_5175;
wire n_7260;
wire n_8855;
wire n_10483;
wire n_11657;
wire n_17000;
wire n_13820;
wire n_12470;
wire n_17976;
wire n_14039;
wire n_8546;
wire n_9878;
wire n_11536;
wire n_11717;
wire n_17584;
wire n_9069;
wire n_8966;
wire n_12154;
wire n_15323;
wire n_8487;
wire n_7263;
wire n_8844;
wire n_14995;
wire n_16312;
wire n_16653;
wire n_5948;
wire n_16570;
wire n_5611;
wire n_10662;
wire n_13471;
wire n_15817;
wire n_16586;
wire n_17992;
wire n_6911;
wire n_9674;
wire n_11512;
wire n_17121;
wire n_11327;
wire n_8533;
wire n_18143;
wire n_12799;
wire n_16438;
wire n_15555;
wire n_13114;
wire n_15002;
wire n_8869;
wire n_5900;
wire n_15860;
wire n_16804;
wire n_14956;
wire n_15731;
wire n_15684;
wire n_9786;
wire n_13976;
wire n_8584;
wire n_6327;
wire n_13200;
wire n_11140;
wire n_8932;
wire n_14862;
wire n_9063;
wire n_8998;
wire n_6607;
wire n_15833;
wire n_9188;
wire n_9467;
wire n_15652;
wire n_9372;
wire n_10960;
wire n_11078;
wire n_9743;
wire n_7850;
wire n_7509;
wire n_16422;
wire n_11620;
wire n_7209;
wire n_5171;
wire n_15592;
wire n_12617;
wire n_6401;
wire n_5554;
wire n_6227;
wire n_12919;
wire n_17260;
wire n_8480;
wire n_9926;
wire n_7240;
wire n_10094;
wire n_12095;
wire n_14620;
wire n_10749;
wire n_17414;
wire n_11907;
wire n_14291;
wire n_15933;
wire n_14092;
wire n_12432;
wire n_12796;
wire n_8911;
wire n_17999;
wire n_11352;
wire n_16591;
wire n_16371;
wire n_5427;
wire n_15876;
wire n_5639;
wire n_14293;
wire n_7725;
wire n_8398;
wire n_10585;
wire n_15039;
wire n_5417;
wire n_8772;
wire n_12279;
wire n_12008;
wire n_9480;
wire n_8307;
wire n_14005;
wire n_14884;
wire n_10896;
wire n_8767;
wire n_16890;
wire n_15273;
wire n_9113;
wire n_9158;
wire n_12156;
wire n_11851;
wire n_13764;
wire n_17217;
wire n_14441;
wire n_16294;
wire n_16545;
wire n_7609;
wire n_14688;
wire n_15827;
wire n_13264;
wire n_8010;
wire n_7278;
wire n_11986;
wire n_12637;
wire n_15878;
wire n_15965;
wire n_17254;
wire n_12301;
wire n_9263;
wire n_18064;
wire n_16959;
wire n_8347;
wire n_17848;
wire n_11734;
wire n_18272;
wire n_7630;
wire n_11517;
wire n_11022;
wire n_14468;
wire n_11831;
wire n_14766;
wire n_10162;
wire n_12302;
wire n_8466;
wire n_6416;
wire n_5488;
wire n_12190;
wire n_14222;
wire n_15054;
wire n_9632;
wire n_17291;
wire n_16370;
wire n_10353;
wire n_17314;
wire n_8813;
wire n_16352;
wire n_8354;
wire n_6695;
wire n_8204;
wire n_14067;
wire n_7741;
wire n_5447;
wire n_5383;
wire n_14598;
wire n_6127;
wire n_7565;
wire n_11259;
wire n_14446;
wire n_11197;
wire n_9282;
wire n_14909;
wire n_14747;
wire n_15635;
wire n_5781;
wire n_15403;
wire n_7883;
wire n_6600;
wire n_10933;
wire n_17171;
wire n_12192;
wire n_7410;
wire n_12010;
wire n_12977;
wire n_10546;
wire n_7097;
wire n_12864;
wire n_13227;
wire n_13869;
wire n_9503;
wire n_6421;
wire n_10724;
wire n_7414;
wire n_5747;
wire n_15486;
wire n_11427;
wire n_10660;
wire n_13348;
wire n_16740;
wire n_16365;
wire n_13166;
wire n_7495;
wire n_9782;
wire n_5969;
wire n_13350;
wire n_9114;
wire n_8312;
wire n_9855;
wire n_15400;
wire n_8040;
wire n_14242;
wire n_11153;
wire n_9347;
wire n_13615;
wire n_9469;
wire n_9680;
wire n_9746;
wire n_10923;
wire n_6079;
wire n_6192;
wire n_9633;
wire n_12746;
wire n_15452;
wire n_10836;
wire n_13266;
wire n_16499;
wire n_6458;
wire n_10884;
wire n_13319;
wire n_13623;
wire n_15062;
wire n_15698;
wire n_8132;
wire n_6746;
wire n_12436;
wire n_7586;
wire n_10780;
wire n_9501;
wire n_12528;
wire n_7720;
wire n_6719;
wire n_13544;
wire n_12792;
wire n_15556;
wire n_16719;
wire n_14586;
wire n_5437;
wire n_9148;
wire n_15417;
wire n_16757;
wire n_15959;
wire n_13530;
wire n_17130;
wire n_11475;
wire n_5826;
wire n_7659;
wire n_17333;
wire n_12973;
wire n_14095;
wire n_11385;
wire n_14191;
wire n_6506;
wire n_14289;
wire n_16588;
wire n_6287;
wire n_13092;
wire n_16354;
wire n_6662;
wire n_17984;
wire n_8650;
wire n_12916;
wire n_10870;
wire n_12923;
wire n_16202;
wire n_9585;
wire n_10267;
wire n_13888;
wire n_8974;
wire n_10379;
wire n_16464;
wire n_17249;
wire n_5245;
wire n_14561;
wire n_7189;
wire n_8688;
wire n_10740;
wire n_10821;
wire n_16891;
wire n_16108;
wire n_17172;
wire n_8983;
wire n_10558;
wire n_6851;
wire n_16450;
wire n_8116;
wire n_12144;
wire n_9338;
wire n_12716;
wire n_6687;
wire n_10297;
wire n_6884;
wire n_8356;
wire n_8013;
wire n_9075;
wire n_13981;
wire n_14614;
wire n_6780;
wire n_6513;
wire n_12463;
wire n_12524;
wire n_16216;
wire n_16928;
wire n_17728;
wire n_8519;
wire n_14484;
wire n_7841;
wire n_15399;
wire n_10497;
wire n_6619;
wire n_10354;
wire n_11456;
wire n_8193;
wire n_17396;
wire n_17072;
wire n_15620;
wire n_14536;
wire n_5603;
wire n_17725;
wire n_10888;
wire n_17883;
wire n_6804;
wire n_9370;
wire n_15717;
wire n_16980;
wire n_11647;
wire n_12392;
wire n_13205;
wire n_13421;
wire n_12173;
wire n_9409;
wire n_17037;
wire n_14140;
wire n_5716;
wire n_16815;
wire n_10138;
wire n_17734;
wire n_18054;
wire n_6516;
wire n_10358;
wire n_5208;
wire n_7490;
wire n_7792;
wire n_10578;
wire n_15902;
wire n_6924;
wire n_13745;
wire n_7492;
wire n_12168;
wire n_12349;
wire n_13349;
wire n_10948;
wire n_5606;
wire n_13730;
wire n_15087;
wire n_12665;
wire n_5231;
wire n_8329;
wire n_5237;
wire n_7809;
wire n_11736;
wire n_14339;
wire n_14804;
wire n_9626;
wire n_14501;
wire n_16073;
wire n_8154;
wire n_15007;
wire n_16812;
wire n_12067;
wire n_17092;
wire n_5456;
wire n_12546;
wire n_7073;
wire n_13489;
wire n_14825;
wire n_11393;
wire n_10007;
wire n_5093;
wire n_10904;
wire n_10386;
wire n_6040;
wire n_15125;
wire n_15479;
wire n_9961;
wire n_13488;
wire n_15542;
wire n_14718;
wire n_5727;
wire n_17643;
wire n_9098;
wire n_11325;
wire n_5390;
wire n_7114;
wire n_5347;
wire n_14612;
wire n_9861;
wire n_6788;
wire n_13638;
wire n_15686;
wire n_17058;
wire n_14869;
wire n_16190;
wire n_11660;
wire n_10448;
wire n_17457;
wire n_14985;
wire n_5115;
wire n_12963;
wire n_14110;
wire n_9536;
wire n_6393;
wire n_8566;
wire n_17878;
wire n_12282;
wire n_8086;
wire n_14316;
wire n_12620;
wire n_8746;
wire n_11411;
wire n_6249;
wire n_14506;
wire n_5833;
wire n_6849;
wire n_13268;
wire n_12431;
wire n_18173;
wire n_18219;
wire n_9593;
wire n_17399;
wire n_18297;
wire n_15613;
wire n_9017;
wire n_5407;
wire n_14595;
wire n_11281;
wire n_15218;
wire n_16874;
wire n_11841;
wire n_11658;
wire n_5232;
wire n_14765;
wire n_18149;
wire n_9703;
wire n_18065;
wire n_14215;
wire n_15437;
wire n_7271;
wire n_12830;
wire n_15991;
wire n_11025;
wire n_6572;
wire n_18125;
wire n_12213;
wire n_6739;
wire n_11372;
wire n_10450;
wire n_13117;
wire n_13510;
wire n_12397;
wire n_14920;
wire n_14781;
wire n_17977;
wire n_13665;
wire n_17190;
wire n_5149;
wire n_7569;
wire n_5151;
wire n_5967;
wire n_7003;
wire n_17572;
wire n_9565;
wire n_7897;
wire n_17160;
wire n_14954;
wire n_7962;
wire n_8942;
wire n_5345;
wire n_5357;
wire n_6666;
wire n_16441;
wire n_13179;
wire n_13429;
wire n_10320;
wire n_17946;
wire n_14835;
wire n_8113;
wire n_6812;
wire n_15284;
wire n_5982;
wire n_10308;
wire n_14216;
wire n_17640;
wire n_17971;
wire n_8652;
wire n_16032;
wire n_13993;
wire n_5135;
wire n_15711;
wire n_17758;
wire n_16092;
wire n_15701;
wire n_7419;
wire n_15025;
wire n_11545;
wire n_12974;
wire n_14078;
wire n_13717;
wire n_5827;
wire n_11465;
wire n_9337;
wire n_5494;
wire n_14314;
wire n_15298;
wire n_15409;
wire n_6200;
wire n_11437;
wire n_15602;
wire n_10304;
wire n_16243;
wire n_11436;
wire n_7784;
wire n_17022;
wire n_13804;
wire n_10902;
wire n_8714;
wire n_6123;
wire n_10607;
wire n_6934;
wire n_7094;
wire n_7500;
wire n_11463;
wire n_14152;
wire n_16320;
wire n_10605;
wire n_11394;
wire n_17081;
wire n_6082;
wire n_10668;
wire n_8944;
wire n_12487;
wire n_13660;
wire n_13861;
wire n_9232;
wire n_12385;
wire n_15471;
wire n_16977;
wire n_17128;
wire n_9320;
wire n_10713;
wire n_16768;
wire n_11191;
wire n_14937;
wire n_17233;
wire n_9167;
wire n_10464;
wire n_5136;
wire n_15451;
wire n_7864;
wire n_5228;
wire n_14580;
wire n_10596;
wire n_14654;
wire n_10034;
wire n_11068;
wire n_15130;
wire n_7129;
wire n_13081;
wire n_5758;
wire n_5323;
wire n_14249;
wire n_7790;
wire n_17884;
wire n_6952;
wire n_17108;
wire n_7062;
wire n_10875;
wire n_15287;
wire n_16166;
wire n_12735;
wire n_9526;
wire n_8107;
wire n_5471;
wire n_7642;
wire n_5434;
wire n_12475;
wire n_15461;
wire n_14300;
wire n_15375;
wire n_9077;
wire n_5941;
wire n_15993;
wire n_16186;
wire n_16794;
wire n_7045;
wire n_12646;
wire n_5879;
wire n_11277;
wire n_15340;
wire n_11665;
wire n_15880;
wire n_15195;
wire n_17458;
wire n_5558;
wire n_11061;
wire n_13800;
wire n_9692;
wire n_13777;
wire n_13444;
wire n_14022;
wire n_5350;
wire n_13267;
wire n_15737;
wire n_13959;
wire n_9141;
wire n_11483;
wire n_5338;
wire n_7238;
wire n_16437;
wire n_12733;
wire n_7126;
wire n_16560;
wire n_9745;
wire n_5669;
wire n_9787;
wire n_8674;
wire n_11073;
wire n_14105;
wire n_12944;
wire n_13362;
wire n_18083;
wire n_14637;
wire n_15120;
wire n_7931;
wire n_10309;
wire n_12061;
wire n_12265;
wire n_13190;
wire n_12380;
wire n_15546;
wire n_8482;
wire n_11462;
wire n_17662;
wire n_8992;
wire n_14703;
wire n_13032;
wire n_6979;
wire n_17199;
wire n_11224;
wire n_10024;
wire n_9892;
wire n_6203;
wire n_7405;
wire n_10762;
wire n_7739;
wire n_16227;
wire n_17231;
wire n_13790;
wire n_10490;
wire n_14357;
wire n_8761;
wire n_9078;
wire n_7207;
wire n_16418;
wire n_8899;
wire n_11127;
wire n_17601;
wire n_7934;
wire n_9015;
wire n_7454;
wire n_14283;
wire n_9012;
wire n_12794;
wire n_5830;
wire n_6796;
wire n_9233;
wire n_12890;
wire n_14492;
wire n_18119;
wire n_9217;
wire n_13576;
wire n_14644;
wire n_5760;
wire n_6368;
wire n_15457;
wire n_6556;
wire n_11632;
wire n_15893;
wire n_10974;
wire n_9435;
wire n_5668;
wire n_17219;
wire n_5878;
wire n_8926;
wire n_5588;
wire n_11692;
wire n_11762;
wire n_14662;
wire n_5765;
wire n_11843;
wire n_14341;
wire n_14470;
wire n_16479;
wire n_17109;
wire n_11344;
wire n_9389;
wire n_11403;
wire n_12926;
wire n_6596;
wire n_15794;
wire n_5090;
wire n_14159;
wire n_6870;
wire n_10520;
wire n_7639;
wire n_13666;
wire n_12247;
wire n_12881;
wire n_5613;
wire n_10914;
wire n_10129;
wire n_16435;
wire n_5104;
wire n_5042;
wire n_13710;
wire n_11510;
wire n_10084;
wire n_14082;
wire n_17711;
wire n_7251;
wire n_15966;
wire n_16193;
wire n_10519;
wire n_7776;
wire n_12966;
wire n_6080;
wire n_10318;
wire n_13785;
wire n_7059;
wire n_13287;
wire n_14665;
wire n_8561;
wire n_10877;
wire n_8255;
wire n_7035;
wire n_10468;
wire n_14752;
wire n_5571;
wire n_11854;
wire n_8029;
wire n_12894;
wire n_10906;
wire n_17493;
wire n_5289;
wire n_6713;
wire n_14632;
wire n_17859;
wire n_5513;
wire n_6747;
wire n_12276;
wire n_6281;
wire n_13588;
wire n_15925;
wire n_17483;
wire n_5972;
wire n_10289;
wire n_14496;
wire n_9381;
wire n_13261;
wire n_13634;
wire n_9873;
wire n_15738;
wire n_16636;
wire n_11925;
wire n_12594;
wire n_10905;
wire n_5916;
wire n_7029;
wire n_5984;
wire n_7317;
wire n_13030;
wire n_14043;
wire n_15855;
wire n_9575;
wire n_5145;
wire n_12529;
wire n_14636;
wire n_11817;
wire n_15887;
wire n_6094;
wire n_15036;
wire n_6444;
wire n_11961;
wire n_12001;
wire n_16941;
wire n_5132;
wire n_15879;
wire n_5191;
wire n_10298;
wire n_12433;
wire n_6333;
wire n_10940;
wire n_6262;
wire n_16103;
wire n_12765;
wire n_13704;
wire n_5869;
wire n_8130;
wire n_5925;
wire n_9023;
wire n_12097;
wire n_6240;
wire n_10723;
wire n_5359;
wire n_13627;
wire n_17325;
wire n_9412;
wire n_6412;
wire n_5293;
wire n_7782;
wire n_7220;
wire n_10293;
wire n_11824;
wire n_15427;
wire n_15228;
wire n_10361;
wire n_7438;
wire n_11269;
wire n_11270;
wire n_9955;
wire n_10161;
wire n_10432;
wire n_15192;
wire n_7515;
wire n_11532;
wire n_7574;
wire n_12402;
wire n_17911;
wire n_12728;
wire n_17357;
wire n_16751;
wire n_16447;
wire n_6684;
wire n_8921;
wire n_13191;
wire n_13784;
wire n_13766;
wire n_10640;
wire n_11546;
wire n_18071;
wire n_7065;
wire n_10271;
wire n_11314;
wire n_5510;
wire n_6046;
wire n_15359;
wire n_7894;
wire n_9418;
wire n_7868;
wire n_16381;
wire n_6973;
wire n_9733;
wire n_14963;
wire n_5363;
wire n_7285;
wire n_17035;
wire n_8286;
wire n_5200;
wire n_9502;
wire n_18164;
wire n_5659;
wire n_5618;
wire n_15045;
wire n_6325;
wire n_15802;
wire n_13374;
wire n_9765;
wire n_9029;
wire n_11130;
wire n_16455;
wire n_10163;
wire n_13824;
wire n_16530;
wire n_6737;
wire n_12262;
wire n_6454;
wire n_5356;
wire n_6721;
wire n_8178;
wire n_14175;
wire n_5369;
wire n_16289;
wire n_11935;
wire n_13452;
wire n_5258;
wire n_12708;
wire n_5255;
wire n_14423;
wire n_15202;
wire n_15919;
wire n_16733;
wire n_18129;
wire n_13656;
wire n_10576;
wire n_9623;
wire n_11822;
wire n_10424;
wire n_12805;
wire n_7008;
wire n_11035;
wire n_8925;
wire n_10404;
wire n_14138;
wire n_16598;
wire n_15318;
wire n_15986;
wire n_8432;
wire n_16040;
wire n_6111;
wire n_16163;
wire n_10130;
wire n_17740;
wire n_12901;
wire n_7505;
wire n_17708;
wire n_8047;
wire n_6260;
wire n_7501;
wire n_17875;
wire n_16515;
wire n_16993;
wire n_10214;
wire n_12971;
wire n_15636;
wire n_5080;
wire n_11389;
wire n_6665;
wire n_9783;
wire n_7566;
wire n_7937;
wire n_12658;
wire n_17766;
wire n_16658;
wire n_7055;
wire n_14568;
wire n_14562;
wire n_12372;
wire n_8268;
wire n_11501;
wire n_12564;
wire n_8053;
wire n_13141;
wire n_17434;
wire n_11015;
wire n_5858;
wire n_16401;
wire n_18274;
wire n_5817;
wire n_10317;
wire n_6690;
wire n_9840;
wire n_5723;
wire n_10491;
wire n_5295;
wire n_6137;
wire n_10712;
wire n_6201;
wire n_10192;
wire n_9909;
wire n_7113;
wire n_12204;
wire n_17287;
wire n_17959;
wire n_14684;
wire n_15055;
wire n_10453;
wire n_11034;
wire n_15852;
wire n_8735;
wire n_11895;
wire n_15291;
wire n_7872;
wire n_12543;
wire n_13895;
wire n_10219;
wire n_15541;
wire n_15722;
wire n_5627;
wire n_16524;
wire n_12888;
wire n_16972;
wire n_13854;
wire n_14062;
wire n_8845;
wire n_7242;
wire n_5155;
wire n_16235;
wire n_14467;
wire n_6461;
wire n_12013;
wire n_8830;
wire n_17098;
wire n_11662;
wire n_17420;
wire n_14706;
wire n_7954;
wire n_6212;
wire n_15703;
wire n_18327;
wire n_6908;
wire n_7819;
wire n_6570;
wire n_15838;
wire n_14362;
wire n_12741;
wire n_8022;
wire n_9532;
wire n_8415;
wire n_9112;
wire n_6498;
wire n_10062;
wire n_16873;
wire n_7228;
wire n_9561;
wire n_6692;
wire n_8547;
wire n_14553;
wire n_16478;
wire n_17930;
wire n_10788;
wire n_11500;
wire n_15092;
wire n_6074;
wire n_10910;
wire n_17229;
wire n_7561;
wire n_6380;
wire n_17709;
wire n_10892;
wire n_17806;
wire n_10216;
wire n_9091;
wire n_14377;
wire n_18290;
wire n_8386;
wire n_5996;
wire n_8426;
wire n_9326;
wire n_8672;
wire n_11977;
wire n_10049;
wire n_5327;
wire n_7994;
wire n_9180;
wire n_10431;
wire n_11215;
wire n_8540;
wire n_6045;
wire n_16737;
wire n_9932;
wire n_15274;
wire n_15421;
wire n_5137;
wire n_6505;
wire n_13705;
wire n_14535;
wire n_15767;
wire n_16097;
wire n_18138;
wire n_14776;
wire n_9220;
wire n_9834;
wire n_17255;
wire n_15814;
wire n_7415;
wire n_13726;
wire n_9474;
wire n_14770;
wire n_14551;
wire n_7793;
wire n_7702;
wire n_5796;
wire n_9542;
wire n_11530;
wire n_7598;
wire n_14406;
wire n_15001;
wire n_6320;
wire n_17465;
wire n_6489;
wire n_6068;
wire n_15000;
wire n_14449;
wire n_12889;
wire n_14290;
wire n_15765;
wire n_14919;
wire n_8192;
wire n_5791;
wire n_17862;
wire n_17366;
wire n_8791;
wire n_17669;
wire n_9458;
wire n_10608;
wire n_15535;
wire n_9642;
wire n_14768;
wire n_5098;
wire n_6877;
wire n_6772;
wire n_9020;
wire n_9910;
wire n_6823;
wire n_6806;
wire n_7426;
wire n_11014;
wire n_15355;
wire n_5906;
wire n_8350;
wire n_11439;
wire n_14744;
wire n_16036;
wire n_12526;
wire n_9100;
wire n_11119;
wire n_11752;
wire n_14081;
wire n_17412;
wire n_14410;
wire n_16944;
wire n_8816;
wire n_7957;
wire n_14549;
wire n_8712;
wire n_16287;
wire n_8048;
wire n_6831;
wire n_17941;
wire n_15058;
wire n_16172;
wire n_10395;
wire n_12255;
wire n_9781;
wire n_13881;
wire n_8663;
wire n_15861;
wire n_7217;
wire n_9940;
wire n_12068;
wire n_10802;
wire n_7058;
wire n_6284;
wire n_6157;
wire n_5423;
wire n_7497;
wire n_18106;
wire n_8503;
wire n_6785;
wire n_8254;
wire n_6374;
wire n_8959;
wire n_13280;
wire n_9117;
wire n_6930;
wire n_12784;
wire n_9198;
wire n_16259;
wire n_6017;
wire n_16623;
wire n_11729;
wire n_8506;
wire n_16624;
wire n_11289;
wire n_11699;
wire n_7735;
wire n_8265;
wire n_8465;
wire n_8049;
wire n_12277;
wire n_16433;
wire n_16821;
wire n_6838;
wire n_11902;
wire n_12212;
wire n_12126;
wire n_5736;
wire n_6937;
wire n_12686;
wire n_15716;
wire n_6443;
wire n_13328;
wire n_6105;
wire n_16236;
wire n_10080;
wire n_16695;
wire n_13554;
wire n_7558;
wire n_12344;
wire n_12250;
wire n_8937;
wire n_12961;
wire n_14142;
wire n_16253;
wire n_17264;
wire n_5069;
wire n_7442;
wire n_10574;
wire n_8272;
wire n_5700;
wire n_6543;
wire n_9249;
wire n_16480;
wire n_15527;
wire n_18281;
wire n_11628;
wire n_10594;
wire n_11784;
wire n_12193;
wire n_16934;
wire n_9398;
wire n_5099;
wire n_16144;
wire n_15748;
wire n_11622;
wire n_14033;
wire n_14269;
wire n_11763;
wire n_13393;
wire n_5052;
wire n_6091;
wire n_17509;
wire n_11606;
wire n_17701;
wire n_12749;
wire n_6674;
wire n_15821;
wire n_18218;
wire n_10155;
wire n_16930;
wire n_17845;
wire n_14585;
wire n_6034;
wire n_16627;
wire n_15683;
wire n_15964;
wire n_15032;
wire n_7499;
wire n_16405;
wire n_17253;
wire n_9751;
wire n_14866;
wire n_13134;
wire n_5579;
wire n_17972;
wire n_8381;
wire n_13399;
wire n_7085;
wire n_16423;
wire n_13413;
wire n_17298;
wire n_12079;
wire n_9579;
wire n_11006;
wire n_10879;
wire n_6652;
wire n_7098;
wire n_6762;
wire n_15090;
wire n_7341;
wire n_7895;
wire n_13602;
wire n_11321;
wire n_13250;
wire n_15980;
wire n_17655;
wire n_17188;
wire n_8366;
wire n_10792;
wire n_16137;
wire n_8101;
wire n_7611;
wire n_16342;
wire n_9925;
wire n_10655;
wire n_14065;
wire n_7391;
wire n_18181;
wire n_17198;
wire n_10890;
wire n_12187;
wire n_16616;
wire n_12093;
wire n_5837;
wire n_14539;
wire n_15963;
wire n_6895;
wire n_7646;
wire n_17276;
wire n_8384;
wire n_13035;
wire n_9889;
wire n_5642;
wire n_14299;
wire n_12705;
wire n_7224;
wire n_5880;
wire n_8728;
wire n_17342;
wire n_6169;
wire n_11133;
wire n_12241;
wire n_14114;
wire n_12211;
wire n_15082;
wire n_17162;
wire n_7524;
wire n_5713;
wire n_6005;
wire n_15100;
wire n_10212;
wire n_8023;
wire n_13770;
wire n_13975;
wire n_17528;
wire n_8052;
wire n_11001;
wire n_7627;
wire n_16391;
wire n_9998;
wire n_11143;
wire n_10654;
wire n_5118;
wire n_5105;
wire n_9729;
wire n_14112;
wire n_15367;
wire n_13833;
wire n_13886;
wire n_15402;
wire n_15934;
wire n_11757;
wire n_13169;
wire n_8614;
wire n_16124;
wire n_5793;
wire n_17855;
wire n_5591;
wire n_13237;
wire n_17367;
wire n_7856;
wire n_16055;
wire n_17716;
wire n_9081;
wire n_7496;
wire n_12446;
wire n_12640;
wire n_15302;
wire n_12699;
wire n_17320;
wire n_9784;
wire n_13354;
wire n_13696;
wire n_15250;
wire n_5623;
wire n_12856;
wire n_14834;
wire n_16106;
wire n_10005;
wire n_17433;
wire n_10544;
wire n_16915;
wire n_10217;
wire n_12231;
wire n_5681;
wire n_11421;
wire n_11780;
wire n_12745;
wire n_14798;
wire n_17760;
wire n_9856;
wire n_15474;
wire n_15768;
wire n_9101;
wire n_7399;
wire n_12841;
wire n_15955;
wire n_8656;
wire n_6213;
wire n_10393;
wire n_6118;
wire n_5256;
wire n_17763;
wire n_11793;
wire n_12527;
wire n_16584;
wire n_18193;
wire n_7605;
wire n_14386;
wire n_11400;
wire n_5220;
wire n_12814;
wire n_5732;
wire n_8897;
wire n_9696;
wire n_12545;
wire n_5178;
wire n_11621;
wire n_15436;
wire n_16380;
wire n_6814;
wire n_13913;
wire n_7342;
wire n_16943;
wire n_12354;
wire n_9825;
wire n_8014;
wire n_13783;
wire n_15493;
wire n_16078;
wire n_5507;
wire n_10093;
wire n_16535;
wire n_18231;
wire n_8564;
wire n_11969;
wire n_14926;
wire n_18023;
wire n_17377;
wire n_7472;
wire n_7214;
wire n_12685;
wire n_5077;
wire n_10850;
wire n_12886;
wire n_13297;
wire n_8371;
wire n_10945;
wire n_5872;
wire n_13564;
wire n_14601;
wire n_15984;
wire n_16679;
wire n_18192;
wire n_11791;
wire n_8231;
wire n_7408;
wire n_9250;
wire n_10541;
wire n_6115;
wire n_9572;
wire n_12196;
wire n_6858;
wire n_10375;
wire n_11948;
wire n_11910;
wire n_8558;
wire n_5735;
wire n_12119;
wire n_9483;
wire n_10275;
wire n_9816;
wire n_17006;
wire n_9253;
wire n_15080;
wire n_8164;
wire n_7254;
wire n_6944;
wire n_7384;
wire n_16981;
wire n_9136;
wire n_14280;
wire n_7837;
wire n_8357;
wire n_10726;
wire n_9426;
wire n_8870;
wire n_9831;
wire n_13434;
wire n_14017;
wire n_14395;
wire n_18171;
wire n_8143;
wire n_11064;
wire n_14187;
wire n_6430;
wire n_14027;
wire n_16510;
wire n_6193;
wire n_17682;
wire n_10614;
wire n_8422;
wire n_6462;
wire n_5314;
wire n_12094;
wire n_15916;
wire n_12096;
wire n_9896;
wire n_9650;
wire n_13657;
wire n_16541;
wire n_12730;
wire n_10002;
wire n_5049;
wire n_6757;
wire n_6822;
wire n_14639;
wire n_5953;
wire n_7599;
wire n_18213;
wire n_16218;
wire n_5277;
wire n_5176;
wire n_11974;
wire n_12202;
wire n_6779;
wire n_6518;
wire n_9767;
wire n_15258;
wire n_16085;
wire n_17772;
wire n_6797;
wire n_11367;
wire n_14094;
wire n_7938;
wire n_8253;
wire n_14730;
wire n_5952;
wire n_15207;
wire n_12534;
wire n_13692;
wire n_5820;
wire n_5483;
wire n_12120;
wire n_16466;
wire n_17488;
wire n_9028;
wire n_9055;
wire n_5718;
wire n_10251;
wire n_14722;
wire n_11562;
wire n_11866;
wire n_13585;
wire n_17159;
wire n_6916;
wire n_17194;
wire n_17951;
wire n_5150;
wire n_11383;
wire n_12854;
wire n_16386;
wire n_16899;
wire n_8563;
wire n_15988;
wire n_9949;
wire n_16168;
wire n_17706;
wire n_5075;
wire n_14906;
wire n_11655;
wire n_12816;
wire n_7812;
wire n_12553;
wire n_18319;
wire n_5051;
wire n_16907;
wire n_18331;
wire n_14486;
wire n_11552;
wire n_14807;
wire n_18259;
wire n_9684;
wire n_15418;
wire n_6152;
wire n_10010;
wire n_9724;
wire n_13430;
wire n_8243;
wire n_10226;
wire n_11117;
wire n_14964;
wire n_8236;
wire n_11046;
wire n_8292;
wire n_17614;
wire n_14640;
wire n_18279;
wire n_14901;
wire n_11547;
wire n_12676;
wire n_13327;
wire n_14412;
wire n_14391;
wire n_5777;
wire n_7949;
wire n_18113;
wire n_8611;
wire n_7046;
wire n_12720;
wire n_17361;
wire n_16760;
wire n_10475;
wire n_13365;
wire n_10020;
wire n_9826;
wire n_5142;
wire n_14195;
wire n_10467;
wire n_18072;
wire n_5156;
wire n_13118;
wire n_5926;
wire n_8011;
wire n_15271;
wire n_9839;
wire n_15816;
wire n_14431;
wire n_9399;
wire n_12535;
wire n_14254;
wire n_13279;
wire n_15497;
wire n_17393;
wire n_17544;
wire n_17522;
wire n_12283;
wire n_12506;
wire n_14044;
wire n_16678;
wire n_6589;
wire n_17672;
wire n_7579;
wire n_16424;
wire n_15393;
wire n_8139;
wire n_12046;
wire n_8123;
wire n_15104;
wire n_10720;
wire n_7173;
wire n_7917;
wire n_5951;
wire n_7092;
wire n_10907;
wire n_6197;
wire n_6971;
wire n_9938;
wire n_8424;
wire n_9776;
wire n_8859;
wire n_13844;
wire n_14462;
wire n_11256;
wire n_7460;
wire n_9658;
wire n_15773;
wire n_16539;
wire n_11914;
wire n_9605;
wire n_12124;
wire n_11934;
wire n_14731;
wire n_15638;
wire n_11047;
wire n_10868;
wire n_17872;
wire n_17829;
wire n_9013;
wire n_8730;
wire n_9417;
wire n_14004;
wire n_13945;
wire n_14841;
wire n_8156;
wire n_9290;
wire n_9212;
wire n_13431;
wire n_15446;
wire n_13342;
wire n_9721;
wire n_14913;
wire n_14789;
wire n_12189;
wire n_10615;
wire n_7698;
wire n_12884;
wire n_13187;
wire n_7886;
wire n_7344;
wire n_6154;
wire n_14504;
wire n_6020;
wire n_15884;
wire n_13082;
wire n_9586;
wire n_7904;
wire n_12310;
wire n_11004;
wire n_10751;
wire n_12683;
wire n_16728;
wire n_13821;
wire n_11287;
wire n_5701;
wire n_10706;
wire n_18142;
wire n_10774;
wire n_11208;
wire n_16467;
wire n_12108;
wire n_12502;
wire n_15267;
wire n_9104;
wire n_7079;
wire n_10225;
wire n_11963;
wire n_10570;
wire n_9293;
wire n_15517;
wire n_16987;
wire n_11860;
wire n_13298;
wire n_5120;
wire n_8645;
wire n_10744;
wire n_16504;
wire n_11625;
wire n_5470;
wire n_17135;
wire n_17595;
wire n_17970;
wire n_16174;
wire n_7675;
wire n_10416;
wire n_16949;
wire n_14933;
wire n_7774;
wire n_17511;
wire n_5797;
wire n_7922;
wire n_8189;
wire n_8618;
wire n_6696;
wire n_11181;
wire n_11787;
wire n_14024;
wire n_5222;
wire n_13810;
wire n_8285;
wire n_17736;
wire n_5743;
wire n_9919;
wire n_10396;
wire n_12899;
wire n_8826;
wire n_6210;
wire n_10123;
wire n_5772;
wire n_14252;
wire n_15790;
wire n_17225;
wire n_8715;
wire n_12761;
wire n_17898;
wire n_14522;
wire n_8782;
wire n_6964;
wire n_14399;
wire n_10083;
wire n_5801;
wire n_6117;
wire n_14331;
wire n_15561;
wire n_8117;
wire n_12918;
wire n_11825;
wire n_17961;
wire n_6202;
wire n_7279;
wire n_7670;
wire n_11364;
wire n_12713;
wire n_15585;
wire n_14126;
wire n_12522;
wire n_12822;
wire n_9445;
wire n_14148;
wire n_18261;
wire n_14031;
wire n_6681;
wire n_13539;
wire n_5971;
wire n_11420;
wire n_12223;
wire n_13532;
wire n_15892;
wire n_11470;
wire n_13089;
wire n_5392;
wire n_8497;
wire n_12082;
wire n_9930;
wire n_6661;
wire n_8018;
wire n_6640;
wire n_12151;
wire n_17278;
wire n_15755;
wire n_17038;
wire n_13335;
wire n_7940;
wire n_14493;
wire n_11230;
wire n_12757;
wire n_7371;
wire n_10731;
wire n_6962;
wire n_13411;
wire n_11063;
wire n_10347;
wire n_11074;
wire n_15468;
wire n_6455;
wire n_17783;
wire n_7721;
wire n_9727;
wire n_17459;
wire n_15034;
wire n_7606;
wire n_16965;
wire n_18159;
wire n_18050;
wire n_5443;
wire n_12025;
wire n_5600;
wire n_15895;
wire n_5169;
wire n_6963;
wire n_10926;
wire n_6644;
wire n_13879;
wire n_13848;
wire n_14534;
wire n_6896;
wire n_14475;
wire n_12183;
wire n_14633;
wire n_17110;
wire n_11669;
wire n_16712;
wire n_10734;
wire n_6832;
wire n_8798;
wire n_7836;
wire n_16823;
wire n_16128;
wire n_16224;
wire n_17174;
wire n_12143;
wire n_6160;
wire n_14473;
wire n_7564;
wire n_11493;
wire n_12158;
wire n_7884;
wire n_8673;
wire n_10281;
wire n_17668;
wire n_6718;
wire n_9685;
wire n_11486;
wire n_8502;
wire n_6542;
wire n_10126;
wire n_10759;
wire n_13293;
wire n_11786;
wire n_17295;
wire n_10650;
wire n_14083;
wire n_16465;
wire n_17906;
wire n_11777;
wire n_6031;
wire n_5502;
wire n_5568;
wire n_9421;
wire n_8577;
wire n_11722;
wire n_14487;
wire n_7653;
wire n_15835;
wire n_16667;
wire n_10092;
wire n_10445;
wire n_15241;
wire n_5656;
wire n_8531;
wire n_16858;
wire n_8635;
wire n_6763;
wire n_5974;
wire n_9567;
wire n_6280;
wire n_9298;
wire n_11941;
wire n_10116;
wire n_6438;
wire n_13614;
wire n_10048;
wire n_9059;
wire n_12937;
wire n_15372;
wire n_8485;
wire n_17352;
wire n_13285;
wire n_6316;
wire n_7383;
wire n_18315;
wire n_18031;
wire n_5474;
wire n_13596;
wire n_8872;
wire n_8752;
wire n_16711;
wire n_18214;
wire n_13609;
wire n_9396;
wire n_17504;
wire n_5413;
wire n_6758;
wire n_12459;
wire n_13715;
wire n_13398;
wire n_7976;
wire n_9234;
wire n_9425;
wire n_12648;
wire n_10364;
wire n_5412;
wire n_17170;
wire n_17402;
wire n_9620;
wire n_6069;
wire n_10963;
wire n_5752;
wire n_10191;
wire n_6874;
wire n_17824;
wire n_13330;
wire n_16127;
wire n_13235;
wire n_15319;
wire n_8341;
wire n_13412;
wire n_13995;
wire n_14867;
wire n_12638;
wire n_16263;
wire n_8521;
wire n_11209;
wire n_6030;
wire n_13561;
wire n_8199;
wire n_12976;
wire n_13091;
wire n_13306;
wire n_18222;
wire n_6077;
wire n_16270;
wire n_17869;
wire n_8005;
wire n_11718;
wire n_7743;
wire n_16961;
wire n_16122;
wire n_17168;
wire n_5201;
wire n_6299;
wire n_9280;
wire n_9517;
wire n_6386;
wire n_9639;
wire n_9192;
wire n_14089;
wire n_12762;
wire n_9102;
wire n_5217;
wire n_10003;
wire n_10025;
wire n_8016;
wire n_10156;
wire n_8669;
wire n_17605;
wire n_5957;
wire n_15603;
wire n_12066;
wire n_11234;
wire n_16101;
wire n_12021;
wire n_14822;
wire n_8283;
wire n_13016;
wire n_13048;
wire n_17804;
wire n_10502;
wire n_16102;
wire n_7655;
wire n_5490;
wire n_8291;
wire n_17209;
wire n_17323;
wire n_16377;
wire n_8176;
wire n_10674;
wire n_16721;
wire n_17334;
wire n_17129;
wire n_15337;
wire n_5158;
wire n_14942;
wire n_6708;
wire n_7737;
wire n_16696;
wire n_10179;
wire n_16470;
wire n_14076;
wire n_7433;
wire n_11000;
wire n_12447;
wire n_13939;
wire n_16856;
wire n_11702;
wire n_10466;
wire n_12667;
wire n_16273;
wire n_15782;
wire n_12221;
wire n_7347;
wire n_8145;
wire n_9487;
wire n_10268;
wire n_13560;
wire n_6792;
wire n_14389;
wire n_12906;
wire n_15392;
wire n_7633;
wire n_12851;
wire n_6177;
wire n_5912;
wire n_11431;
wire n_10679;
wire n_12691;
wire n_7798;
wire n_10492;
wire n_11177;
wire n_12980;
wire n_12416;
wire n_16284;
wire n_17699;
wire n_13436;
wire n_17842;
wire n_13023;
wire n_13985;
wire n_11454;
wire n_9221;
wire n_6033;
wire n_12989;
wire n_11418;
wire n_18161;
wire n_7397;
wire n_5557;
wire n_12739;
wire n_7389;
wire n_13074;
wire n_12791;
wire n_5472;
wire n_16860;
wire n_7602;
wire n_13920;
wire n_13795;
wire n_14483;
wire n_8069;
wire n_6002;
wire n_14696;
wire n_14571;
wire n_17018;
wire n_14753;
wire n_5711;
wire n_7554;
wire n_18118;
wire n_16471;
wire n_14903;
wire n_5396;
wire n_7693;
wire n_14052;
wire n_16562;
wire n_5335;
wire n_8888;
wire n_12650;
wire n_12319;
wire n_15661;
wire n_15391;
wire n_6557;
wire n_7300;
wire n_17503;
wire n_18013;
wire n_15515;
wire n_9566;
wire n_17550;
wire n_12692;
wire n_12403;
wire n_14908;
wire n_17426;
wire n_15522;
wire n_9578;
wire n_8483;
wire n_15534;
wire n_14820;
wire n_8797;
wire n_5960;
wire n_8605;
wire n_8041;
wire n_18122;
wire n_18325;
wire n_9868;
wire n_13451;
wire n_18014;
wire n_14778;
wire n_15225;
wire n_11750;
wire n_14124;
wire n_18249;
wire n_14442;
wire n_15386;
wire n_11572;
wire n_18238;
wire n_7532;
wire n_11038;
wire n_11049;
wire n_9292;
wire n_10460;
wire n_13363;
wire n_5143;
wire n_7724;
wire n_18002;
wire n_12669;
wire n_15492;
wire n_15508;
wire n_11491;
wire n_14838;
wire n_6142;
wire n_6917;
wire n_7510;
wire n_11109;
wire n_5859;
wire n_16833;
wire n_10968;
wire n_8760;
wire n_10004;
wire n_8928;
wire n_11894;
wire n_10729;
wire n_16305;
wire n_17558;
wire n_13689;
wire n_8374;
wire n_17076;
wire n_14276;
wire n_8917;
wire n_6163;
wire n_10811;
wire n_14540;
wire n_7118;
wire n_16509;
wire n_8006;
wire n_11806;
wire n_17680;
wire n_9884;
wire n_11504;
wire n_11737;
wire n_6778;
wire n_7946;
wire n_8723;
wire n_6285;
wire n_9857;
wire n_12127;
wire n_11637;
wire n_14622;
wire n_6025;
wire n_13769;
wire n_8957;
wire n_12058;
wire n_7257;
wire n_11799;
wire n_10944;
wire n_11788;
wire n_13537;
wire n_16999;
wire n_17395;
wire n_15809;
wire n_16521;
wire n_6862;
wire n_7067;
wire n_6319;
wire n_13143;
wire n_13808;
wire n_10140;
wire n_12868;
wire n_14226;
wire n_17774;
wire n_12642;
wire n_10013;
wire n_14106;
wire n_17073;
wire n_12600;
wire n_7933;
wire n_5283;
wire n_8409;
wire n_9815;
wire n_9110;
wire n_7669;
wire n_5268;
wire n_10110;
wire n_13909;
wire n_6318;
wire n_10133;
wire n_14531;
wire n_14720;
wire n_17126;
wire n_8215;
wire n_11453;
wire n_16234;
wire n_11184;
wire n_8220;
wire n_9471;
wire n_9048;
wire n_7927;
wire n_11356;
wire n_6089;
wire n_18052;
wire n_8629;
wire n_13045;
wire n_5122;
wire n_7910;
wire n_11955;
wire n_12005;
wire n_13426;
wire n_14596;
wire n_6315;
wire n_10592;
wire n_14887;
wire n_7970;
wire n_14172;
wire n_15518;
wire n_15985;
wire n_10476;
wire n_8407;
wire n_5556;
wire n_5462;
wire n_16100;
wire n_15153;
wire n_14147;
wire n_12953;
wire n_14593;
wire n_13507;
wire n_15159;
wire n_11488;
wire n_13040;
wire n_18280;
wire n_17622;
wire n_15432;
wire n_12369;
wire n_9394;
wire n_8991;
wire n_12300;
wire n_5840;
wire n_13015;
wire n_14934;
wire n_6343;
wire n_10186;
wire n_11938;
wire n_17100;
wire n_15505;
wire n_14988;
wire n_11946;
wire n_17538;
wire n_9191;
wire n_11918;
wire n_16404;
wire n_17557;
wire n_18205;
wire n_9004;
wire n_12832;
wire n_13839;
wire n_6049;
wire n_6919;
wire n_7423;
wire n_17773;
wire n_17673;
wire n_7865;
wire n_6052;
wire n_17565;
wire n_11412;
wire n_13522;
wire n_10700;
wire n_5330;
wire n_15690;
wire n_15746;
wire n_7069;
wire n_12290;
wire n_13208;
wire n_6886;
wire n_13761;
wire n_18295;
wire n_14219;
wire n_12169;
wire n_8783;
wire n_6912;
wire n_8326;
wire n_10496;
wire n_11249;
wire n_13538;
wire n_10521;
wire n_12838;
wire n_5914;
wire n_14523;
wire n_11464;
wire n_12325;
wire n_15465;
wire n_8504;
wire n_10695;
wire n_14763;
wire n_8445;
wire n_11950;
wire n_13847;
wire n_11648;
wire n_8250;
wire n_18283;
wire n_10994;
wire n_11576;
wire n_5039;
wire n_9118;
wire n_13950;
wire n_6061;
wire n_14025;
wire n_15006;
wire n_12969;
wire n_13214;
wire n_5378;
wire n_10758;
wire n_13559;
wire n_8408;
wire n_10120;
wire n_11410;
wire n_15499;
wire n_11251;
wire n_7252;
wire n_17411;
wire n_5542;
wire n_15450;
wire n_9051;
wire n_16159;
wire n_17241;
wire n_7133;
wire n_6883;
wire n_10345;
wire n_13065;
wire n_5519;
wire n_12809;
wire n_9908;
wire n_12748;
wire n_17095;
wire n_18123;
wire n_13639;
wire n_16691;
wire n_6009;
wire n_7061;
wire n_8155;
wire n_5278;
wire n_8818;
wire n_12264;
wire n_11633;
wire n_11641;
wire n_16592;
wire n_16840;
wire n_17372;
wire n_7518;
wire n_9123;
wire n_12352;
wire n_17041;
wire n_5586;
wire n_13221;
wire n_15297;
wire n_10232;
wire n_17182;
wire n_6378;
wire n_8660;
wire n_5187;
wire n_13619;
wire n_15581;
wire n_12054;
wire n_5675;
wire n_14055;
wire n_18202;
wire n_8275;
wire n_9327;
wire n_6601;
wire n_5771;
wire n_7216;
wire n_6407;
wire n_15488;
wire n_11555;
wire n_9687;
wire n_14552;
wire n_17222;
wire n_8297;
wire n_9828;
wire n_6749;
wire n_13921;
wire n_11984;
wire n_14355;
wire n_6839;
wire n_10533;
wire n_13053;
wire n_14448;
wire n_9519;
wire n_10611;
wire n_7711;
wire n_15431;
wire n_13635;
wire n_12368;
wire n_10089;
wire n_15206;
wire n_12137;
wire n_15538;
wire n_17569;
wire n_11651;
wire n_14038;
wire n_7705;
wire n_10455;
wire n_15259;
wire n_8590;
wire n_6051;
wire n_12538;
wire n_6217;
wire n_13671;
wire n_6680;
wire n_5844;
wire n_12016;
wire n_15610;
wire n_7972;
wire n_16537;
wire n_17602;
wire n_15075;
wire n_6532;
wire n_13517;
wire n_15837;
wire n_17815;
wire n_6155;
wire n_17817;
wire n_6446;
wire n_8072;
wire n_12644;
wire n_17187;
wire n_6738;
wire n_6250;
wire n_7458;
wire n_7614;
wire n_7854;
wire n_12017;
wire n_7707;
wire n_10632;
wire n_13428;
wire n_17422;
wire n_11672;
wire n_16016;
wire n_11696;
wire n_8050;
wire n_6736;
wire n_5344;
wire n_16730;
wire n_15398;
wire n_6526;
wire n_8142;
wire n_10820;
wire n_14914;
wire n_10601;
wire n_13455;
wire n_6339;
wire n_17451;
wire n_14594;
wire n_17424;
wire n_12197;
wire n_5225;
wire n_8151;
wire n_6350;
wire n_7013;
wire n_12892;
wire n_5662;
wire n_17371;
wire n_16061;
wire n_14213;
wire n_9802;
wire n_9315;
wire n_9296;
wire n_8599;
wire n_10447;
wire n_12373;
wire n_12660;
wire n_14393;
wire n_10022;
wire n_14526;
wire n_15278;
wire n_18263;
wire n_5265;
wire n_14184;
wire n_11567;
wire n_10305;
wire n_14769;
wire n_12855;
wire n_17211;
wire n_15777;
wire n_14795;
wire n_16880;
wire n_10031;
wire n_12877;
wire n_5705;
wire n_12350;
wire n_14691;
wire n_15730;
wire n_14576;
wire n_15944;
wire n_13137;
wire n_10798;
wire n_12388;
wire n_7656;
wire n_10760;
wire n_11202;
wire n_6845;
wire n_9405;
wire n_14647;
wire n_12891;
wire n_9302;
wire n_7105;
wire n_18264;
wire n_12836;
wire n_5196;
wire n_13892;
wire n_16298;
wire n_5181;
wire n_17313;
wire n_13636;
wire n_16057;
wire n_11779;
wire n_11888;
wire n_10166;
wire n_14317;
wire n_16489;
wire n_15024;
wire n_6829;
wire n_11684;
wire n_11879;
wire n_16866;
wire n_5574;
wire n_15843;
wire n_11054;
wire n_16272;
wire n_5126;
wire n_6508;
wire n_9977;
wire n_9842;
wire n_9887;
wire n_15820;
wire n_14893;
wire n_15370;
wire n_7570;
wire n_5553;
wire n_11116;
wire n_8246;
wire n_15220;
wire n_9524;
wire n_16346;
wire n_11129;
wire n_7771;
wire n_13742;
wire n_7052;
wire n_7262;
wire n_5368;
wire n_9322;
wire n_11937;
wire n_17793;
wire n_10098;
wire n_15079;
wire n_10510;
wire n_13934;
wire n_13905;
wire n_10848;
wire n_10042;
wire n_8057;
wire n_9122;
wire n_8349;
wire n_5626;
wire n_9333;
wire n_13240;
wire n_16131;
wire n_15947;
wire n_8743;
wire n_6603;
wire n_6114;
wire n_14073;
wire n_16136;
wire n_9590;
wire n_13515;
wire n_6576;
wire n_15915;
wire n_17097;
wire n_7943;
wire n_17590;
wire n_18032;
wire n_7364;
wire n_8473;
wire n_10993;
wire n_13838;
wire n_10342;
wire n_7208;
wire n_12286;
wire n_6245;
wire n_15353;
wire n_12992;
wire n_14132;
wire n_10439;
wire n_16918;
wire n_11923;
wire n_12844;
wire n_14284;
wire n_5499;
wire n_6703;
wire n_18287;
wire n_5604;
wire n_13868;
wire n_9676;
wire n_15103;
wire n_10444;
wire n_7714;
wire n_10054;
wire n_9902;
wire n_17966;
wire n_12759;
wire n_16430;
wire n_8535;
wire n_17627;
wire n_16726;
wire n_10728;
wire n_17537;
wire n_9621;
wire n_13175;
wire n_7202;
wire n_9140;
wire n_9604;
wire n_18144;
wire n_7011;
wire n_18194;
wire n_13759;
wire n_7621;
wire n_5291;
wire n_8068;
wire n_10565;
wire n_10540;
wire n_14444;
wire n_12935;
wire n_16230;
wire n_9821;
wire n_11943;
wire n_14158;
wire n_10748;
wire n_5876;
wire n_17042;
wire n_10178;
wire n_11995;
wire n_15294;
wire n_11058;
wire n_16955;
wire n_17270;
wire n_6970;
wire n_11842;
wire n_12076;
wire n_12790;
wire n_12979;
wire n_5114;
wire n_6704;
wire n_6409;
wire n_16191;
wire n_6876;
wire n_12659;
wire n_7778;
wire n_9343;
wire n_15563;
wire n_7028;
wire n_12532;
wire n_7320;
wire n_7313;
wire n_6255;
wire n_14437;
wire n_7343;
wire n_5288;
wire n_5540;
wire n_5699;
wire n_11473;
wire n_7525;
wire n_13735;
wire n_7875;
wire n_16065;
wire n_5810;
wire n_11568;
wire n_14384;
wire n_16113;
wire n_13258;
wire n_15784;
wire n_15891;
wire n_13617;
wire n_12702;
wire n_16077;
wire n_17207;
wire n_16350;
wire n_17715;
wire n_6938;
wire n_12050;
wire n_12138;
wire n_5762;
wire n_16672;
wire n_16705;
wire n_13713;
wire n_5218;
wire n_8785;
wire n_9952;
wire n_12473;
wire n_13013;
wire n_14577;
wire n_15175;
wire n_10686;
wire n_15975;
wire n_8327;
wire n_12606;
wire n_9219;
wire n_7337;
wire n_6989;
wire n_8512;
wire n_13625;
wire n_5408;
wire n_10971;
wire n_6427;
wire n_15810;
wire n_13051;
wire n_13054;
wire n_7753;
wire n_10076;
wire n_11924;
wire n_15410;
wire n_12374;
wire n_8168;
wire n_14837;
wire n_16099;
wire n_14266;
wire n_14064;
wire n_8392;
wire n_17043;
wire n_7038;
wire n_12967;
wire n_15440;
wire n_14745;
wire n_15383;
wire n_5366;
wire n_17702;
wire n_10132;
wire n_10282;
wire n_13649;
wire n_9872;
wire n_16080;
wire n_15354;
wire n_12956;
wire n_6360;
wire n_18145;
wire n_11203;
wire n_18314;
wire n_13026;
wire n_18020;
wire n_9553;
wire n_10900;
wire n_6146;
wire n_10616;
wire n_18248;
wire n_9447;
wire n_6270;
wire n_11585;
wire n_9150;
wire n_17674;
wire n_18190;
wire n_16717;
wire n_5477;
wire n_9592;
wire n_9984;
wire n_5451;
wire n_12695;
wire n_14111;
wire n_11416;
wire n_17398;
wire n_11526;
wire n_11742;
wire n_13855;
wire n_12179;
wire n_18067;
wire n_8419;
wire n_16280;
wire n_11809;
wire n_15187;
wire n_5086;
wire n_9814;
wire n_10858;
wire n_12038;
wire n_17535;
wire n_5901;
wire n_6353;
wire n_16989;
wire n_14359;
wire n_17530;
wire n_10769;
wire n_15513;
wire n_16739;
wire n_9446;
wire n_14689;
wire n_17513;
wire n_15088;
wire n_17733;
wire n_10211;
wire n_10023;
wire n_15335;
wire n_11877;
wire n_15384;
wire n_17841;
wire n_6345;
wire n_12105;
wire n_9461;
wire n_16336;
wire n_10772;
wire n_9793;
wire n_6691;
wire n_8997;
wire n_14324;
wire n_16895;
wire n_17571;
wire n_15939;
wire n_13184;
wire n_15641;
wire n_12360;
wire n_15330;
wire n_15361;
wire n_12297;
wire n_12952;
wire n_9874;
wire n_13332;
wire n_7392;
wire n_5053;
wire n_7912;
wire n_8245;
wire n_14567;
wire n_6239;
wire n_6803;
wire n_16931;
wire n_10446;
wire n_11735;
wire n_14981;
wire n_7919;
wire n_15050;
wire n_6340;
wire n_7583;
wire n_14281;
wire n_14876;
wire n_8109;
wire n_5226;
wire n_7657;
wire n_14129;
wire n_15936;
wire n_17505;
wire n_7995;
wire n_11405;
wire n_15382;
wire n_5867;
wire n_8985;
wire n_6048;
wire n_13318;
wire n_18098;
wire n_14733;
wire n_5079;
wire n_5590;
wire n_16994;
wire n_10331;
wire n_12103;
wire n_6773;
wire n_9403;
wire n_5632;
wire n_14515;
wire n_8390;
wire n_15252;
wire n_11480;
wire n_17840;
wire n_16268;
wire n_11874;
wire n_12115;
wire n_6336;
wire n_8463;
wire n_14120;
wire n_7041;
wire n_15324;
wire n_17096;
wire n_7802;
wire n_15489;
wire n_14243;
wire n_7370;
wire n_13366;
wire n_10181;
wire n_10074;
wire n_9731;
wire n_5660;
wire n_11104;
wire n_17988;
wire n_13677;
wire n_7557;
wire n_11862;
wire n_16885;
wire n_11952;
wire n_14529;
wire n_6174;
wire n_12828;
wire n_13322;
wire n_6023;
wire n_18299;
wire n_6776;
wire n_18300;
wire n_14894;
wire n_18038;
wire n_13078;
wire n_5426;
wire n_18077;
wire n_17730;
wire n_15496;
wire n_9947;
wire n_15758;
wire n_6463;
wire n_15423;
wire n_13387;
wire n_14370;
wire n_7896;
wire n_16836;
wire n_13226;
wire n_9699;
wire n_6372;
wire n_10962;
wire n_11037;
wire n_9305;
wire n_10481;
wire n_14624;
wire n_7176;
wire n_12003;
wire n_14194;
wire n_14868;
wire n_15770;
wire n_18270;
wire n_10220;
wire n_13917;
wire n_17324;
wire n_10381;
wire n_15237;
wire n_8517;
wire n_12332;
wire n_5625;
wire n_5778;
wire n_6396;
wire n_10642;
wire n_9218;
wire n_13317;
wire n_11556;
wire n_17816;
wire n_6669;
wire n_9096;
wire n_10634;
wire n_13480;
wire n_17541;
wire n_10170;
wire n_10142;
wire n_10569;
wire n_12326;
wire n_15449;
wire n_14489;
wire n_15830;
wire n_5531;
wire n_15321;
wire n_16867;
wire n_9534;
wire n_7826;
wire n_18203;
wire n_18021;
wire n_5429;
wire n_11044;
wire n_5818;
wire n_5646;
wire n_6940;
wire n_5248;
wire n_11042;
wire n_17404;
wire n_12141;
wire n_6394;
wire n_9164;
wire n_9546;
wire n_12622;
wire n_11226;
wire n_5448;
wire n_7590;
wire n_5432;
wire n_14977;
wire n_16126;
wire n_13732;
wire n_15804;
wire n_9358;
wire n_11985;
wire n_16606;
wire n_5160;
wire n_11328;
wire n_13545;
wire n_16756;
wire n_8208;
wire n_15117;
wire n_6995;
wire n_7185;
wire n_10127;
wire n_14214;
wire n_11525;
wire n_16472;
wire n_9730;
wire n_6254;
wire n_6161;
wire n_13246;
wire n_9066;
wire n_16209;
wire n_10800;
wire n_11020;
wire n_9185;
wire n_15233;
wire n_17768;
wire n_16444;
wire n_9318;
wire n_18112;
wire n_10374;
wire n_7987;
wire n_8134;
wire n_14367;
wire n_10328;
wire n_14542;
wire n_8631;
wire n_5445;
wire n_8694;
wire n_11892;
wire n_8965;
wire n_16550;
wire n_8647;
wire n_13288;
wire n_11013;
wire n_17704;
wire n_12343;
wire n_7332;
wire n_6660;
wire n_15396;
wire n_5719;
wire n_17598;
wire n_15422;
wire n_7225;
wire n_10529;
wire n_12396;
wire n_13823;
wire n_6128;
wire n_7037;
wire n_11820;
wire n_14900;
wire n_11587;
wire n_15350;
wire n_14863;
wire n_12081;
wire n_17046;
wire n_13157;
wire n_10314;
wire n_14966;
wire n_15982;
wire n_17449;
wire n_15646;
wire n_5749;
wire n_12296;
wire n_11697;
wire n_18329;
wire n_8427;
wire n_9339;
wire n_5332;
wire n_16554;
wire n_13038;
wire n_9596;
wire n_16495;
wire n_5108;
wire n_7409;
wire n_10006;
wire n_18196;
wire n_10667;
wire n_7258;
wire n_7432;
wire n_9156;
wire n_11441;
wire n_11242;
wire n_11916;
wire n_15209;
wire n_14591;
wire n_15818;
wire n_16832;
wire n_11435;
wire n_12804;
wire n_13999;
wire n_11471;
wire n_17064;
wire n_6334;
wire n_16765;
wire n_10346;
wire n_17607;
wire n_13236;
wire n_8984;
wire n_6848;
wire n_14502;
wire n_10539;
wire n_8345;
wire n_15590;
wire n_10414;
wire n_6321;
wire n_7765;
wire n_17948;
wire n_9708;
wire n_9268;
wire n_8764;
wire n_17666;
wire n_6794;
wire n_10340;
wire n_13310;
wire n_16865;
wire n_18225;
wire n_10245;
wire n_14479;
wire n_17761;
wire n_11644;
wire n_7761;
wire n_17165;
wire n_7197;
wire n_17477;
wire n_12466;
wire n_12701;
wire n_16585;
wire n_5489;
wire n_17886;
wire n_15560;
wire n_12106;
wire n_6400;
wire n_17192;
wire n_12560;
wire n_9097;
wire n_5057;
wire n_10280;
wire n_15909;
wire n_12895;
wire n_17498;
wire n_16066;
wire n_11432;
wire n_12342;
wire n_6705;
wire n_7775;
wire n_9636;
wire n_10256;
wire n_14559;
wire n_14676;
wire n_7619;
wire n_12125;
wire n_5436;
wire n_5907;
wire n_11120;
wire n_5072;
wire n_11391;
wire n_11164;
wire n_6044;
wire n_17113;
wire n_11527;
wire n_17374;
wire n_17667;
wire n_18277;
wire n_5286;
wire n_8083;
wire n_8853;
wire n_18292;
wire n_16736;
wire n_11371;
wire n_6495;
wire n_10917;
wire n_7403;
wire n_13933;
wire n_6902;
wire n_6470;
wire n_14619;
wire n_9473;
wire n_10727;
wire n_11591;
wire n_10145;
wire n_12341;
wire n_9560;
wire n_8038;
wire n_5569;
wire n_10938;
wire n_15631;
wire n_15525;
wire n_9175;
wire n_8711;
wire n_10976;
wire n_5439;
wire n_8229;
wire n_8949;
wire n_14248;
wire n_17776;
wire n_14928;
wire n_10612;
wire n_5619;
wire n_15127;
wire n_6481;
wire n_9810;
wire n_14079;
wire n_7548;
wire n_9244;
wire n_14878;
wire n_15444;
wire n_9584;
wire n_12047;
wire n_6534;
wire n_11460;
wire n_15112;
wire n_13289;
wire n_8567;
wire n_10797;
wire n_13320;
wire n_9439;
wire n_11915;
wire n_17056;
wire n_14224;
wire n_13210;
wire n_14015;
wire n_8655;
wire n_9235;
wire n_6181;
wire n_8705;
wire n_6728;
wire n_11642;
wire n_15313;
wire n_9043;
wire n_17430;
wire n_9768;
wire n_11306;
wire n_17176;
wire n_14566;
wire n_16796;
wire n_13549;
wire n_5119;
wire n_9037;
wire n_15334;
wire n_5715;
wire n_9085;
wire n_12434;
wire n_8085;
wire n_14874;
wire n_8777;
wire n_6133;
wire n_11891;
wire n_14951;
wire n_8852;
wire n_9264;
wire n_6528;
wire n_10114;
wire n_16546;
wire n_7604;
wire n_7407;
wire n_17050;
wire n_17790;
wire n_14499;
wire n_8185;
wire n_12998;
wire n_13427;
wire n_10845;
wire n_15942;
wire n_8513;
wire n_6670;
wire n_12248;
wire n_14155;
wire n_16226;
wire n_6774;
wire n_8365;
wire n_11007;
wire n_16909;
wire n_14229;
wire n_17047;
wire n_5887;
wire n_6741;
wire n_17562;
wire n_7424;
wire n_11557;
wire n_12405;
wire n_6038;
wire n_15320;
wire n_18305;
wire n_7727;
wire n_10599;
wire n_11231;
wire n_9550;
wire n_9836;
wire n_13228;
wire n_6282;
wire n_13244;
wire n_9929;
wire n_18217;
wire n_12134;
wire n_15877;
wire n_8035;
wire n_8505;
wire n_16317;
wire n_11399;
wire n_11092;
wire n_11163;
wire n_8874;
wire n_11542;
wire n_10008;
wire n_16195;
wire n_16446;
wire n_6700;
wire n_15362;
wire n_15742;
wire n_7334;
wire n_7684;
wire n_7755;
wire n_8098;
wire n_10623;
wire n_9187;
wire n_13880;
wire n_11276;
wire n_12770;
wire n_10511;
wire n_14418;
wire n_5932;
wire n_13011;
wire n_15629;
wire n_6178;
wire n_11575;
wire n_10503;
wire n_6234;
wire n_15226;
wire n_15180;
wire n_14880;
wire n_11732;
wire n_6012;
wire n_14518;
wire n_16630;
wire n_9406;
wire n_10857;
wire n_9342;
wire n_14119;
wire n_13222;
wire n_13323;
wire n_13604;
wire n_14321;
wire n_15146;
wire n_15279;
wire n_18087;
wire n_17678;
wire n_7787;
wire n_14808;
wire n_15750;
wire n_8067;
wire n_12421;
wire n_5092;
wire n_10708;
wire n_14136;
wire n_13106;
wire n_14950;
wire n_16946;
wire n_18139;
wire n_15961;
wire n_17349;
wire n_7849;
wire n_12550;
wire n_5186;
wire n_13126;
wire n_17520;
wire n_15772;
wire n_11045;
wire n_18239;
wire n_7367;
wire n_8619;
wire n_9851;
wire n_9559;
wire n_11993;
wire n_14818;
wire n_18114;
wire n_15448;
wire n_11508;
wire n_12755;
wire n_8679;
wire n_9806;
wire n_8644;
wire n_12306;
wire n_12965;
wire n_11982;
wire n_10516;
wire n_6715;
wire n_11395;
wire n_5828;
wire n_11634;
wire n_7200;
wire n_13068;
wire n_9860;
wire n_16668;
wire n_11887;
wire n_11301;
wire n_15031;
wire n_7582;
wire n_13402;
wire n_6337;
wire n_13997;
wire n_8923;
wire n_8970;
wire n_10119;
wire n_8332;
wire n_14302;
wire n_16938;
wire n_17547;
wire n_10548;
wire n_11010;
wire n_11408;
wire n_15182;
wire n_17223;
wire n_8632;
wire n_14829;
wire n_6770;
wire n_7745;
wire n_6743;
wire n_8876;
wire n_11670;
wire n_10733;
wire n_10547;
wire n_13218;
wire n_14011;
wire n_5238;
wire n_10067;
wire n_14646;
wire n_13958;
wire n_13239;
wire n_8856;
wire n_12603;
wire n_14230;
wire n_11604;
wire n_15907;
wire n_9240;
wire n_16575;
wire n_16926;
wire n_7877;
wire n_11506;
wire n_11666;
wire n_8945;
wire n_18115;
wire n_11503;
wire n_8918;
wire n_14433;
wire n_16140;
wire n_7799;
wire n_16022;
wire n_6682;
wire n_5054;
wire n_7673;
wire n_11857;
wire n_15886;
wire n_5631;
wire n_8028;
wire n_6539;
wire n_17844;
wire n_16925;
wire n_17239;
wire n_16035;
wire n_7243;
wire n_18294;
wire n_7179;
wire n_9345;
wire n_5399;
wire n_6314;
wire n_6617;
wire n_10222;
wire n_11193;
wire n_17084;
wire n_13983;
wire n_11293;
wire n_12439;
wire n_5694;
wire n_8774;
wire n_7274;
wire n_5326;
wire n_17808;
wire n_12072;
wire n_14199;
wire n_15920;
wire n_8779;
wire n_13949;
wire n_8968;
wire n_13941;
wire n_17021;
wire n_7608;
wire n_8404;
wire n_13090;
wire n_6595;
wire n_12558;
wire n_12244;
wire n_12199;
wire n_11214;
wire n_5459;
wire n_14986;
wire n_7738;
wire n_13851;
wire n_14209;
wire n_9223;
wire n_16971;
wire n_9499;
wire n_10647;
wire n_14177;
wire n_14495;
wire n_11362;
wire n_17597;
wire n_11288;
wire n_16788;
wire n_11409;
wire n_15091;
wire n_5528;
wire n_18186;
wire n_13036;
wire n_11027;
wire n_12996;
wire n_16283;
wire n_5391;
wire n_12873;
wire n_8073;
wire n_7785;
wire n_5422;
wire n_13225;
wire n_16129;
wire n_16448;
wire n_6385;
wire n_14485;
wire n_6289;
wire n_12591;
wire n_16518;
wire n_5267;
wire n_10581;
wire n_13587;
wire n_5523;
wire n_16205;
wire n_7373;
wire n_9576;
wire n_9120;
wire n_14832;
wire n_17415;
wire n_14917;
wire n_10097;
wire n_10405;
wire n_15009;
wire n_6186;
wire n_16356;
wire n_5153;
wire n_12726;
wire n_9651;
wire n_12833;
wire n_14206;
wire n_6257;
wire n_14240;
wire n_12690;
wire n_11031;
wire n_16574;
wire n_14080;
wire n_13076;
wire n_15787;
wire n_9386;
wire n_17592;
wire n_11285;
wire n_10813;
wire n_6852;
wire n_6346;
wire n_11346;
wire n_12618;
wire n_16087;
wire n_9779;
wire n_16475;
wire n_5044;
wire n_5809;
wire n_12414;
wire n_11513;
wire n_17802;
wire n_16142;
wire n_5365;
wire n_14888;
wire n_16743;
wire n_17116;
wire n_7587;
wire n_13729;
wire n_5045;
wire n_17175;
wire n_11250;
wire n_7874;
wire n_15992;
wire n_11340;
wire n_5354;
wire n_16882;
wire n_6274;
wire n_14381;
wire n_14739;
wire n_7372;
wire n_7760;
wire n_10588;
wire n_15699;
wire n_17609;
wire n_9635;
wire n_6818;
wire n_5915;
wire n_9444;
wire n_11190;
wire n_10943;
wire n_7226;
wire n_5452;
wire n_8930;
wire n_13992;
wire n_7057;
wire n_12736;
wire n_7685;
wire n_8031;
wire n_11818;
wire n_8750;
wire n_14193;
wire n_15840;
wire n_14649;
wire n_5595;
wire n_18015;
wire n_6609;
wire n_6815;
wire n_6753;
wire n_9364;
wire n_16334;
wire n_9512;
wire n_9581;
wire n_17274;
wire n_9317;
wire n_14625;
wire n_14661;
wire n_14968;
wire n_16811;
wire n_8593;
wire n_14047;
wire n_18258;
wire n_17548;
wire n_17529;
wire n_13592;
wire n_7730;
wire n_14262;
wire n_16970;
wire n_14723;
wire n_13165;
wire n_8509;
wire n_9314;
wire n_9459;
wire n_16773;
wire n_8405;
wire n_13659;
wire n_14558;
wire n_9549;
wire n_17299;
wire n_11564;
wire n_10641;
wire n_7913;
wire n_11719;
wire n_8492;
wire n_6764;
wire n_14569;
wire n_5535;
wire n_15795;
wire n_9275;
wire n_17453;
wire n_13670;
wire n_15245;
wire n_15598;
wire n_15102;
wire n_10210;
wire n_5370;
wire n_11944;
wire n_13967;
wire n_7706;
wire n_7891;
wire n_6391;
wire n_13248;
wire n_16093;
wire n_11785;
wire n_8088;
wire n_5372;
wire n_5299;
wire n_5594;
wire n_17359;
wire n_11754;
wire n_14369;
wire n_17991;
wire n_17040;
wire n_17066;
wire n_14301;
wire n_9865;
wire n_18191;
wire n_6471;
wire n_16816;
wire n_11075;
wire n_15960;
wire n_11511;
wire n_17370;
wire n_12981;
wire n_13061;
wire n_13546;
wire n_6627;
wire n_10027;
wire n_5761;
wire n_10263;
wire n_10722;
wire n_14422;
wire n_13005;
wire n_13978;
wire n_11771;
wire n_17940;
wire n_17224;
wire n_18177;
wire n_7203;
wire n_8429;
wire n_8854;
wire n_9757;
wire n_15121;
wire n_7512;
wire n_5550;
wire n_12333;
wire n_11912;
wire n_15405;
wire n_5082;
wire n_9656;
wire n_15442;
wire n_10426;
wire n_11284;
wire n_7215;
wire n_5209;
wire n_15033;
wire n_10246;
wire n_13500;
wire n_6636;
wire n_13004;
wire n_10617;
wire n_5929;
wire n_16146;
wire n_16662;
wire n_10909;
wire n_15347;
wire n_5559;
wire n_12694;
wire n_13972;
wire n_14295;
wire n_5478;
wire n_11298;
wire n_15733;
wire n_7388;
wire n_16225;
wire n_7694;
wire n_6243;
wire n_6488;
wire n_9629;
wire n_13864;
wire n_11185;
wire n_16532;
wire n_5102;
wire n_16590;
wire n_16347;
wire n_11498;
wire n_6022;
wire n_8686;
wire n_6457;
wire n_10299;
wire n_17312;
wire n_12904;
wire n_16900;
wire n_16571;
wire n_7982;
wire n_13874;
wire n_11384;
wire n_10763;
wire n_10494;
wire n_13520;
wire n_8773;
wire n_16772;
wire n_18296;
wire n_10743;
wire n_8225;
wire n_18047;
wire n_8583;
wire n_6867;
wire n_8887;
wire n_9556;
wire n_15494;
wire n_17646;
wire n_6538;
wire n_6230;
wire n_5868;
wire n_17517;
wire n_15524;
wire n_12810;
wire n_15989;
wire n_9259;
wire n_9995;
wire n_14680;
wire n_15946;
wire n_12820;
wire n_6633;
wire n_9371;
wire n_8080;
wire n_11496;
wire n_6187;
wire n_15662;
wire n_6172;
wire n_13274;
wire n_10050;
wire n_13827;
wire n_18273;
wire n_5275;
wire n_14927;
wire n_15196;
wire n_10702;
wire n_13572;
wire n_14236;
wire n_17864;
wire n_5071;
wire n_7311;
wire n_17315;
wire n_15606;
wire n_8964;
wire n_5989;
wire n_11768;
wire n_15051;
wire n_17385;
wire n_12085;
wire n_17173;
wire n_14748;
wire n_18080;
wire n_9008;
wire n_6574;
wire n_11388;
wire n_11683;
wire n_13786;
wire n_8929;
wire n_8539;
wire n_17075;
wire n_6395;
wire n_17932;
wire n_9484;
wire n_15660;
wire n_8745;
wire n_6854;
wire n_7996;
wire n_6233;
wire n_6456;
wire n_8776;
wire n_8588;
wire n_8554;
wire n_9319;
wire n_15568;
wire n_18313;
wire n_17282;
wire n_11748;
wire n_7488;
wire n_5227;
wire n_13463;
wire n_9442;
wire n_14351;
wire n_16564;
wire n_10165;
wire n_18095;
wire n_14385;
wire n_7198;
wire n_17240;
wire n_10366;
wire n_12207;
wire n_8802;
wire n_13242;
wire n_13194;
wire n_9587;
wire n_6784;
wire n_14915;
wire n_6168;
wire n_16076;
wire n_13871;
wire n_14168;
wire n_9904;
wire n_9157;
wire n_16781;
wire n_17754;
wire n_8431;
wire n_8453;
wire n_6766;
wire n_18197;
wire n_5242;
wire n_8955;
wire n_12510;
wire n_17608;
wire n_8634;
wire n_14575;
wire n_6330;
wire n_15978;
wire n_5520;
wire n_8896;
wire n_14695;
wire n_16706;
wire n_17310;
wire n_7950;
wire n_7249;
wire n_13741;
wire n_9713;
wire n_17462;
wire n_11210;
wire n_9452;
wire n_10104;
wire n_16111;
wire n_15539;
wire n_14186;
wire n_16771;
wire n_7336;
wire n_5947;
wire n_8837;
wire n_16439;
wire n_7031;
wire n_8907;
wire n_17082;
wire n_6799;
wire n_18073;
wire n_10115;
wire n_17085;
wire n_14514;
wire n_14853;
wire n_13654;
wire n_16400;
wire n_8015;
wire n_14149;
wire n_10397;
wire n_16417;
wire n_14454;
wire n_9974;
wire n_13245;
wire n_15221;
wire n_10398;
wire n_5920;
wire n_17030;
wire n_17480;
wire n_6672;
wire n_17851;
wire n_17563;
wire n_13193;
wire n_6149;
wire n_8256;
wire n_13739;
wire n_14578;
wire n_10065;
wire n_11156;
wire n_12628;
wire n_10087;
wire n_14003;
wire n_7142;
wire n_11598;
wire n_13977;
wire n_15692;
wire n_5808;
wire n_6054;
wire n_17710;
wire n_17247;
wire n_7089;
wire n_11176;
wire n_17336;
wire n_12687;
wire n_7916;
wire n_12260;
wire n_6450;
wire n_5294;
wire n_5353;
wire n_12445;
wire n_13776;
wire n_16920;
wire n_16990;
wire n_17463;
wire n_17665;
wire n_8074;
wire n_12878;
wire n_14023;
wire n_10174;
wire n_12281;
wire n_10266;
wire n_12879;
wire n_16050;
wire n_10509;
wire n_12355;
wire n_16819;
wire n_5458;
wire n_7042;
wire n_5617;
wire n_8778;
wire n_8039;
wire n_10415;
wire n_5244;
wire n_17907;
wire n_6523;
wire n_16639;
wire n_13127;
wire n_5382;
wire n_14581;
wire n_8065;
wire n_6107;
wire n_16282;
wire n_9634;
wire n_12601;
wire n_12004;
wire n_11893;
wire n_17023;
wire n_11828;
wire n_6775;
wire n_5274;
wire n_10873;
wire n_8194;
wire n_12291;
wire n_14125;
wire n_11582;
wire n_8207;
wire n_13109;
wire n_17428;
wire n_10106;
wire n_12474;
wire n_13414;
wire n_9241;
wire n_6232;
wire n_13688;
wire n_6445;
wire n_10422;
wire n_17955;
wire n_10736;
wire n_7181;
wire n_6134;
wire n_5384;
wire n_9903;
wire n_15712;
wire n_8582;
wire n_10378;
wire n_17063;
wire n_6056;
wire n_8537;
wire n_6932;
wire n_17438;
wire n_13425;
wire n_7036;
wire n_16922;
wire n_17341;
wire n_9615;
wire n_17516;
wire n_8951;
wire n_7759;
wire n_9600;
wire n_17425;
wire n_11095;
wire n_7818;
wire n_11180;
wire n_9748;
wire n_9945;
wire n_5125;
wire n_12024;
wire n_9927;
wire n_17145;
wire n_15574;
wire n_5587;
wire n_6855;
wire n_14072;
wire n_11876;
wire n_5789;
wire n_8217;
wire n_10046;
wire n_15157;
wire n_17392;
wire n_13182;
wire n_18158;
wire n_16525;
wire n_16952;
wire n_14787;
wire n_16237;
wire n_18157;
wire n_13911;
wire n_16165;
wire n_6585;
wire n_5787;
wire n_6369;
wire n_5056;
wire n_17201;
wire n_10954;
wire n_10388;
wire n_14883;
wire n_8437;
wire n_5249;
wire n_8849;
wire n_7447;
wire n_10659;
wire n_13124;
wire n_13956;
wire n_14617;
wire n_7944;
wire n_5198;
wire n_11709;
wire n_5360;
wire n_10804;
wire n_7455;
wire n_5829;
wire n_5233;
wire n_9295;
wire n_5269;
wire n_13819;
wire n_11602;
wire n_11304;
wire n_18255;
wire n_6252;
wire n_12934;
wire n_6493;
wire n_5866;
wire n_14843;
wire n_8568;
wire n_10239;
wire n_12723;
wire n_7947;
wire n_12428;
wire n_12857;
wire n_10841;
wire n_13566;
wire n_14315;
wire n_9916;
wire n_18167;
wire n_8980;
wire n_13682;
wire n_5899;
wire n_11630;
wire n_13339;
wire n_16702;
wire n_7629;
wire n_13478;
wire n_8051;
wire n_17580;
wire n_7104;
wire n_8716;
wire n_11461;
wire n_9844;
wire n_15376;
wire n_7601;
wire n_11135;
wire n_15467;
wire n_12520;
wire n_14303;
wire n_11994;
wire n_15998;
wire n_17346;
wire n_12457;
wire n_12743;
wire n_6026;
wire n_15177;
wire n_5247;
wire n_8030;
wire n_7757;
wire n_9316;
wire n_9663;
wire n_13918;
wire n_15714;
wire n_17117;
wire n_10168;
wire n_13526;
wire n_18267;
wire n_5865;
wire n_13019;
wire n_14335;
wire n_10075;
wire n_15275;
wire n_17811;
wire n_17386;
wire n_5317;
wire n_6544;
wire n_14848;
wire n_14989;
wire n_10068;
wire n_11596;
wire n_10276;
wire n_15332;
wire n_12533;
wire n_8749;
wire n_11024;
wire n_16877;
wire n_7138;
wire n_7290;
wire n_14424;
wire n_8544;
wire n_13077;
wire n_15419;
wire n_13524;
wire n_8249;
wire n_12555;
wire n_9628;
wire n_14560;
wire n_6679;
wire n_8496;
wire n_9789;
wire n_14273;
wire n_13296;
wire n_18324;
wire n_13891;
wire n_14090;
wire n_5380;
wire n_5924;
wire n_12839;
wire n_7625;
wire n_5822;
wire n_10495;
wire n_9299;
wire n_12251;
wire n_6259;
wire n_7284;
wire n_11246;
wire n_14693;
wire n_16551;
wire n_17545;
wire n_11715;
wire n_12766;
wire n_12983;
wire n_16830;
wire n_6390;
wire n_16361;
wire n_16266;
wire n_17596;
wire n_12573;
wire n_12945;
wire n_11970;
wire n_15047;
wire n_17567;
wire n_14839;
wire n_5786;
wire n_13466;
wire n_5182;
wire n_11113;
wire n_12451;
wire n_7971;
wire n_15310;
wire n_12542;
wire n_18033;
wire n_12376;
wire n_9022;
wire n_10927;
wire n_17834;
wire n_6630;
wire n_15463;
wire n_13116;
wire n_12585;
wire n_10704;
wire n_5658;
wire n_16133;
wire n_16817;
wire n_11613;
wire n_5388;
wire n_18108;
wire n_13256;
wire n_13968;
wire n_13942;
wire n_9427;
wire n_17003;
wire n_13231;
wire n_8698;
wire n_6279;
wire n_8695;
wire n_9344;
wire n_14461;
wire n_12530;
wire n_13718;
wire n_8751;
wire n_15618;
wire n_15671;
wire n_15789;
wire n_15979;
wire n_10603;
wire n_12875;
wire n_15864;
wire n_11085;
wire n_17156;
wire n_6813;
wire n_9764;
wire n_17292;
wire n_15720;
wire n_17164;
wire n_12808;
wire n_5564;
wire n_11294;
wire n_13024;
wire n_8273;
wire n_14897;
wire n_17485;
wire n_11021;
wire n_15918;
wire n_14041;
wire n_14817;
wire n_16490;
wire n_15675;
wire n_9242;
wire n_9498;
wire n_8442;
wire n_14799;
wire n_7106;
wire n_8472;
wire n_9535;
wire n_6042;
wire n_7644;
wire n_12494;
wire n_10011;
wire n_6057;
wire n_7529;
wire n_8986;
wire n_12488;
wire n_11905;
wire n_6675;
wire n_13147;
wire n_18289;
wire n_12229;
wire n_13740;
wire n_6476;
wire n_16576;
wire n_8200;
wire n_14397;
wire n_10055;
wire n_7907;
wire n_13064;
wire n_10982;
wire n_8188;
wire n_11951;
wire n_12219;
wire n_8528;
wire n_11926;
wire n_13041;
wire n_14879;
wire n_6207;
wire n_17814;
wire n_17749;
wire n_5539;
wire n_10764;
wire n_16894;
wire n_16177;
wire n_14333;
wire n_6268;
wire n_17660;
wire n_6878;
wire n_6286;
wire n_9088;
wire n_15490;
wire n_12630;
wire n_6524;
wire n_10787;
wire n_17964;
wire n_18320;
wire n_12910;
wire n_5547;
wire n_6225;
wire n_8920;
wire n_8267;
wire n_12758;
wire n_13302;
wire n_10972;
wire n_7297;
wire n_6291;
wire n_5893;
wire n_16587;
wire n_17794;
wire n_12883;
wire n_17507;
wire n_17865;
wire n_16042;
wire n_9734;
wire n_9505;
wire n_9664;
wire n_12672;
wire n_7199;
wire n_14167;
wire n_17094;
wire n_5273;
wire n_10262;
wire n_10826;
wire n_8360;
wire n_13828;
wire n_17527;
wire n_17916;
wire n_18221;
wire n_8036;
wire n_9510;
wire n_5261;
wire n_16121;
wire n_11423;
wire n_6520;
wire n_14162;
wire n_7853;
wire n_7648;
wire n_9413;
wire n_17616;
wire n_9888;
wire n_14085;
wire n_17818;
wire n_8393;
wire n_16932;
wire n_11484;
wire n_18056;
wire n_8821;
wire n_11760;
wire n_18088;
wire n_9863;
wire n_12946;
wire n_13397;
wire n_10881;
wire n_8160;
wire n_9199;
wire n_11370;
wire n_5193;
wire n_17214;
wire n_10707;
wire n_9014;
wire n_10204;
wire n_9411;
wire n_12394;
wire n_12613;
wire n_12706;
wire n_11909;
wire n_13882;
wire n_17423;
wire n_9336;
wire n_9360;
wire n_10556;
wire n_9543;
wire n_15374;
wire n_17303;
wire n_6024;
wire n_7866;
wire n_17742;
wire n_18172;
wire n_13252;
wire n_14783;
wire n_18317;
wire n_13174;
wire n_7487;
wire n_15553;
wire n_10717;
wire n_16640;
wire n_6425;
wire n_13931;
wire n_5993;
wire n_16293;
wire n_17784;
wire n_13541;
wire n_12978;
wire n_14201;
wire n_12253;
wire n_14710;
wire n_7638;
wire n_8833;
wire n_14296;
wire n_17890;
wire n_5703;
wire n_15169;
wire n_8240;
wire n_12450;
wire n_14857;
wire n_17134;
wire n_7988;
wire n_13579;
wire n_9404;
wire n_14643;
wire n_8579;
wire n_16331;
wire n_6432;
wire n_5534;
wire n_14354;
wire n_9678;
wire n_16104;
wire n_12444;
wire n_8258;
wire n_9854;
wire n_7259;
wire n_11071;
wire n_11979;
wire n_15414;
wire n_13050;
wire n_8626;
wire n_13384;
wire n_12289;
wire n_6540;
wire n_6955;
wire n_9481;
wire n_5174;
wire n_10862;
wire n_12583;
wire n_15872;
wire n_16375;
wire n_5157;
wire n_13936;
wire n_17897;
wire n_9672;
wire n_14009;
wire n_17591;
wire n_9893;
wire n_7237;
wire n_8935;
wire n_11928;
wire n_17339;
wire n_5087;
wire n_12590;
wire n_12596;
wire n_6388;
wire n_17472;
wire n_10240;
wire n_5904;
wire n_9478;
wire n_13465;
wire n_11792;
wire n_9266;
wire n_9813;
wire n_12551;
wire n_14026;
wire n_6760;
wire n_13817;
wire n_17868;
wire n_8009;
wire n_11329;
wire n_17519;
wire n_15700;
wire n_15929;
wire n_5620;
wire n_5061;
wire n_5750;
wire n_7063;
wire n_5572;
wire n_10338;
wire n_10205;
wire n_12034;
wire n_14275;
wire n_11573;
wire n_11703;
wire n_9042;
wire n_11671;
wire n_8012;
wire n_11445;
wire n_14692;
wire n_7576;
wire n_9506;
wire n_8608;
wire n_13946;
wire n_15655;
wire n_8008;
wire n_17142;
wire n_12498;
wire n_10285;
wire n_14040;
wire n_6795;
wire n_14464;
wire n_5881;
wire n_8079;
wire n_6664;
wire n_15695;
wire n_16090;
wire n_12228;
wire n_5815;
wire n_12378;
wire n_11832;
wire n_6261;
wire n_15953;
wire n_5873;
wire n_17195;
wire n_13926;
wire n_9666;
wire n_10112;
wire n_15200;
wire n_14163;
wire n_6487;
wire n_9146;
wire n_18140;
wire n_7734;
wire n_6729;
wire n_18271;
wire n_17016;
wire n_15046;
wire n_10056;
wire n_17309;
wire n_9862;
wire n_17408;
wire n_5755;
wire n_10283;
wire n_9274;
wire n_15407;
wire n_15680;
wire n_8702;
wire n_5949;
wire n_16302;
wire n_10469;
wire n_15999;
wire n_13944;
wire n_5195;
wire n_7483;
wire n_17277;
wire n_15926;
wire n_6608;
wire n_17722;
wire n_15498;
wire n_14145;
wire n_7858;
wire n_9619;
wire n_12742;
wire n_15172;
wire n_7385;
wire n_11088;
wire n_12423;
wire n_10618;
wire n_13902;
wire n_8576;
wire n_18241;
wire n_9508;
wire n_10105;
wire n_7668;
wire n_13008;
wire n_8662;
wire n_17839;
wire n_16567;
wire n_15694;
wire n_16577;
wire n_6663;
wire n_13504;
wire n_7476;
wire n_5955;
wire n_15022;
wire n_7327;
wire n_18084;
wire n_5763;
wire n_6656;
wire n_8436;
wire n_11154;
wire n_17803;
wire n_13491;
wire n_9987;
wire n_8124;
wire n_8148;
wire n_14135;
wire n_12518;
wire n_15519;
wire n_8033;
wire n_6843;
wire n_12764;
wire n_7953;
wire n_8343;
wire n_16599;
wire n_5246;
wire n_5964;
wire n_16322;
wire n_11065;
wire n_13812;
wire n_12417;
wire n_8118;
wire n_14182;
wire n_13751;
wire n_15850;
wire n_12209;
wire n_15143;
wire n_12882;
wire n_16809;
wire n_7266;
wire n_5164;
wire n_11449;
wire n_17786;
wire n_6969;
wire n_11447;
wire n_16445;
wire n_18302;
wire n_8741;
wire n_12427;
wire n_17908;
wire n_13894;
wire n_14217;
wire n_16700;
wire n_5665;
wire n_6485;
wire n_5340;
wire n_14882;
wire n_5498;
wire n_7100;
wire n_15173;
wire n_15012;
wire n_14541;
wire n_5783;
wire n_11123;
wire n_8478;
wire n_5183;
wire n_11319;
wire n_11676;
wire n_6075;
wire n_7082;
wire n_9569;
wire n_15439;
wire n_17375;
wire n_18030;
wire n_6120;
wire n_16878;
wire n_6659;
wire n_17322;
wire n_13513;
wire n_6750;
wire n_15685;
wire n_15808;
wire n_11018;
wire n_5549;
wire n_9935;
wire n_14477;
wire n_18212;
wire n_9707;
wire n_13663;
wire n_16410;
wire n_14664;
wire n_8376;
wire n_9827;
wire n_7689;
wire n_13858;
wire n_15674;
wire n_7132;
wire n_11537;
wire n_8763;
wire n_13361;
wire n_5442;
wire n_13792;
wire n_5739;
wire n_7824;
wire n_8996;
wire n_12707;
wire n_15832;
wire n_15949;
wire n_16112;
wire n_13161;
wire n_9007;
wire n_9797;
wire n_13132;
wire n_17713;
wire n_6003;
wire n_16167;
wire n_5385;
wire n_8726;
wire n_13662;
wire n_8799;
wire n_7796;
wire n_10670;
wire n_9053;
wire n_6478;
wire n_6066;
wire n_15607;
wire n_15232;
wire n_9450;
wire n_13272;
wire n_15512;
wire n_12437;
wire n_7034;
wire n_6086;
wire n_18025;
wire n_17645;
wire n_9121;
wire n_16797;
wire n_6650;
wire n_6224;
wire n_10789;
wire n_14725;
wire n_10387;
wire n_8303;
wire n_8796;
wire n_12941;
wire n_10661;
wire n_13859;
wire n_11638;
wire n_14476;
wire n_10088;
wire n_12026;
wire n_10629;
wire n_15246;
wire n_14208;
wire n_13898;
wire n_7084;
wire n_16442;
wire n_5845;
wire n_9617;
wire n_9089;
wire n_8883;
wire n_7293;
wire n_10505;
wire n_16634;
wire n_8251;
wire n_10247;
wire n_9236;
wire n_5990;
wire n_6175;
wire n_10860;
wire n_15464;
wire n_15387;
wire n_6060;
wire n_7253;
wire n_6891;
wire n_17687;
wire n_5663;
wire n_12537;
wire n_14547;
wire n_9493;
wire n_8860;
wire n_14364;
wire n_8003;
wire n_6410;
wire n_16927;
wire n_12607;
wire n_16746;
wire n_5973;
wire n_17283;
wire n_15184;
wire n_17471;
wire n_12958;
wire n_12849;
wire n_17421;
wire n_16185;
wire n_16633;
wire n_14849;
wire n_15822;
wire n_5537;
wire n_5304;
wire n_17143;
wire n_8524;
wire n_13835;
wire n_13863;
wire n_6059;
wire n_15713;
wire n_16200;
wire n_5130;
wire n_16985;
wire n_12329;
wire n_13650;
wire n_17220;
wire n_8914;
wire n_10524;
wire n_7520;
wire n_12032;
wire n_12159;
wire n_5162;
wire n_8520;
wire n_9490;
wire n_16686;
wire n_6103;
wire n_6809;
wire n_10376;
wire n_12737;
wire n_16991;
wire n_17895;
wire n_15328;
wire n_11213;
wire n_10986;
wire n_12504;
wire n_12987;
wire n_14780;
wire n_6267;
wire n_8165;
wire n_15163;
wire n_11523;
wire n_9525;
wire n_9127;
wire n_9119;
wire n_12521;
wire n_5855;
wire n_11903;
wire n_9002;
wire n_16645;
wire n_10069;
wire n_10697;
wire n_15300;
wire n_11100;
wire n_17752;
wire n_13695;
wire n_12866;
wire n_14030;
wire n_8330;
wire n_12226;
wire n_8682;
wire n_5757;
wire n_6437;
wire n_17389;
wire n_7331;
wire n_6610;
wire n_7918;
wire n_12170;
wire n_11440;
wire n_10259;
wire n_8467;
wire n_13216;
wire n_8775;
wire n_8886;
wire n_10844;
wire n_16692;
wire n_15371;
wire n_16613;
wire n_12482;
wire n_11476;
wire n_8696;
wire n_16002;
wire n_14742;
wire n_15600;
wire n_6957;
wire n_14658;
wire n_17994;
wire n_7514;
wire n_5704;
wire n_11966;
wire n_10330;
wire n_15571;
wire n_7163;
wire n_7620;
wire n_11115;
wire n_16105;
wire n_16443;
wire n_9867;
wire n_17186;
wire n_5473;
wire n_15113;
wire n_17354;
wire n_11765;
wire n_5946;
wire n_10197;
wire n_16372;
wire n_6711;
wire n_14648;
wire n_15501;
wire n_8464;
wire n_12440;
wire n_15580;
wire n_13313;
wire n_16249;
wire n_16847;
wire n_7445;
wire n_10584;
wire n_17514;
wire n_6847;
wire n_9131;
wire n_9790;
wire n_5177;
wire n_10522;
wire n_15011;
wire n_11200;
wire n_16072;
wire n_16291;
wire n_10752;
wire n_16188;
wire n_15152;
wire n_11332;
wire n_15426;
wire n_7123;
wire n_6384;
wire n_10854;
wire n_16118;
wire n_15244;
wire n_15122;
wire n_11189;
wire n_12834;
wire n_10768;
wire n_14791;
wire n_8720;
wire n_14779;
wire n_7959;
wire n_16269;
wire n_17380;
wire n_16806;
wire n_10542;
wire n_9611;
wire n_15203;
wire n_15352;
wire n_7563;
wire n_15217;
wire n_6298;
wire n_11170;
wire n_11337;
wire n_13987;
wire n_17300;
wire n_9032;
wire n_14218;
wire n_14982;
wire n_9428;
wire n_9990;
wire n_18146;
wire n_16062;
wire n_7361;
wire n_12929;
wire n_11278;
wire n_16029;
wire n_5172;
wire n_8186;
wire n_18062;
wire n_9705;
wire n_8890;
wire n_13497;
wire n_7322;
wire n_16979;
wire n_8219;
wire n_5710;
wire n_7453;
wire n_6067;
wire n_9774;
wire n_5070;
wire n_14941;
wire n_17326;
wire n_16986;
wire n_18321;
wire n_12022;
wire n_15725;
wire n_6377;
wire n_12358;
wire n_13793;
wire n_12242;
wire n_17775;
wire n_14010;
wire n_5566;
wire n_10419;
wire n_5414;
wire n_8738;
wire n_16084;
wire n_13186;
wire n_10645;
wire n_11713;
wire n_15691;
wire n_17487;
wire n_18107;
wire n_12214;
wire n_13282;
wire n_13988;
wire n_6348;
wire n_7713;
wire n_16427;
wire n_18210;
wire n_10412;
wire n_15545;
wire n_17748;
wire n_5296;
wire n_6129;
wire n_5450;
wire n_15147;
wire n_17167;
wire n_11195;
wire n_17251;
wire n_6834;
wire n_10124;
wire n_17331;
wire n_11975;
wire n_5313;
wire n_12254;
wire n_13073;
wire n_13580;
wire n_18053;
wire n_14178;
wire n_14816;
wire n_12320;
wire n_9374;
wire n_16421;
wire n_16462;
wire n_16536;
wire n_16419;
wire n_14960;
wire n_10737;
wire n_9792;
wire n_6136;
wire n_7261;
wire n_6723;
wire n_5834;
wire n_14008;
wire n_8066;
wire n_5874;
wire n_14459;
wire n_16229;
wire n_7977;
wire n_14582;
wire n_14970;
wire n_10294;
wire n_14063;
wire n_10687;
wire n_16643;
wire n_12763;
wire n_11402;
wire n_14597;
wire n_14976;
wire n_18310;
wire n_8342;
wire n_13527;
wire n_7508;
wire n_9771;
wire n_17985;
wire n_10480;
wire n_15549;
wire n_9712;
wire n_7021;
wire n_13831;
wire n_12627;
wire n_5270;
wire n_11345;
wire n_5956;
wire n_7834;
wire n_14670;
wire n_16147;
wire n_14349;
wire n_5188;
wire n_9905;
wire n_8571;
wire n_9308;
wire n_9163;
wire n_7000;
wire n_6078;
wire n_10243;
wire n_17684;
wire n_17431;
wire n_15627;
wire n_10721;
wire n_10038;
wire n_15905;
wire n_7921;
wire n_18126;
wire n_17482;
wire n_17579;
wire n_8877;
wire n_16178;
wire n_8862;
wire n_16247;
wire n_10144;
wire n_16414;
wire n_8402;
wire n_10410;
wire n_16364;
wire n_7130;
wire n_10823;
wire n_15070;
wire n_10176;
wire n_11714;
wire n_17356;
wire n_5823;
wire n_13687;
wire n_16355;
wire n_5465;
wire n_16605;
wire n_9387;
wire n_7538;
wire n_11778;
wire n_12492;
wire n_13794;
wire n_7517;
wire n_14948;
wire n_17905;
wire n_5853;
wire n_16436;
wire n_15504;
wire n_17343;
wire n_14758;
wire n_10799;
wire n_17724;
wire n_15994;
wire n_17467;
wire n_10315;
wire n_7077;
wire n_11300;
wire n_12561;
wire n_14497;
wire n_17009;
wire n_13382;
wire n_17692;
wire n_17677;
wire n_11338;
wire n_12359;
wire n_15528;
wire n_6642;
wire n_11577;
wire n_15276;
wire n_5467;
wire n_5522;
wire n_17093;
wire n_7346;
wire n_10525;
wire n_11930;
wire n_5148;
wire n_13353;
wire n_15076;
wire n_17065;
wire n_7333;
wire n_11334;
wire n_16158;
wire n_7546;
wire n_16779;
wire n_17494;
wire n_9847;
wire n_12688;
wire n_5934;
wire n_6942;
wire n_8418;
wire n_10932;
wire n_10227;
wire n_18291;
wire n_11096;
wire n_17099;
wire n_17554;
wire n_9577;
wire n_10951;
wire n_18278;
wire n_9111;
wire n_8805;
wire n_10646;
wire n_6511;
wire n_15219;
wire n_12635;
wire n_6507;
wire n_12677;
wire n_14338;
wire n_9513;
wire n_12568;
wire n_11482;
wire n_14819;
wire n_9853;
wire n_11759;
wire n_17639;
wire n_10710;
wire n_15137;
wire n_17044;
wire n_7319;
wire n_7997;
wire n_12610;
wire n_6497;
wire n_12639;
wire n_6001;
wire n_6007;
wire n_9130;
wire n_10409;
wire n_9941;
wire n_9135;
wire n_14414;
wire n_6606;
wire n_10709;
wire n_10633;
wire n_5318;
wire n_11829;
wire n_5395;
wire n_14327;
wire n_13901;
wire n_15346;
wire n_7078;
wire n_15292;
wire n_7047;
wire n_8144;
wire n_17304;
wire n_5067;
wire n_7107;
wire n_10606;
wire n_16360;
wire n_13047;
wire n_14077;
wire n_16070;
wire n_13049;
wire n_11936;
wire n_18208;
wire n_17476;
wire n_16758;
wire n_17689;
wire n_10325;
wire n_7469;
wire n_15668;
wire n_13055;
wire n_17968;
wire n_14786;
wire n_8111;
wire n_11308;

CKINVDCx5p33_ASAP7_75t_R g5039 ( 
.A(n_136),
.Y(n_5039)
);

CKINVDCx5p33_ASAP7_75t_R g5040 ( 
.A(n_913),
.Y(n_5040)
);

BUFx2_ASAP7_75t_L g5041 ( 
.A(n_3017),
.Y(n_5041)
);

CKINVDCx5p33_ASAP7_75t_R g5042 ( 
.A(n_229),
.Y(n_5042)
);

BUFx2_ASAP7_75t_L g5043 ( 
.A(n_1205),
.Y(n_5043)
);

CKINVDCx5p33_ASAP7_75t_R g5044 ( 
.A(n_4983),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_997),
.Y(n_5045)
);

CKINVDCx5p33_ASAP7_75t_R g5046 ( 
.A(n_1540),
.Y(n_5046)
);

CKINVDCx5p33_ASAP7_75t_R g5047 ( 
.A(n_1080),
.Y(n_5047)
);

INVx1_ASAP7_75t_SL g5048 ( 
.A(n_4232),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_3526),
.Y(n_5049)
);

CKINVDCx5p33_ASAP7_75t_R g5050 ( 
.A(n_2767),
.Y(n_5050)
);

CKINVDCx5p33_ASAP7_75t_R g5051 ( 
.A(n_4838),
.Y(n_5051)
);

INVxp67_ASAP7_75t_SL g5052 ( 
.A(n_346),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_3044),
.Y(n_5053)
);

BUFx3_ASAP7_75t_L g5054 ( 
.A(n_1186),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_4888),
.Y(n_5055)
);

CKINVDCx5p33_ASAP7_75t_R g5056 ( 
.A(n_3999),
.Y(n_5056)
);

BUFx6f_ASAP7_75t_L g5057 ( 
.A(n_1978),
.Y(n_5057)
);

CKINVDCx5p33_ASAP7_75t_R g5058 ( 
.A(n_4609),
.Y(n_5058)
);

CKINVDCx5p33_ASAP7_75t_R g5059 ( 
.A(n_2076),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_1146),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_1977),
.Y(n_5061)
);

CKINVDCx5p33_ASAP7_75t_R g5062 ( 
.A(n_123),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_4128),
.Y(n_5063)
);

CKINVDCx5p33_ASAP7_75t_R g5064 ( 
.A(n_3685),
.Y(n_5064)
);

CKINVDCx5p33_ASAP7_75t_R g5065 ( 
.A(n_4348),
.Y(n_5065)
);

CKINVDCx5p33_ASAP7_75t_R g5066 ( 
.A(n_4294),
.Y(n_5066)
);

INVx1_ASAP7_75t_L g5067 ( 
.A(n_4568),
.Y(n_5067)
);

INVx2_ASAP7_75t_L g5068 ( 
.A(n_577),
.Y(n_5068)
);

CKINVDCx5p33_ASAP7_75t_R g5069 ( 
.A(n_3814),
.Y(n_5069)
);

CKINVDCx5p33_ASAP7_75t_R g5070 ( 
.A(n_4229),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_2361),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4115),
.Y(n_5072)
);

BUFx10_ASAP7_75t_L g5073 ( 
.A(n_2208),
.Y(n_5073)
);

CKINVDCx5p33_ASAP7_75t_R g5074 ( 
.A(n_4152),
.Y(n_5074)
);

INVx1_ASAP7_75t_L g5075 ( 
.A(n_3154),
.Y(n_5075)
);

CKINVDCx5p33_ASAP7_75t_R g5076 ( 
.A(n_4159),
.Y(n_5076)
);

CKINVDCx5p33_ASAP7_75t_R g5077 ( 
.A(n_4388),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_3882),
.Y(n_5078)
);

CKINVDCx5p33_ASAP7_75t_R g5079 ( 
.A(n_1672),
.Y(n_5079)
);

CKINVDCx14_ASAP7_75t_R g5080 ( 
.A(n_2835),
.Y(n_5080)
);

CKINVDCx5p33_ASAP7_75t_R g5081 ( 
.A(n_1172),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_97),
.Y(n_5082)
);

CKINVDCx5p33_ASAP7_75t_R g5083 ( 
.A(n_3597),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4221),
.Y(n_5084)
);

INVx1_ASAP7_75t_SL g5085 ( 
.A(n_1608),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4244),
.Y(n_5086)
);

BUFx2_ASAP7_75t_L g5087 ( 
.A(n_1678),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_1962),
.Y(n_5088)
);

BUFx3_ASAP7_75t_L g5089 ( 
.A(n_3370),
.Y(n_5089)
);

CKINVDCx5p33_ASAP7_75t_R g5090 ( 
.A(n_4276),
.Y(n_5090)
);

CKINVDCx5p33_ASAP7_75t_R g5091 ( 
.A(n_3411),
.Y(n_5091)
);

CKINVDCx5p33_ASAP7_75t_R g5092 ( 
.A(n_1635),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_2425),
.Y(n_5093)
);

CKINVDCx5p33_ASAP7_75t_R g5094 ( 
.A(n_396),
.Y(n_5094)
);

CKINVDCx5p33_ASAP7_75t_R g5095 ( 
.A(n_3324),
.Y(n_5095)
);

CKINVDCx5p33_ASAP7_75t_R g5096 ( 
.A(n_3700),
.Y(n_5096)
);

CKINVDCx5p33_ASAP7_75t_R g5097 ( 
.A(n_611),
.Y(n_5097)
);

INVx1_ASAP7_75t_L g5098 ( 
.A(n_3134),
.Y(n_5098)
);

HB1xp67_ASAP7_75t_L g5099 ( 
.A(n_3745),
.Y(n_5099)
);

CKINVDCx5p33_ASAP7_75t_R g5100 ( 
.A(n_604),
.Y(n_5100)
);

CKINVDCx5p33_ASAP7_75t_R g5101 ( 
.A(n_4378),
.Y(n_5101)
);

CKINVDCx5p33_ASAP7_75t_R g5102 ( 
.A(n_3151),
.Y(n_5102)
);

INVx1_ASAP7_75t_SL g5103 ( 
.A(n_2646),
.Y(n_5103)
);

CKINVDCx5p33_ASAP7_75t_R g5104 ( 
.A(n_4965),
.Y(n_5104)
);

BUFx3_ASAP7_75t_L g5105 ( 
.A(n_1008),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_1284),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_1418),
.Y(n_5107)
);

CKINVDCx5p33_ASAP7_75t_R g5108 ( 
.A(n_1524),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_2944),
.Y(n_5109)
);

CKINVDCx5p33_ASAP7_75t_R g5110 ( 
.A(n_2096),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_4522),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_4880),
.Y(n_5112)
);

CKINVDCx5p33_ASAP7_75t_R g5113 ( 
.A(n_4227),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_4048),
.Y(n_5114)
);

CKINVDCx5p33_ASAP7_75t_R g5115 ( 
.A(n_1679),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_3827),
.Y(n_5116)
);

CKINVDCx5p33_ASAP7_75t_R g5117 ( 
.A(n_2317),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_3229),
.Y(n_5118)
);

CKINVDCx5p33_ASAP7_75t_R g5119 ( 
.A(n_3373),
.Y(n_5119)
);

INVx2_ASAP7_75t_L g5120 ( 
.A(n_4122),
.Y(n_5120)
);

INVx1_ASAP7_75t_SL g5121 ( 
.A(n_4220),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_1214),
.Y(n_5122)
);

CKINVDCx5p33_ASAP7_75t_R g5123 ( 
.A(n_1630),
.Y(n_5123)
);

CKINVDCx5p33_ASAP7_75t_R g5124 ( 
.A(n_4123),
.Y(n_5124)
);

INVx1_ASAP7_75t_L g5125 ( 
.A(n_3912),
.Y(n_5125)
);

CKINVDCx5p33_ASAP7_75t_R g5126 ( 
.A(n_757),
.Y(n_5126)
);

CKINVDCx5p33_ASAP7_75t_R g5127 ( 
.A(n_3851),
.Y(n_5127)
);

CKINVDCx5p33_ASAP7_75t_R g5128 ( 
.A(n_565),
.Y(n_5128)
);

CKINVDCx5p33_ASAP7_75t_R g5129 ( 
.A(n_3640),
.Y(n_5129)
);

CKINVDCx5p33_ASAP7_75t_R g5130 ( 
.A(n_692),
.Y(n_5130)
);

CKINVDCx5p33_ASAP7_75t_R g5131 ( 
.A(n_100),
.Y(n_5131)
);

CKINVDCx5p33_ASAP7_75t_R g5132 ( 
.A(n_3498),
.Y(n_5132)
);

BUFx3_ASAP7_75t_L g5133 ( 
.A(n_5018),
.Y(n_5133)
);

BUFx2_ASAP7_75t_L g5134 ( 
.A(n_3439),
.Y(n_5134)
);

CKINVDCx5p33_ASAP7_75t_R g5135 ( 
.A(n_1076),
.Y(n_5135)
);

HB1xp67_ASAP7_75t_L g5136 ( 
.A(n_4476),
.Y(n_5136)
);

CKINVDCx5p33_ASAP7_75t_R g5137 ( 
.A(n_4131),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_4259),
.Y(n_5138)
);

CKINVDCx5p33_ASAP7_75t_R g5139 ( 
.A(n_1575),
.Y(n_5139)
);

CKINVDCx20_ASAP7_75t_R g5140 ( 
.A(n_3733),
.Y(n_5140)
);

CKINVDCx5p33_ASAP7_75t_R g5141 ( 
.A(n_210),
.Y(n_5141)
);

CKINVDCx5p33_ASAP7_75t_R g5142 ( 
.A(n_2131),
.Y(n_5142)
);

CKINVDCx5p33_ASAP7_75t_R g5143 ( 
.A(n_3677),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_3862),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_4234),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_4655),
.Y(n_5146)
);

INVx1_ASAP7_75t_L g5147 ( 
.A(n_4226),
.Y(n_5147)
);

INVx2_ASAP7_75t_SL g5148 ( 
.A(n_2355),
.Y(n_5148)
);

INVx1_ASAP7_75t_L g5149 ( 
.A(n_3475),
.Y(n_5149)
);

BUFx3_ASAP7_75t_L g5150 ( 
.A(n_4291),
.Y(n_5150)
);

CKINVDCx16_ASAP7_75t_R g5151 ( 
.A(n_2840),
.Y(n_5151)
);

CKINVDCx5p33_ASAP7_75t_R g5152 ( 
.A(n_4242),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_961),
.Y(n_5153)
);

CKINVDCx5p33_ASAP7_75t_R g5154 ( 
.A(n_3088),
.Y(n_5154)
);

CKINVDCx20_ASAP7_75t_R g5155 ( 
.A(n_3058),
.Y(n_5155)
);

CKINVDCx5p33_ASAP7_75t_R g5156 ( 
.A(n_4465),
.Y(n_5156)
);

CKINVDCx5p33_ASAP7_75t_R g5157 ( 
.A(n_759),
.Y(n_5157)
);

CKINVDCx5p33_ASAP7_75t_R g5158 ( 
.A(n_78),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_405),
.Y(n_5159)
);

CKINVDCx5p33_ASAP7_75t_R g5160 ( 
.A(n_1099),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_4485),
.Y(n_5161)
);

CKINVDCx20_ASAP7_75t_R g5162 ( 
.A(n_4153),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_1515),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_1095),
.Y(n_5164)
);

CKINVDCx5p33_ASAP7_75t_R g5165 ( 
.A(n_538),
.Y(n_5165)
);

CKINVDCx5p33_ASAP7_75t_R g5166 ( 
.A(n_2158),
.Y(n_5166)
);

CKINVDCx5p33_ASAP7_75t_R g5167 ( 
.A(n_4425),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_4191),
.Y(n_5168)
);

CKINVDCx5p33_ASAP7_75t_R g5169 ( 
.A(n_2214),
.Y(n_5169)
);

BUFx6f_ASAP7_75t_L g5170 ( 
.A(n_3351),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_3797),
.Y(n_5171)
);

INVx2_ASAP7_75t_SL g5172 ( 
.A(n_1167),
.Y(n_5172)
);

CKINVDCx5p33_ASAP7_75t_R g5173 ( 
.A(n_4156),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_712),
.Y(n_5174)
);

BUFx5_ASAP7_75t_L g5175 ( 
.A(n_2393),
.Y(n_5175)
);

INVx3_ASAP7_75t_L g5176 ( 
.A(n_1490),
.Y(n_5176)
);

BUFx6f_ASAP7_75t_L g5177 ( 
.A(n_1718),
.Y(n_5177)
);

BUFx2_ASAP7_75t_SL g5178 ( 
.A(n_1075),
.Y(n_5178)
);

CKINVDCx5p33_ASAP7_75t_R g5179 ( 
.A(n_4269),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_1531),
.Y(n_5180)
);

CKINVDCx5p33_ASAP7_75t_R g5181 ( 
.A(n_4145),
.Y(n_5181)
);

CKINVDCx5p33_ASAP7_75t_R g5182 ( 
.A(n_3724),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_3858),
.Y(n_5183)
);

CKINVDCx14_ASAP7_75t_R g5184 ( 
.A(n_172),
.Y(n_5184)
);

CKINVDCx20_ASAP7_75t_R g5185 ( 
.A(n_2067),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_4296),
.Y(n_5186)
);

CKINVDCx5p33_ASAP7_75t_R g5187 ( 
.A(n_4288),
.Y(n_5187)
);

CKINVDCx5p33_ASAP7_75t_R g5188 ( 
.A(n_2353),
.Y(n_5188)
);

CKINVDCx5p33_ASAP7_75t_R g5189 ( 
.A(n_4773),
.Y(n_5189)
);

CKINVDCx5p33_ASAP7_75t_R g5190 ( 
.A(n_442),
.Y(n_5190)
);

CKINVDCx5p33_ASAP7_75t_R g5191 ( 
.A(n_4061),
.Y(n_5191)
);

CKINVDCx20_ASAP7_75t_R g5192 ( 
.A(n_3307),
.Y(n_5192)
);

INVx2_ASAP7_75t_L g5193 ( 
.A(n_1870),
.Y(n_5193)
);

BUFx2_ASAP7_75t_L g5194 ( 
.A(n_3564),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_3741),
.Y(n_5195)
);

CKINVDCx5p33_ASAP7_75t_R g5196 ( 
.A(n_3425),
.Y(n_5196)
);

CKINVDCx5p33_ASAP7_75t_R g5197 ( 
.A(n_2338),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_2175),
.Y(n_5198)
);

CKINVDCx5p33_ASAP7_75t_R g5199 ( 
.A(n_726),
.Y(n_5199)
);

CKINVDCx5p33_ASAP7_75t_R g5200 ( 
.A(n_181),
.Y(n_5200)
);

CKINVDCx5p33_ASAP7_75t_R g5201 ( 
.A(n_4263),
.Y(n_5201)
);

BUFx2_ASAP7_75t_SL g5202 ( 
.A(n_4300),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_1474),
.Y(n_5203)
);

CKINVDCx5p33_ASAP7_75t_R g5204 ( 
.A(n_2169),
.Y(n_5204)
);

CKINVDCx5p33_ASAP7_75t_R g5205 ( 
.A(n_3348),
.Y(n_5205)
);

BUFx3_ASAP7_75t_L g5206 ( 
.A(n_319),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_3661),
.Y(n_5207)
);

INVx2_ASAP7_75t_L g5208 ( 
.A(n_1123),
.Y(n_5208)
);

INVx2_ASAP7_75t_L g5209 ( 
.A(n_1917),
.Y(n_5209)
);

BUFx10_ASAP7_75t_L g5210 ( 
.A(n_1290),
.Y(n_5210)
);

CKINVDCx5p33_ASAP7_75t_R g5211 ( 
.A(n_621),
.Y(n_5211)
);

CKINVDCx5p33_ASAP7_75t_R g5212 ( 
.A(n_2370),
.Y(n_5212)
);

CKINVDCx5p33_ASAP7_75t_R g5213 ( 
.A(n_2114),
.Y(n_5213)
);

HB1xp67_ASAP7_75t_L g5214 ( 
.A(n_1304),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_2894),
.Y(n_5215)
);

BUFx10_ASAP7_75t_L g5216 ( 
.A(n_4012),
.Y(n_5216)
);

CKINVDCx5p33_ASAP7_75t_R g5217 ( 
.A(n_296),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_490),
.Y(n_5218)
);

INVx1_ASAP7_75t_L g5219 ( 
.A(n_1601),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_3799),
.Y(n_5220)
);

BUFx6f_ASAP7_75t_L g5221 ( 
.A(n_4086),
.Y(n_5221)
);

CKINVDCx5p33_ASAP7_75t_R g5222 ( 
.A(n_3185),
.Y(n_5222)
);

CKINVDCx5p33_ASAP7_75t_R g5223 ( 
.A(n_1946),
.Y(n_5223)
);

BUFx6f_ASAP7_75t_L g5224 ( 
.A(n_3210),
.Y(n_5224)
);

INVx1_ASAP7_75t_L g5225 ( 
.A(n_3147),
.Y(n_5225)
);

CKINVDCx5p33_ASAP7_75t_R g5226 ( 
.A(n_1312),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_2262),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_2684),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_2846),
.Y(n_5229)
);

CKINVDCx5p33_ASAP7_75t_R g5230 ( 
.A(n_3345),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_979),
.Y(n_5231)
);

CKINVDCx5p33_ASAP7_75t_R g5232 ( 
.A(n_1975),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_4467),
.Y(n_5233)
);

CKINVDCx5p33_ASAP7_75t_R g5234 ( 
.A(n_1733),
.Y(n_5234)
);

CKINVDCx20_ASAP7_75t_R g5235 ( 
.A(n_3350),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_4142),
.Y(n_5236)
);

INVx1_ASAP7_75t_L g5237 ( 
.A(n_1411),
.Y(n_5237)
);

CKINVDCx5p33_ASAP7_75t_R g5238 ( 
.A(n_3881),
.Y(n_5238)
);

CKINVDCx5p33_ASAP7_75t_R g5239 ( 
.A(n_4250),
.Y(n_5239)
);

CKINVDCx5p33_ASAP7_75t_R g5240 ( 
.A(n_4531),
.Y(n_5240)
);

CKINVDCx5p33_ASAP7_75t_R g5241 ( 
.A(n_3758),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_4192),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_4800),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_4030),
.Y(n_5244)
);

CKINVDCx5p33_ASAP7_75t_R g5245 ( 
.A(n_3911),
.Y(n_5245)
);

CKINVDCx5p33_ASAP7_75t_R g5246 ( 
.A(n_4273),
.Y(n_5246)
);

CKINVDCx5p33_ASAP7_75t_R g5247 ( 
.A(n_1778),
.Y(n_5247)
);

CKINVDCx5p33_ASAP7_75t_R g5248 ( 
.A(n_2867),
.Y(n_5248)
);

CKINVDCx5p33_ASAP7_75t_R g5249 ( 
.A(n_85),
.Y(n_5249)
);

CKINVDCx5p33_ASAP7_75t_R g5250 ( 
.A(n_15),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_4798),
.Y(n_5251)
);

CKINVDCx14_ASAP7_75t_R g5252 ( 
.A(n_4300),
.Y(n_5252)
);

CKINVDCx5p33_ASAP7_75t_R g5253 ( 
.A(n_3957),
.Y(n_5253)
);

CKINVDCx5p33_ASAP7_75t_R g5254 ( 
.A(n_4081),
.Y(n_5254)
);

CKINVDCx5p33_ASAP7_75t_R g5255 ( 
.A(n_2845),
.Y(n_5255)
);

INVxp67_ASAP7_75t_L g5256 ( 
.A(n_4134),
.Y(n_5256)
);

CKINVDCx5p33_ASAP7_75t_R g5257 ( 
.A(n_364),
.Y(n_5257)
);

CKINVDCx20_ASAP7_75t_R g5258 ( 
.A(n_1136),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_3198),
.Y(n_5259)
);

INVx1_ASAP7_75t_SL g5260 ( 
.A(n_4551),
.Y(n_5260)
);

CKINVDCx5p33_ASAP7_75t_R g5261 ( 
.A(n_2463),
.Y(n_5261)
);

INVxp67_ASAP7_75t_SL g5262 ( 
.A(n_869),
.Y(n_5262)
);

CKINVDCx5p33_ASAP7_75t_R g5263 ( 
.A(n_4256),
.Y(n_5263)
);

CKINVDCx16_ASAP7_75t_R g5264 ( 
.A(n_1497),
.Y(n_5264)
);

CKINVDCx5p33_ASAP7_75t_R g5265 ( 
.A(n_3474),
.Y(n_5265)
);

CKINVDCx5p33_ASAP7_75t_R g5266 ( 
.A(n_2189),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_5021),
.Y(n_5267)
);

CKINVDCx5p33_ASAP7_75t_R g5268 ( 
.A(n_2455),
.Y(n_5268)
);

BUFx2_ASAP7_75t_L g5269 ( 
.A(n_1098),
.Y(n_5269)
);

CKINVDCx5p33_ASAP7_75t_R g5270 ( 
.A(n_4105),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_4562),
.Y(n_5271)
);

CKINVDCx20_ASAP7_75t_R g5272 ( 
.A(n_3694),
.Y(n_5272)
);

BUFx5_ASAP7_75t_L g5273 ( 
.A(n_4884),
.Y(n_5273)
);

CKINVDCx5p33_ASAP7_75t_R g5274 ( 
.A(n_2891),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_894),
.Y(n_5275)
);

CKINVDCx5p33_ASAP7_75t_R g5276 ( 
.A(n_433),
.Y(n_5276)
);

CKINVDCx5p33_ASAP7_75t_R g5277 ( 
.A(n_4276),
.Y(n_5277)
);

CKINVDCx5p33_ASAP7_75t_R g5278 ( 
.A(n_653),
.Y(n_5278)
);

CKINVDCx20_ASAP7_75t_R g5279 ( 
.A(n_3113),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_499),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_4113),
.Y(n_5281)
);

CKINVDCx5p33_ASAP7_75t_R g5282 ( 
.A(n_2961),
.Y(n_5282)
);

CKINVDCx5p33_ASAP7_75t_R g5283 ( 
.A(n_1707),
.Y(n_5283)
);

CKINVDCx5p33_ASAP7_75t_R g5284 ( 
.A(n_3168),
.Y(n_5284)
);

CKINVDCx5p33_ASAP7_75t_R g5285 ( 
.A(n_1086),
.Y(n_5285)
);

BUFx3_ASAP7_75t_L g5286 ( 
.A(n_1749),
.Y(n_5286)
);

BUFx2_ASAP7_75t_L g5287 ( 
.A(n_4134),
.Y(n_5287)
);

CKINVDCx5p33_ASAP7_75t_R g5288 ( 
.A(n_4201),
.Y(n_5288)
);

CKINVDCx20_ASAP7_75t_R g5289 ( 
.A(n_3953),
.Y(n_5289)
);

BUFx10_ASAP7_75t_L g5290 ( 
.A(n_3777),
.Y(n_5290)
);

CKINVDCx5p33_ASAP7_75t_R g5291 ( 
.A(n_1893),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_2273),
.Y(n_5292)
);

CKINVDCx5p33_ASAP7_75t_R g5293 ( 
.A(n_1131),
.Y(n_5293)
);

CKINVDCx5p33_ASAP7_75t_R g5294 ( 
.A(n_2190),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_1396),
.Y(n_5295)
);

CKINVDCx5p33_ASAP7_75t_R g5296 ( 
.A(n_263),
.Y(n_5296)
);

INVx1_ASAP7_75t_SL g5297 ( 
.A(n_2325),
.Y(n_5297)
);

CKINVDCx5p33_ASAP7_75t_R g5298 ( 
.A(n_1371),
.Y(n_5298)
);

INVx1_ASAP7_75t_L g5299 ( 
.A(n_1646),
.Y(n_5299)
);

CKINVDCx5p33_ASAP7_75t_R g5300 ( 
.A(n_1330),
.Y(n_5300)
);

CKINVDCx5p33_ASAP7_75t_R g5301 ( 
.A(n_1731),
.Y(n_5301)
);

CKINVDCx16_ASAP7_75t_R g5302 ( 
.A(n_362),
.Y(n_5302)
);

CKINVDCx5p33_ASAP7_75t_R g5303 ( 
.A(n_1133),
.Y(n_5303)
);

CKINVDCx5p33_ASAP7_75t_R g5304 ( 
.A(n_1026),
.Y(n_5304)
);

CKINVDCx20_ASAP7_75t_R g5305 ( 
.A(n_1222),
.Y(n_5305)
);

INVx1_ASAP7_75t_L g5306 ( 
.A(n_385),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_3703),
.Y(n_5307)
);

INVx3_ASAP7_75t_L g5308 ( 
.A(n_4281),
.Y(n_5308)
);

CKINVDCx5p33_ASAP7_75t_R g5309 ( 
.A(n_1818),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_2806),
.Y(n_5310)
);

CKINVDCx5p33_ASAP7_75t_R g5311 ( 
.A(n_4197),
.Y(n_5311)
);

BUFx10_ASAP7_75t_L g5312 ( 
.A(n_4787),
.Y(n_5312)
);

INVx2_ASAP7_75t_L g5313 ( 
.A(n_3091),
.Y(n_5313)
);

CKINVDCx20_ASAP7_75t_R g5314 ( 
.A(n_3094),
.Y(n_5314)
);

CKINVDCx5p33_ASAP7_75t_R g5315 ( 
.A(n_4969),
.Y(n_5315)
);

CKINVDCx5p33_ASAP7_75t_R g5316 ( 
.A(n_1817),
.Y(n_5316)
);

CKINVDCx20_ASAP7_75t_R g5317 ( 
.A(n_1087),
.Y(n_5317)
);

CKINVDCx16_ASAP7_75t_R g5318 ( 
.A(n_3852),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_1407),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_3920),
.Y(n_5320)
);

CKINVDCx5p33_ASAP7_75t_R g5321 ( 
.A(n_4219),
.Y(n_5321)
);

CKINVDCx5p33_ASAP7_75t_R g5322 ( 
.A(n_3087),
.Y(n_5322)
);

INVx1_ASAP7_75t_SL g5323 ( 
.A(n_4422),
.Y(n_5323)
);

CKINVDCx5p33_ASAP7_75t_R g5324 ( 
.A(n_4181),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_4138),
.Y(n_5325)
);

CKINVDCx5p33_ASAP7_75t_R g5326 ( 
.A(n_1529),
.Y(n_5326)
);

BUFx3_ASAP7_75t_L g5327 ( 
.A(n_796),
.Y(n_5327)
);

BUFx3_ASAP7_75t_L g5328 ( 
.A(n_785),
.Y(n_5328)
);

CKINVDCx20_ASAP7_75t_R g5329 ( 
.A(n_1169),
.Y(n_5329)
);

BUFx2_ASAP7_75t_L g5330 ( 
.A(n_130),
.Y(n_5330)
);

CKINVDCx5p33_ASAP7_75t_R g5331 ( 
.A(n_2992),
.Y(n_5331)
);

INVx2_ASAP7_75t_L g5332 ( 
.A(n_4301),
.Y(n_5332)
);

BUFx8_ASAP7_75t_SL g5333 ( 
.A(n_1473),
.Y(n_5333)
);

CKINVDCx5p33_ASAP7_75t_R g5334 ( 
.A(n_4972),
.Y(n_5334)
);

CKINVDCx5p33_ASAP7_75t_R g5335 ( 
.A(n_1903),
.Y(n_5335)
);

CKINVDCx5p33_ASAP7_75t_R g5336 ( 
.A(n_2982),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_1563),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_4774),
.Y(n_5338)
);

INVx1_ASAP7_75t_SL g5339 ( 
.A(n_15),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_1144),
.Y(n_5340)
);

INVx1_ASAP7_75t_L g5341 ( 
.A(n_1373),
.Y(n_5341)
);

BUFx2_ASAP7_75t_L g5342 ( 
.A(n_201),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_4214),
.Y(n_5343)
);

CKINVDCx5p33_ASAP7_75t_R g5344 ( 
.A(n_3544),
.Y(n_5344)
);

CKINVDCx5p33_ASAP7_75t_R g5345 ( 
.A(n_3252),
.Y(n_5345)
);

CKINVDCx5p33_ASAP7_75t_R g5346 ( 
.A(n_1188),
.Y(n_5346)
);

CKINVDCx5p33_ASAP7_75t_R g5347 ( 
.A(n_1655),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_1416),
.Y(n_5348)
);

CKINVDCx5p33_ASAP7_75t_R g5349 ( 
.A(n_1933),
.Y(n_5349)
);

INVx2_ASAP7_75t_L g5350 ( 
.A(n_852),
.Y(n_5350)
);

CKINVDCx5p33_ASAP7_75t_R g5351 ( 
.A(n_351),
.Y(n_5351)
);

INVx1_ASAP7_75t_SL g5352 ( 
.A(n_1836),
.Y(n_5352)
);

CKINVDCx5p33_ASAP7_75t_R g5353 ( 
.A(n_2614),
.Y(n_5353)
);

CKINVDCx5p33_ASAP7_75t_R g5354 ( 
.A(n_12),
.Y(n_5354)
);

CKINVDCx5p33_ASAP7_75t_R g5355 ( 
.A(n_3433),
.Y(n_5355)
);

CKINVDCx16_ASAP7_75t_R g5356 ( 
.A(n_977),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_4271),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_4486),
.Y(n_5358)
);

CKINVDCx5p33_ASAP7_75t_R g5359 ( 
.A(n_4231),
.Y(n_5359)
);

CKINVDCx5p33_ASAP7_75t_R g5360 ( 
.A(n_309),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_4746),
.Y(n_5361)
);

INVx2_ASAP7_75t_L g5362 ( 
.A(n_4227),
.Y(n_5362)
);

BUFx10_ASAP7_75t_L g5363 ( 
.A(n_1233),
.Y(n_5363)
);

CKINVDCx5p33_ASAP7_75t_R g5364 ( 
.A(n_4756),
.Y(n_5364)
);

CKINVDCx5p33_ASAP7_75t_R g5365 ( 
.A(n_578),
.Y(n_5365)
);

CKINVDCx5p33_ASAP7_75t_R g5366 ( 
.A(n_2933),
.Y(n_5366)
);

INVx2_ASAP7_75t_L g5367 ( 
.A(n_3609),
.Y(n_5367)
);

CKINVDCx20_ASAP7_75t_R g5368 ( 
.A(n_510),
.Y(n_5368)
);

INVx1_ASAP7_75t_L g5369 ( 
.A(n_2380),
.Y(n_5369)
);

INVx1_ASAP7_75t_L g5370 ( 
.A(n_2211),
.Y(n_5370)
);

CKINVDCx5p33_ASAP7_75t_R g5371 ( 
.A(n_4149),
.Y(n_5371)
);

CKINVDCx5p33_ASAP7_75t_R g5372 ( 
.A(n_3799),
.Y(n_5372)
);

INVx2_ASAP7_75t_SL g5373 ( 
.A(n_1079),
.Y(n_5373)
);

BUFx3_ASAP7_75t_L g5374 ( 
.A(n_4360),
.Y(n_5374)
);

CKINVDCx5p33_ASAP7_75t_R g5375 ( 
.A(n_2973),
.Y(n_5375)
);

INVxp67_ASAP7_75t_L g5376 ( 
.A(n_4160),
.Y(n_5376)
);

CKINVDCx5p33_ASAP7_75t_R g5377 ( 
.A(n_2069),
.Y(n_5377)
);

CKINVDCx5p33_ASAP7_75t_R g5378 ( 
.A(n_2792),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_1276),
.Y(n_5379)
);

CKINVDCx5p33_ASAP7_75t_R g5380 ( 
.A(n_3376),
.Y(n_5380)
);

CKINVDCx5p33_ASAP7_75t_R g5381 ( 
.A(n_1071),
.Y(n_5381)
);

HB1xp67_ASAP7_75t_L g5382 ( 
.A(n_4021),
.Y(n_5382)
);

CKINVDCx5p33_ASAP7_75t_R g5383 ( 
.A(n_2909),
.Y(n_5383)
);

CKINVDCx20_ASAP7_75t_R g5384 ( 
.A(n_2801),
.Y(n_5384)
);

CKINVDCx5p33_ASAP7_75t_R g5385 ( 
.A(n_2608),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_593),
.Y(n_5386)
);

CKINVDCx20_ASAP7_75t_R g5387 ( 
.A(n_3339),
.Y(n_5387)
);

CKINVDCx20_ASAP7_75t_R g5388 ( 
.A(n_1844),
.Y(n_5388)
);

CKINVDCx5p33_ASAP7_75t_R g5389 ( 
.A(n_4287),
.Y(n_5389)
);

CKINVDCx5p33_ASAP7_75t_R g5390 ( 
.A(n_4199),
.Y(n_5390)
);

CKINVDCx5p33_ASAP7_75t_R g5391 ( 
.A(n_1058),
.Y(n_5391)
);

CKINVDCx5p33_ASAP7_75t_R g5392 ( 
.A(n_2439),
.Y(n_5392)
);

CKINVDCx5p33_ASAP7_75t_R g5393 ( 
.A(n_1454),
.Y(n_5393)
);

CKINVDCx5p33_ASAP7_75t_R g5394 ( 
.A(n_3712),
.Y(n_5394)
);

BUFx2_ASAP7_75t_SL g5395 ( 
.A(n_3474),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_4187),
.Y(n_5396)
);

INVx1_ASAP7_75t_L g5397 ( 
.A(n_4162),
.Y(n_5397)
);

INVx1_ASAP7_75t_SL g5398 ( 
.A(n_412),
.Y(n_5398)
);

CKINVDCx5p33_ASAP7_75t_R g5399 ( 
.A(n_3269),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_4474),
.Y(n_5400)
);

CKINVDCx5p33_ASAP7_75t_R g5401 ( 
.A(n_2464),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_8),
.Y(n_5402)
);

CKINVDCx5p33_ASAP7_75t_R g5403 ( 
.A(n_887),
.Y(n_5403)
);

CKINVDCx5p33_ASAP7_75t_R g5404 ( 
.A(n_4297),
.Y(n_5404)
);

BUFx10_ASAP7_75t_L g5405 ( 
.A(n_3611),
.Y(n_5405)
);

CKINVDCx5p33_ASAP7_75t_R g5406 ( 
.A(n_646),
.Y(n_5406)
);

CKINVDCx5p33_ASAP7_75t_R g5407 ( 
.A(n_195),
.Y(n_5407)
);

CKINVDCx5p33_ASAP7_75t_R g5408 ( 
.A(n_4151),
.Y(n_5408)
);

BUFx3_ASAP7_75t_L g5409 ( 
.A(n_1420),
.Y(n_5409)
);

CKINVDCx5p33_ASAP7_75t_R g5410 ( 
.A(n_189),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_648),
.Y(n_5411)
);

CKINVDCx5p33_ASAP7_75t_R g5412 ( 
.A(n_2902),
.Y(n_5412)
);

INVx2_ASAP7_75t_SL g5413 ( 
.A(n_4212),
.Y(n_5413)
);

INVx1_ASAP7_75t_L g5414 ( 
.A(n_1939),
.Y(n_5414)
);

CKINVDCx5p33_ASAP7_75t_R g5415 ( 
.A(n_2719),
.Y(n_5415)
);

INVx2_ASAP7_75t_L g5416 ( 
.A(n_4769),
.Y(n_5416)
);

CKINVDCx5p33_ASAP7_75t_R g5417 ( 
.A(n_2389),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_1591),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_2809),
.Y(n_5419)
);

CKINVDCx20_ASAP7_75t_R g5420 ( 
.A(n_212),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_2453),
.Y(n_5421)
);

CKINVDCx5p33_ASAP7_75t_R g5422 ( 
.A(n_4278),
.Y(n_5422)
);

CKINVDCx5p33_ASAP7_75t_R g5423 ( 
.A(n_4149),
.Y(n_5423)
);

CKINVDCx5p33_ASAP7_75t_R g5424 ( 
.A(n_2449),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_4163),
.Y(n_5425)
);

BUFx3_ASAP7_75t_L g5426 ( 
.A(n_3389),
.Y(n_5426)
);

INVx1_ASAP7_75t_L g5427 ( 
.A(n_4187),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_2874),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_3035),
.Y(n_5429)
);

CKINVDCx5p33_ASAP7_75t_R g5430 ( 
.A(n_4724),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_2757),
.Y(n_5431)
);

CKINVDCx5p33_ASAP7_75t_R g5432 ( 
.A(n_1783),
.Y(n_5432)
);

CKINVDCx5p33_ASAP7_75t_R g5433 ( 
.A(n_1924),
.Y(n_5433)
);

CKINVDCx16_ASAP7_75t_R g5434 ( 
.A(n_4215),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_2126),
.Y(n_5435)
);

CKINVDCx5p33_ASAP7_75t_R g5436 ( 
.A(n_2276),
.Y(n_5436)
);

INVx1_ASAP7_75t_L g5437 ( 
.A(n_986),
.Y(n_5437)
);

INVx1_ASAP7_75t_L g5438 ( 
.A(n_2470),
.Y(n_5438)
);

BUFx10_ASAP7_75t_L g5439 ( 
.A(n_2578),
.Y(n_5439)
);

INVx1_ASAP7_75t_SL g5440 ( 
.A(n_1578),
.Y(n_5440)
);

CKINVDCx5p33_ASAP7_75t_R g5441 ( 
.A(n_4167),
.Y(n_5441)
);

CKINVDCx5p33_ASAP7_75t_R g5442 ( 
.A(n_331),
.Y(n_5442)
);

CKINVDCx5p33_ASAP7_75t_R g5443 ( 
.A(n_1542),
.Y(n_5443)
);

CKINVDCx5p33_ASAP7_75t_R g5444 ( 
.A(n_4228),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_636),
.Y(n_5445)
);

CKINVDCx5p33_ASAP7_75t_R g5446 ( 
.A(n_2569),
.Y(n_5446)
);

INVx2_ASAP7_75t_L g5447 ( 
.A(n_247),
.Y(n_5447)
);

CKINVDCx5p33_ASAP7_75t_R g5448 ( 
.A(n_1118),
.Y(n_5448)
);

CKINVDCx5p33_ASAP7_75t_R g5449 ( 
.A(n_1532),
.Y(n_5449)
);

INVx1_ASAP7_75t_SL g5450 ( 
.A(n_2877),
.Y(n_5450)
);

CKINVDCx5p33_ASAP7_75t_R g5451 ( 
.A(n_3047),
.Y(n_5451)
);

CKINVDCx5p33_ASAP7_75t_R g5452 ( 
.A(n_1634),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_4049),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_3391),
.Y(n_5454)
);

CKINVDCx20_ASAP7_75t_R g5455 ( 
.A(n_732),
.Y(n_5455)
);

INVx1_ASAP7_75t_L g5456 ( 
.A(n_3185),
.Y(n_5456)
);

BUFx5_ASAP7_75t_L g5457 ( 
.A(n_2919),
.Y(n_5457)
);

CKINVDCx5p33_ASAP7_75t_R g5458 ( 
.A(n_4460),
.Y(n_5458)
);

CKINVDCx5p33_ASAP7_75t_R g5459 ( 
.A(n_2544),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_4190),
.Y(n_5460)
);

INVx2_ASAP7_75t_SL g5461 ( 
.A(n_3733),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_4173),
.Y(n_5462)
);

CKINVDCx5p33_ASAP7_75t_R g5463 ( 
.A(n_4669),
.Y(n_5463)
);

CKINVDCx5p33_ASAP7_75t_R g5464 ( 
.A(n_255),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_3116),
.Y(n_5465)
);

CKINVDCx5p33_ASAP7_75t_R g5466 ( 
.A(n_2431),
.Y(n_5466)
);

HB1xp67_ASAP7_75t_L g5467 ( 
.A(n_4302),
.Y(n_5467)
);

CKINVDCx20_ASAP7_75t_R g5468 ( 
.A(n_2248),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_214),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_509),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_4185),
.Y(n_5471)
);

CKINVDCx5p33_ASAP7_75t_R g5472 ( 
.A(n_4131),
.Y(n_5472)
);

INVx1_ASAP7_75t_L g5473 ( 
.A(n_4139),
.Y(n_5473)
);

CKINVDCx5p33_ASAP7_75t_R g5474 ( 
.A(n_4788),
.Y(n_5474)
);

CKINVDCx5p33_ASAP7_75t_R g5475 ( 
.A(n_4136),
.Y(n_5475)
);

BUFx2_ASAP7_75t_L g5476 ( 
.A(n_228),
.Y(n_5476)
);

CKINVDCx5p33_ASAP7_75t_R g5477 ( 
.A(n_4738),
.Y(n_5477)
);

CKINVDCx5p33_ASAP7_75t_R g5478 ( 
.A(n_3063),
.Y(n_5478)
);

INVx1_ASAP7_75t_SL g5479 ( 
.A(n_4176),
.Y(n_5479)
);

CKINVDCx5p33_ASAP7_75t_R g5480 ( 
.A(n_3727),
.Y(n_5480)
);

CKINVDCx5p33_ASAP7_75t_R g5481 ( 
.A(n_1783),
.Y(n_5481)
);

CKINVDCx5p33_ASAP7_75t_R g5482 ( 
.A(n_4241),
.Y(n_5482)
);

CKINVDCx20_ASAP7_75t_R g5483 ( 
.A(n_400),
.Y(n_5483)
);

CKINVDCx5p33_ASAP7_75t_R g5484 ( 
.A(n_1903),
.Y(n_5484)
);

CKINVDCx5p33_ASAP7_75t_R g5485 ( 
.A(n_771),
.Y(n_5485)
);

INVx2_ASAP7_75t_L g5486 ( 
.A(n_4290),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_3231),
.Y(n_5487)
);

CKINVDCx5p33_ASAP7_75t_R g5488 ( 
.A(n_4458),
.Y(n_5488)
);

CKINVDCx5p33_ASAP7_75t_R g5489 ( 
.A(n_2850),
.Y(n_5489)
);

CKINVDCx5p33_ASAP7_75t_R g5490 ( 
.A(n_3794),
.Y(n_5490)
);

CKINVDCx20_ASAP7_75t_R g5491 ( 
.A(n_1372),
.Y(n_5491)
);

CKINVDCx5p33_ASAP7_75t_R g5492 ( 
.A(n_457),
.Y(n_5492)
);

CKINVDCx5p33_ASAP7_75t_R g5493 ( 
.A(n_1140),
.Y(n_5493)
);

CKINVDCx5p33_ASAP7_75t_R g5494 ( 
.A(n_4278),
.Y(n_5494)
);

INVx2_ASAP7_75t_L g5495 ( 
.A(n_2102),
.Y(n_5495)
);

CKINVDCx5p33_ASAP7_75t_R g5496 ( 
.A(n_4126),
.Y(n_5496)
);

CKINVDCx5p33_ASAP7_75t_R g5497 ( 
.A(n_4239),
.Y(n_5497)
);

CKINVDCx5p33_ASAP7_75t_R g5498 ( 
.A(n_641),
.Y(n_5498)
);

CKINVDCx20_ASAP7_75t_R g5499 ( 
.A(n_4061),
.Y(n_5499)
);

CKINVDCx5p33_ASAP7_75t_R g5500 ( 
.A(n_106),
.Y(n_5500)
);

INVx1_ASAP7_75t_SL g5501 ( 
.A(n_1320),
.Y(n_5501)
);

CKINVDCx5p33_ASAP7_75t_R g5502 ( 
.A(n_4253),
.Y(n_5502)
);

CKINVDCx5p33_ASAP7_75t_R g5503 ( 
.A(n_4560),
.Y(n_5503)
);

INVx2_ASAP7_75t_L g5504 ( 
.A(n_1499),
.Y(n_5504)
);

CKINVDCx5p33_ASAP7_75t_R g5505 ( 
.A(n_4286),
.Y(n_5505)
);

CKINVDCx5p33_ASAP7_75t_R g5506 ( 
.A(n_4797),
.Y(n_5506)
);

INVx2_ASAP7_75t_L g5507 ( 
.A(n_358),
.Y(n_5507)
);

CKINVDCx5p33_ASAP7_75t_R g5508 ( 
.A(n_2038),
.Y(n_5508)
);

CKINVDCx5p33_ASAP7_75t_R g5509 ( 
.A(n_3010),
.Y(n_5509)
);

INVx1_ASAP7_75t_L g5510 ( 
.A(n_2726),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_4171),
.Y(n_5511)
);

CKINVDCx5p33_ASAP7_75t_R g5512 ( 
.A(n_3131),
.Y(n_5512)
);

CKINVDCx5p33_ASAP7_75t_R g5513 ( 
.A(n_2269),
.Y(n_5513)
);

CKINVDCx5p33_ASAP7_75t_R g5514 ( 
.A(n_2830),
.Y(n_5514)
);

BUFx10_ASAP7_75t_L g5515 ( 
.A(n_4100),
.Y(n_5515)
);

INVx1_ASAP7_75t_SL g5516 ( 
.A(n_3847),
.Y(n_5516)
);

CKINVDCx20_ASAP7_75t_R g5517 ( 
.A(n_651),
.Y(n_5517)
);

CKINVDCx5p33_ASAP7_75t_R g5518 ( 
.A(n_1163),
.Y(n_5518)
);

CKINVDCx20_ASAP7_75t_R g5519 ( 
.A(n_10),
.Y(n_5519)
);

INVx2_ASAP7_75t_L g5520 ( 
.A(n_3451),
.Y(n_5520)
);

INVx2_ASAP7_75t_SL g5521 ( 
.A(n_2547),
.Y(n_5521)
);

CKINVDCx5p33_ASAP7_75t_R g5522 ( 
.A(n_1229),
.Y(n_5522)
);

CKINVDCx16_ASAP7_75t_R g5523 ( 
.A(n_2906),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_1381),
.Y(n_5524)
);

INVx1_ASAP7_75t_L g5525 ( 
.A(n_2385),
.Y(n_5525)
);

INVx2_ASAP7_75t_L g5526 ( 
.A(n_570),
.Y(n_5526)
);

INVx1_ASAP7_75t_SL g5527 ( 
.A(n_4044),
.Y(n_5527)
);

CKINVDCx5p33_ASAP7_75t_R g5528 ( 
.A(n_3440),
.Y(n_5528)
);

INVx1_ASAP7_75t_SL g5529 ( 
.A(n_3752),
.Y(n_5529)
);

INVx1_ASAP7_75t_L g5530 ( 
.A(n_4164),
.Y(n_5530)
);

CKINVDCx5p33_ASAP7_75t_R g5531 ( 
.A(n_1132),
.Y(n_5531)
);

CKINVDCx5p33_ASAP7_75t_R g5532 ( 
.A(n_2587),
.Y(n_5532)
);

CKINVDCx20_ASAP7_75t_R g5533 ( 
.A(n_2360),
.Y(n_5533)
);

CKINVDCx5p33_ASAP7_75t_R g5534 ( 
.A(n_121),
.Y(n_5534)
);

CKINVDCx5p33_ASAP7_75t_R g5535 ( 
.A(n_2393),
.Y(n_5535)
);

BUFx3_ASAP7_75t_L g5536 ( 
.A(n_1553),
.Y(n_5536)
);

CKINVDCx5p33_ASAP7_75t_R g5537 ( 
.A(n_1018),
.Y(n_5537)
);

BUFx10_ASAP7_75t_L g5538 ( 
.A(n_2831),
.Y(n_5538)
);

INVxp67_ASAP7_75t_L g5539 ( 
.A(n_825),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_2519),
.Y(n_5540)
);

INVx2_ASAP7_75t_SL g5541 ( 
.A(n_1475),
.Y(n_5541)
);

INVx2_ASAP7_75t_L g5542 ( 
.A(n_4613),
.Y(n_5542)
);

CKINVDCx5p33_ASAP7_75t_R g5543 ( 
.A(n_3170),
.Y(n_5543)
);

CKINVDCx5p33_ASAP7_75t_R g5544 ( 
.A(n_2352),
.Y(n_5544)
);

CKINVDCx5p33_ASAP7_75t_R g5545 ( 
.A(n_2728),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_2917),
.Y(n_5546)
);

CKINVDCx5p33_ASAP7_75t_R g5547 ( 
.A(n_4819),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_1637),
.Y(n_5548)
);

INVx1_ASAP7_75t_L g5549 ( 
.A(n_4574),
.Y(n_5549)
);

CKINVDCx5p33_ASAP7_75t_R g5550 ( 
.A(n_3278),
.Y(n_5550)
);

CKINVDCx20_ASAP7_75t_R g5551 ( 
.A(n_1987),
.Y(n_5551)
);

INVx2_ASAP7_75t_SL g5552 ( 
.A(n_27),
.Y(n_5552)
);

CKINVDCx5p33_ASAP7_75t_R g5553 ( 
.A(n_9),
.Y(n_5553)
);

CKINVDCx5p33_ASAP7_75t_R g5554 ( 
.A(n_1221),
.Y(n_5554)
);

CKINVDCx5p33_ASAP7_75t_R g5555 ( 
.A(n_4900),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_2977),
.Y(n_5556)
);

CKINVDCx5p33_ASAP7_75t_R g5557 ( 
.A(n_4148),
.Y(n_5557)
);

CKINVDCx5p33_ASAP7_75t_R g5558 ( 
.A(n_1162),
.Y(n_5558)
);

CKINVDCx5p33_ASAP7_75t_R g5559 ( 
.A(n_1896),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_2681),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_2759),
.Y(n_5561)
);

CKINVDCx5p33_ASAP7_75t_R g5562 ( 
.A(n_2917),
.Y(n_5562)
);

CKINVDCx5p33_ASAP7_75t_R g5563 ( 
.A(n_218),
.Y(n_5563)
);

CKINVDCx5p33_ASAP7_75t_R g5564 ( 
.A(n_2671),
.Y(n_5564)
);

CKINVDCx5p33_ASAP7_75t_R g5565 ( 
.A(n_2687),
.Y(n_5565)
);

INVx1_ASAP7_75t_L g5566 ( 
.A(n_2438),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_3615),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_2286),
.Y(n_5568)
);

CKINVDCx5p33_ASAP7_75t_R g5569 ( 
.A(n_303),
.Y(n_5569)
);

CKINVDCx5p33_ASAP7_75t_R g5570 ( 
.A(n_2741),
.Y(n_5570)
);

CKINVDCx5p33_ASAP7_75t_R g5571 ( 
.A(n_723),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_951),
.Y(n_5572)
);

INVx1_ASAP7_75t_L g5573 ( 
.A(n_1274),
.Y(n_5573)
);

CKINVDCx20_ASAP7_75t_R g5574 ( 
.A(n_2646),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_3158),
.Y(n_5575)
);

CKINVDCx5p33_ASAP7_75t_R g5576 ( 
.A(n_4133),
.Y(n_5576)
);

HB1xp67_ASAP7_75t_L g5577 ( 
.A(n_4143),
.Y(n_5577)
);

CKINVDCx5p33_ASAP7_75t_R g5578 ( 
.A(n_2193),
.Y(n_5578)
);

CKINVDCx5p33_ASAP7_75t_R g5579 ( 
.A(n_1708),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_4979),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_3503),
.Y(n_5581)
);

CKINVDCx5p33_ASAP7_75t_R g5582 ( 
.A(n_4054),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_3260),
.Y(n_5583)
);

CKINVDCx5p33_ASAP7_75t_R g5584 ( 
.A(n_1276),
.Y(n_5584)
);

CKINVDCx5p33_ASAP7_75t_R g5585 ( 
.A(n_1043),
.Y(n_5585)
);

CKINVDCx5p33_ASAP7_75t_R g5586 ( 
.A(n_2147),
.Y(n_5586)
);

BUFx10_ASAP7_75t_L g5587 ( 
.A(n_4126),
.Y(n_5587)
);

INVx2_ASAP7_75t_SL g5588 ( 
.A(n_781),
.Y(n_5588)
);

CKINVDCx5p33_ASAP7_75t_R g5589 ( 
.A(n_1134),
.Y(n_5589)
);

CKINVDCx5p33_ASAP7_75t_R g5590 ( 
.A(n_4398),
.Y(n_5590)
);

CKINVDCx5p33_ASAP7_75t_R g5591 ( 
.A(n_4100),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_520),
.Y(n_5592)
);

CKINVDCx5p33_ASAP7_75t_R g5593 ( 
.A(n_371),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_2478),
.Y(n_5594)
);

BUFx10_ASAP7_75t_L g5595 ( 
.A(n_3599),
.Y(n_5595)
);

BUFx8_ASAP7_75t_SL g5596 ( 
.A(n_3521),
.Y(n_5596)
);

INVx1_ASAP7_75t_SL g5597 ( 
.A(n_3745),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_4998),
.Y(n_5598)
);

CKINVDCx5p33_ASAP7_75t_R g5599 ( 
.A(n_1374),
.Y(n_5599)
);

CKINVDCx5p33_ASAP7_75t_R g5600 ( 
.A(n_4261),
.Y(n_5600)
);

CKINVDCx5p33_ASAP7_75t_R g5601 ( 
.A(n_749),
.Y(n_5601)
);

CKINVDCx5p33_ASAP7_75t_R g5602 ( 
.A(n_4251),
.Y(n_5602)
);

CKINVDCx5p33_ASAP7_75t_R g5603 ( 
.A(n_512),
.Y(n_5603)
);

CKINVDCx5p33_ASAP7_75t_R g5604 ( 
.A(n_4595),
.Y(n_5604)
);

CKINVDCx5p33_ASAP7_75t_R g5605 ( 
.A(n_4516),
.Y(n_5605)
);

CKINVDCx5p33_ASAP7_75t_R g5606 ( 
.A(n_3360),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_4254),
.Y(n_5607)
);

CKINVDCx5p33_ASAP7_75t_R g5608 ( 
.A(n_85),
.Y(n_5608)
);

INVx1_ASAP7_75t_L g5609 ( 
.A(n_1516),
.Y(n_5609)
);

INVx1_ASAP7_75t_L g5610 ( 
.A(n_4022),
.Y(n_5610)
);

CKINVDCx5p33_ASAP7_75t_R g5611 ( 
.A(n_2819),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_872),
.Y(n_5612)
);

BUFx6f_ASAP7_75t_L g5613 ( 
.A(n_4948),
.Y(n_5613)
);

CKINVDCx5p33_ASAP7_75t_R g5614 ( 
.A(n_3704),
.Y(n_5614)
);

CKINVDCx5p33_ASAP7_75t_R g5615 ( 
.A(n_1149),
.Y(n_5615)
);

INVx1_ASAP7_75t_SL g5616 ( 
.A(n_28),
.Y(n_5616)
);

CKINVDCx20_ASAP7_75t_R g5617 ( 
.A(n_2477),
.Y(n_5617)
);

CKINVDCx5p33_ASAP7_75t_R g5618 ( 
.A(n_3117),
.Y(n_5618)
);

CKINVDCx5p33_ASAP7_75t_R g5619 ( 
.A(n_487),
.Y(n_5619)
);

CKINVDCx20_ASAP7_75t_R g5620 ( 
.A(n_3288),
.Y(n_5620)
);

BUFx3_ASAP7_75t_L g5621 ( 
.A(n_1965),
.Y(n_5621)
);

CKINVDCx5p33_ASAP7_75t_R g5622 ( 
.A(n_4897),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_1963),
.Y(n_5623)
);

CKINVDCx5p33_ASAP7_75t_R g5624 ( 
.A(n_3848),
.Y(n_5624)
);

CKINVDCx5p33_ASAP7_75t_R g5625 ( 
.A(n_737),
.Y(n_5625)
);

CKINVDCx5p33_ASAP7_75t_R g5626 ( 
.A(n_3988),
.Y(n_5626)
);

BUFx10_ASAP7_75t_L g5627 ( 
.A(n_3211),
.Y(n_5627)
);

CKINVDCx5p33_ASAP7_75t_R g5628 ( 
.A(n_923),
.Y(n_5628)
);

CKINVDCx5p33_ASAP7_75t_R g5629 ( 
.A(n_1852),
.Y(n_5629)
);

CKINVDCx5p33_ASAP7_75t_R g5630 ( 
.A(n_1626),
.Y(n_5630)
);

CKINVDCx5p33_ASAP7_75t_R g5631 ( 
.A(n_4117),
.Y(n_5631)
);

INVx1_ASAP7_75t_L g5632 ( 
.A(n_2777),
.Y(n_5632)
);

CKINVDCx5p33_ASAP7_75t_R g5633 ( 
.A(n_1036),
.Y(n_5633)
);

INVx1_ASAP7_75t_L g5634 ( 
.A(n_4274),
.Y(n_5634)
);

CKINVDCx5p33_ASAP7_75t_R g5635 ( 
.A(n_4193),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_3434),
.Y(n_5636)
);

CKINVDCx5p33_ASAP7_75t_R g5637 ( 
.A(n_246),
.Y(n_5637)
);

CKINVDCx5p33_ASAP7_75t_R g5638 ( 
.A(n_2390),
.Y(n_5638)
);

CKINVDCx20_ASAP7_75t_R g5639 ( 
.A(n_4195),
.Y(n_5639)
);

BUFx2_ASAP7_75t_L g5640 ( 
.A(n_1780),
.Y(n_5640)
);

INVx1_ASAP7_75t_L g5641 ( 
.A(n_4327),
.Y(n_5641)
);

CKINVDCx5p33_ASAP7_75t_R g5642 ( 
.A(n_2102),
.Y(n_5642)
);

CKINVDCx20_ASAP7_75t_R g5643 ( 
.A(n_1581),
.Y(n_5643)
);

CKINVDCx5p33_ASAP7_75t_R g5644 ( 
.A(n_2437),
.Y(n_5644)
);

INVx1_ASAP7_75t_L g5645 ( 
.A(n_1684),
.Y(n_5645)
);

CKINVDCx5p33_ASAP7_75t_R g5646 ( 
.A(n_2371),
.Y(n_5646)
);

INVx2_ASAP7_75t_L g5647 ( 
.A(n_2725),
.Y(n_5647)
);

INVx1_ASAP7_75t_L g5648 ( 
.A(n_705),
.Y(n_5648)
);

INVx1_ASAP7_75t_SL g5649 ( 
.A(n_1064),
.Y(n_5649)
);

INVx1_ASAP7_75t_L g5650 ( 
.A(n_3472),
.Y(n_5650)
);

INVx1_ASAP7_75t_L g5651 ( 
.A(n_4299),
.Y(n_5651)
);

CKINVDCx5p33_ASAP7_75t_R g5652 ( 
.A(n_3640),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_3069),
.Y(n_5653)
);

INVx2_ASAP7_75t_L g5654 ( 
.A(n_4166),
.Y(n_5654)
);

CKINVDCx5p33_ASAP7_75t_R g5655 ( 
.A(n_327),
.Y(n_5655)
);

CKINVDCx5p33_ASAP7_75t_R g5656 ( 
.A(n_5027),
.Y(n_5656)
);

CKINVDCx5p33_ASAP7_75t_R g5657 ( 
.A(n_1073),
.Y(n_5657)
);

CKINVDCx20_ASAP7_75t_R g5658 ( 
.A(n_1167),
.Y(n_5658)
);

CKINVDCx20_ASAP7_75t_R g5659 ( 
.A(n_518),
.Y(n_5659)
);

CKINVDCx5p33_ASAP7_75t_R g5660 ( 
.A(n_1811),
.Y(n_5660)
);

CKINVDCx20_ASAP7_75t_R g5661 ( 
.A(n_1383),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_2011),
.Y(n_5662)
);

CKINVDCx5p33_ASAP7_75t_R g5663 ( 
.A(n_230),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_2253),
.Y(n_5664)
);

CKINVDCx5p33_ASAP7_75t_R g5665 ( 
.A(n_4911),
.Y(n_5665)
);

CKINVDCx5p33_ASAP7_75t_R g5666 ( 
.A(n_1937),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_2014),
.Y(n_5667)
);

CKINVDCx5p33_ASAP7_75t_R g5668 ( 
.A(n_4648),
.Y(n_5668)
);

CKINVDCx5p33_ASAP7_75t_R g5669 ( 
.A(n_1075),
.Y(n_5669)
);

CKINVDCx5p33_ASAP7_75t_R g5670 ( 
.A(n_4132),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_897),
.Y(n_5671)
);

INVx2_ASAP7_75t_L g5672 ( 
.A(n_433),
.Y(n_5672)
);

INVx2_ASAP7_75t_L g5673 ( 
.A(n_340),
.Y(n_5673)
);

CKINVDCx5p33_ASAP7_75t_R g5674 ( 
.A(n_2030),
.Y(n_5674)
);

CKINVDCx5p33_ASAP7_75t_R g5675 ( 
.A(n_249),
.Y(n_5675)
);

BUFx6f_ASAP7_75t_L g5676 ( 
.A(n_3686),
.Y(n_5676)
);

CKINVDCx5p33_ASAP7_75t_R g5677 ( 
.A(n_362),
.Y(n_5677)
);

CKINVDCx5p33_ASAP7_75t_R g5678 ( 
.A(n_3885),
.Y(n_5678)
);

CKINVDCx5p33_ASAP7_75t_R g5679 ( 
.A(n_5030),
.Y(n_5679)
);

CKINVDCx5p33_ASAP7_75t_R g5680 ( 
.A(n_1658),
.Y(n_5680)
);

CKINVDCx5p33_ASAP7_75t_R g5681 ( 
.A(n_4429),
.Y(n_5681)
);

CKINVDCx5p33_ASAP7_75t_R g5682 ( 
.A(n_1027),
.Y(n_5682)
);

CKINVDCx5p33_ASAP7_75t_R g5683 ( 
.A(n_218),
.Y(n_5683)
);

CKINVDCx5p33_ASAP7_75t_R g5684 ( 
.A(n_3395),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_4157),
.Y(n_5685)
);

BUFx10_ASAP7_75t_L g5686 ( 
.A(n_2882),
.Y(n_5686)
);

CKINVDCx5p33_ASAP7_75t_R g5687 ( 
.A(n_3910),
.Y(n_5687)
);

CKINVDCx20_ASAP7_75t_R g5688 ( 
.A(n_4667),
.Y(n_5688)
);

CKINVDCx5p33_ASAP7_75t_R g5689 ( 
.A(n_2458),
.Y(n_5689)
);

BUFx6f_ASAP7_75t_L g5690 ( 
.A(n_3100),
.Y(n_5690)
);

INVx1_ASAP7_75t_L g5691 ( 
.A(n_3932),
.Y(n_5691)
);

CKINVDCx20_ASAP7_75t_R g5692 ( 
.A(n_2626),
.Y(n_5692)
);

CKINVDCx5p33_ASAP7_75t_R g5693 ( 
.A(n_4497),
.Y(n_5693)
);

CKINVDCx20_ASAP7_75t_R g5694 ( 
.A(n_2700),
.Y(n_5694)
);

INVx2_ASAP7_75t_L g5695 ( 
.A(n_1786),
.Y(n_5695)
);

CKINVDCx5p33_ASAP7_75t_R g5696 ( 
.A(n_4298),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_4289),
.Y(n_5697)
);

BUFx5_ASAP7_75t_L g5698 ( 
.A(n_3920),
.Y(n_5698)
);

CKINVDCx5p33_ASAP7_75t_R g5699 ( 
.A(n_4211),
.Y(n_5699)
);

CKINVDCx5p33_ASAP7_75t_R g5700 ( 
.A(n_1210),
.Y(n_5700)
);

CKINVDCx5p33_ASAP7_75t_R g5701 ( 
.A(n_4941),
.Y(n_5701)
);

CKINVDCx5p33_ASAP7_75t_R g5702 ( 
.A(n_2928),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_2499),
.Y(n_5703)
);

CKINVDCx5p33_ASAP7_75t_R g5704 ( 
.A(n_4223),
.Y(n_5704)
);

CKINVDCx5p33_ASAP7_75t_R g5705 ( 
.A(n_2778),
.Y(n_5705)
);

CKINVDCx5p33_ASAP7_75t_R g5706 ( 
.A(n_2472),
.Y(n_5706)
);

BUFx3_ASAP7_75t_L g5707 ( 
.A(n_4848),
.Y(n_5707)
);

CKINVDCx5p33_ASAP7_75t_R g5708 ( 
.A(n_4292),
.Y(n_5708)
);

INVxp67_ASAP7_75t_L g5709 ( 
.A(n_1740),
.Y(n_5709)
);

CKINVDCx5p33_ASAP7_75t_R g5710 ( 
.A(n_2206),
.Y(n_5710)
);

CKINVDCx5p33_ASAP7_75t_R g5711 ( 
.A(n_4755),
.Y(n_5711)
);

CKINVDCx5p33_ASAP7_75t_R g5712 ( 
.A(n_2746),
.Y(n_5712)
);

CKINVDCx5p33_ASAP7_75t_R g5713 ( 
.A(n_768),
.Y(n_5713)
);

CKINVDCx5p33_ASAP7_75t_R g5714 ( 
.A(n_4612),
.Y(n_5714)
);

CKINVDCx5p33_ASAP7_75t_R g5715 ( 
.A(n_3666),
.Y(n_5715)
);

INVx1_ASAP7_75t_L g5716 ( 
.A(n_494),
.Y(n_5716)
);

CKINVDCx5p33_ASAP7_75t_R g5717 ( 
.A(n_58),
.Y(n_5717)
);

CKINVDCx5p33_ASAP7_75t_R g5718 ( 
.A(n_1012),
.Y(n_5718)
);

CKINVDCx5p33_ASAP7_75t_R g5719 ( 
.A(n_4125),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_462),
.Y(n_5720)
);

CKINVDCx5p33_ASAP7_75t_R g5721 ( 
.A(n_1914),
.Y(n_5721)
);

INVx1_ASAP7_75t_L g5722 ( 
.A(n_2984),
.Y(n_5722)
);

CKINVDCx5p33_ASAP7_75t_R g5723 ( 
.A(n_3908),
.Y(n_5723)
);

CKINVDCx5p33_ASAP7_75t_R g5724 ( 
.A(n_368),
.Y(n_5724)
);

CKINVDCx5p33_ASAP7_75t_R g5725 ( 
.A(n_4140),
.Y(n_5725)
);

CKINVDCx5p33_ASAP7_75t_R g5726 ( 
.A(n_175),
.Y(n_5726)
);

CKINVDCx5p33_ASAP7_75t_R g5727 ( 
.A(n_498),
.Y(n_5727)
);

INVx2_ASAP7_75t_L g5728 ( 
.A(n_2674),
.Y(n_5728)
);

CKINVDCx5p33_ASAP7_75t_R g5729 ( 
.A(n_4257),
.Y(n_5729)
);

CKINVDCx5p33_ASAP7_75t_R g5730 ( 
.A(n_4272),
.Y(n_5730)
);

CKINVDCx20_ASAP7_75t_R g5731 ( 
.A(n_1569),
.Y(n_5731)
);

CKINVDCx20_ASAP7_75t_R g5732 ( 
.A(n_748),
.Y(n_5732)
);

CKINVDCx5p33_ASAP7_75t_R g5733 ( 
.A(n_643),
.Y(n_5733)
);

CKINVDCx5p33_ASAP7_75t_R g5734 ( 
.A(n_383),
.Y(n_5734)
);

CKINVDCx5p33_ASAP7_75t_R g5735 ( 
.A(n_4260),
.Y(n_5735)
);

CKINVDCx5p33_ASAP7_75t_R g5736 ( 
.A(n_1916),
.Y(n_5736)
);

CKINVDCx5p33_ASAP7_75t_R g5737 ( 
.A(n_3574),
.Y(n_5737)
);

CKINVDCx5p33_ASAP7_75t_R g5738 ( 
.A(n_4771),
.Y(n_5738)
);

CKINVDCx20_ASAP7_75t_R g5739 ( 
.A(n_3913),
.Y(n_5739)
);

CKINVDCx5p33_ASAP7_75t_R g5740 ( 
.A(n_3438),
.Y(n_5740)
);

CKINVDCx16_ASAP7_75t_R g5741 ( 
.A(n_1135),
.Y(n_5741)
);

HB1xp67_ASAP7_75t_L g5742 ( 
.A(n_2573),
.Y(n_5742)
);

CKINVDCx5p33_ASAP7_75t_R g5743 ( 
.A(n_4686),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_4642),
.Y(n_5744)
);

INVx2_ASAP7_75t_SL g5745 ( 
.A(n_4189),
.Y(n_5745)
);

CKINVDCx5p33_ASAP7_75t_R g5746 ( 
.A(n_3784),
.Y(n_5746)
);

CKINVDCx5p33_ASAP7_75t_R g5747 ( 
.A(n_451),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_4580),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_883),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_4406),
.Y(n_5750)
);

INVx1_ASAP7_75t_L g5751 ( 
.A(n_2285),
.Y(n_5751)
);

CKINVDCx5p33_ASAP7_75t_R g5752 ( 
.A(n_145),
.Y(n_5752)
);

CKINVDCx5p33_ASAP7_75t_R g5753 ( 
.A(n_3270),
.Y(n_5753)
);

INVx1_ASAP7_75t_SL g5754 ( 
.A(n_879),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_761),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_633),
.Y(n_5756)
);

CKINVDCx5p33_ASAP7_75t_R g5757 ( 
.A(n_2681),
.Y(n_5757)
);

CKINVDCx20_ASAP7_75t_R g5758 ( 
.A(n_3804),
.Y(n_5758)
);

INVx1_ASAP7_75t_L g5759 ( 
.A(n_4710),
.Y(n_5759)
);

INVxp33_ASAP7_75t_L g5760 ( 
.A(n_78),
.Y(n_5760)
);

CKINVDCx5p33_ASAP7_75t_R g5761 ( 
.A(n_125),
.Y(n_5761)
);

CKINVDCx14_ASAP7_75t_R g5762 ( 
.A(n_783),
.Y(n_5762)
);

CKINVDCx5p33_ASAP7_75t_R g5763 ( 
.A(n_2606),
.Y(n_5763)
);

CKINVDCx5p33_ASAP7_75t_R g5764 ( 
.A(n_4386),
.Y(n_5764)
);

INVx1_ASAP7_75t_SL g5765 ( 
.A(n_4535),
.Y(n_5765)
);

CKINVDCx5p33_ASAP7_75t_R g5766 ( 
.A(n_545),
.Y(n_5766)
);

CKINVDCx5p33_ASAP7_75t_R g5767 ( 
.A(n_1109),
.Y(n_5767)
);

CKINVDCx5p33_ASAP7_75t_R g5768 ( 
.A(n_4950),
.Y(n_5768)
);

CKINVDCx5p33_ASAP7_75t_R g5769 ( 
.A(n_3480),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_1078),
.Y(n_5770)
);

CKINVDCx20_ASAP7_75t_R g5771 ( 
.A(n_4466),
.Y(n_5771)
);

CKINVDCx5p33_ASAP7_75t_R g5772 ( 
.A(n_2279),
.Y(n_5772)
);

BUFx2_ASAP7_75t_L g5773 ( 
.A(n_840),
.Y(n_5773)
);

CKINVDCx5p33_ASAP7_75t_R g5774 ( 
.A(n_3928),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_4119),
.Y(n_5775)
);

CKINVDCx5p33_ASAP7_75t_R g5776 ( 
.A(n_3024),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_3171),
.Y(n_5777)
);

CKINVDCx5p33_ASAP7_75t_R g5778 ( 
.A(n_877),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_1387),
.Y(n_5779)
);

INVx1_ASAP7_75t_L g5780 ( 
.A(n_4224),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_2327),
.Y(n_5781)
);

CKINVDCx5p33_ASAP7_75t_R g5782 ( 
.A(n_1340),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_3573),
.Y(n_5783)
);

INVx2_ASAP7_75t_L g5784 ( 
.A(n_3892),
.Y(n_5784)
);

CKINVDCx5p33_ASAP7_75t_R g5785 ( 
.A(n_552),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_3682),
.Y(n_5786)
);

INVx2_ASAP7_75t_L g5787 ( 
.A(n_3036),
.Y(n_5787)
);

INVx1_ASAP7_75t_SL g5788 ( 
.A(n_4235),
.Y(n_5788)
);

CKINVDCx14_ASAP7_75t_R g5789 ( 
.A(n_2500),
.Y(n_5789)
);

CKINVDCx5p33_ASAP7_75t_R g5790 ( 
.A(n_639),
.Y(n_5790)
);

INVx1_ASAP7_75t_L g5791 ( 
.A(n_112),
.Y(n_5791)
);

INVx1_ASAP7_75t_SL g5792 ( 
.A(n_370),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_219),
.Y(n_5793)
);

CKINVDCx5p33_ASAP7_75t_R g5794 ( 
.A(n_3896),
.Y(n_5794)
);

CKINVDCx5p33_ASAP7_75t_R g5795 ( 
.A(n_312),
.Y(n_5795)
);

CKINVDCx5p33_ASAP7_75t_R g5796 ( 
.A(n_603),
.Y(n_5796)
);

INVx2_ASAP7_75t_SL g5797 ( 
.A(n_4611),
.Y(n_5797)
);

CKINVDCx5p33_ASAP7_75t_R g5798 ( 
.A(n_1874),
.Y(n_5798)
);

CKINVDCx5p33_ASAP7_75t_R g5799 ( 
.A(n_4242),
.Y(n_5799)
);

CKINVDCx5p33_ASAP7_75t_R g5800 ( 
.A(n_4118),
.Y(n_5800)
);

CKINVDCx5p33_ASAP7_75t_R g5801 ( 
.A(n_839),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_2718),
.Y(n_5802)
);

CKINVDCx5p33_ASAP7_75t_R g5803 ( 
.A(n_3545),
.Y(n_5803)
);

CKINVDCx5p33_ASAP7_75t_R g5804 ( 
.A(n_463),
.Y(n_5804)
);

INVx1_ASAP7_75t_L g5805 ( 
.A(n_4243),
.Y(n_5805)
);

INVx1_ASAP7_75t_L g5806 ( 
.A(n_2304),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_3916),
.Y(n_5807)
);

CKINVDCx5p33_ASAP7_75t_R g5808 ( 
.A(n_1969),
.Y(n_5808)
);

CKINVDCx5p33_ASAP7_75t_R g5809 ( 
.A(n_1886),
.Y(n_5809)
);

INVx1_ASAP7_75t_L g5810 ( 
.A(n_4636),
.Y(n_5810)
);

CKINVDCx5p33_ASAP7_75t_R g5811 ( 
.A(n_414),
.Y(n_5811)
);

INVx1_ASAP7_75t_SL g5812 ( 
.A(n_3723),
.Y(n_5812)
);

INVx1_ASAP7_75t_L g5813 ( 
.A(n_4155),
.Y(n_5813)
);

INVxp67_ASAP7_75t_L g5814 ( 
.A(n_4980),
.Y(n_5814)
);

CKINVDCx5p33_ASAP7_75t_R g5815 ( 
.A(n_720),
.Y(n_5815)
);

BUFx3_ASAP7_75t_L g5816 ( 
.A(n_4154),
.Y(n_5816)
);

CKINVDCx5p33_ASAP7_75t_R g5817 ( 
.A(n_1890),
.Y(n_5817)
);

CKINVDCx5p33_ASAP7_75t_R g5818 ( 
.A(n_1461),
.Y(n_5818)
);

CKINVDCx5p33_ASAP7_75t_R g5819 ( 
.A(n_3828),
.Y(n_5819)
);

BUFx2_ASAP7_75t_L g5820 ( 
.A(n_2633),
.Y(n_5820)
);

BUFx6f_ASAP7_75t_L g5821 ( 
.A(n_4144),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_4249),
.Y(n_5822)
);

INVx1_ASAP7_75t_L g5823 ( 
.A(n_2018),
.Y(n_5823)
);

INVx1_ASAP7_75t_L g5824 ( 
.A(n_1745),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_1807),
.Y(n_5825)
);

INVx2_ASAP7_75t_SL g5826 ( 
.A(n_148),
.Y(n_5826)
);

CKINVDCx5p33_ASAP7_75t_R g5827 ( 
.A(n_4238),
.Y(n_5827)
);

CKINVDCx5p33_ASAP7_75t_R g5828 ( 
.A(n_504),
.Y(n_5828)
);

BUFx3_ASAP7_75t_L g5829 ( 
.A(n_4127),
.Y(n_5829)
);

CKINVDCx14_ASAP7_75t_R g5830 ( 
.A(n_4161),
.Y(n_5830)
);

INVx1_ASAP7_75t_L g5831 ( 
.A(n_59),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_3220),
.Y(n_5832)
);

INVxp67_ASAP7_75t_L g5833 ( 
.A(n_916),
.Y(n_5833)
);

CKINVDCx20_ASAP7_75t_R g5834 ( 
.A(n_3567),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_2939),
.Y(n_5835)
);

CKINVDCx5p33_ASAP7_75t_R g5836 ( 
.A(n_2579),
.Y(n_5836)
);

CKINVDCx5p33_ASAP7_75t_R g5837 ( 
.A(n_4218),
.Y(n_5837)
);

CKINVDCx20_ASAP7_75t_R g5838 ( 
.A(n_3651),
.Y(n_5838)
);

CKINVDCx20_ASAP7_75t_R g5839 ( 
.A(n_3708),
.Y(n_5839)
);

CKINVDCx5p33_ASAP7_75t_R g5840 ( 
.A(n_2493),
.Y(n_5840)
);

CKINVDCx5p33_ASAP7_75t_R g5841 ( 
.A(n_611),
.Y(n_5841)
);

HB1xp67_ASAP7_75t_L g5842 ( 
.A(n_3855),
.Y(n_5842)
);

CKINVDCx5p33_ASAP7_75t_R g5843 ( 
.A(n_2050),
.Y(n_5843)
);

CKINVDCx5p33_ASAP7_75t_R g5844 ( 
.A(n_3674),
.Y(n_5844)
);

CKINVDCx5p33_ASAP7_75t_R g5845 ( 
.A(n_261),
.Y(n_5845)
);

INVx2_ASAP7_75t_L g5846 ( 
.A(n_624),
.Y(n_5846)
);

CKINVDCx20_ASAP7_75t_R g5847 ( 
.A(n_790),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_4714),
.Y(n_5848)
);

BUFx3_ASAP7_75t_L g5849 ( 
.A(n_4255),
.Y(n_5849)
);

CKINVDCx5p33_ASAP7_75t_R g5850 ( 
.A(n_749),
.Y(n_5850)
);

CKINVDCx5p33_ASAP7_75t_R g5851 ( 
.A(n_3149),
.Y(n_5851)
);

CKINVDCx20_ASAP7_75t_R g5852 ( 
.A(n_576),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_4957),
.Y(n_5853)
);

CKINVDCx5p33_ASAP7_75t_R g5854 ( 
.A(n_4784),
.Y(n_5854)
);

INVx1_ASAP7_75t_SL g5855 ( 
.A(n_4175),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_4599),
.Y(n_5856)
);

CKINVDCx5p33_ASAP7_75t_R g5857 ( 
.A(n_1493),
.Y(n_5857)
);

CKINVDCx5p33_ASAP7_75t_R g5858 ( 
.A(n_2127),
.Y(n_5858)
);

CKINVDCx5p33_ASAP7_75t_R g5859 ( 
.A(n_1223),
.Y(n_5859)
);

CKINVDCx5p33_ASAP7_75t_R g5860 ( 
.A(n_2018),
.Y(n_5860)
);

CKINVDCx5p33_ASAP7_75t_R g5861 ( 
.A(n_4319),
.Y(n_5861)
);

INVx1_ASAP7_75t_L g5862 ( 
.A(n_767),
.Y(n_5862)
);

CKINVDCx5p33_ASAP7_75t_R g5863 ( 
.A(n_3495),
.Y(n_5863)
);

INVx2_ASAP7_75t_L g5864 ( 
.A(n_4172),
.Y(n_5864)
);

CKINVDCx5p33_ASAP7_75t_R g5865 ( 
.A(n_4891),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_1427),
.Y(n_5866)
);

CKINVDCx5p33_ASAP7_75t_R g5867 ( 
.A(n_1329),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_3788),
.Y(n_5868)
);

CKINVDCx5p33_ASAP7_75t_R g5869 ( 
.A(n_1382),
.Y(n_5869)
);

CKINVDCx20_ASAP7_75t_R g5870 ( 
.A(n_2871),
.Y(n_5870)
);

CKINVDCx5p33_ASAP7_75t_R g5871 ( 
.A(n_3180),
.Y(n_5871)
);

INVx1_ASAP7_75t_L g5872 ( 
.A(n_1240),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_2157),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_3329),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_4391),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_4309),
.Y(n_5876)
);

CKINVDCx5p33_ASAP7_75t_R g5877 ( 
.A(n_4529),
.Y(n_5877)
);

CKINVDCx5p33_ASAP7_75t_R g5878 ( 
.A(n_289),
.Y(n_5878)
);

CKINVDCx5p33_ASAP7_75t_R g5879 ( 
.A(n_2339),
.Y(n_5879)
);

CKINVDCx5p33_ASAP7_75t_R g5880 ( 
.A(n_1511),
.Y(n_5880)
);

INVx1_ASAP7_75t_L g5881 ( 
.A(n_3258),
.Y(n_5881)
);

CKINVDCx5p33_ASAP7_75t_R g5882 ( 
.A(n_2523),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_4619),
.Y(n_5883)
);

CKINVDCx5p33_ASAP7_75t_R g5884 ( 
.A(n_1154),
.Y(n_5884)
);

CKINVDCx5p33_ASAP7_75t_R g5885 ( 
.A(n_2755),
.Y(n_5885)
);

BUFx10_ASAP7_75t_L g5886 ( 
.A(n_3429),
.Y(n_5886)
);

INVx1_ASAP7_75t_L g5887 ( 
.A(n_4997),
.Y(n_5887)
);

CKINVDCx5p33_ASAP7_75t_R g5888 ( 
.A(n_1631),
.Y(n_5888)
);

INVx1_ASAP7_75t_L g5889 ( 
.A(n_1485),
.Y(n_5889)
);

INVx1_ASAP7_75t_SL g5890 ( 
.A(n_3509),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_4211),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_4169),
.Y(n_5892)
);

INVx1_ASAP7_75t_SL g5893 ( 
.A(n_4288),
.Y(n_5893)
);

CKINVDCx5p33_ASAP7_75t_R g5894 ( 
.A(n_4208),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_2219),
.Y(n_5895)
);

CKINVDCx5p33_ASAP7_75t_R g5896 ( 
.A(n_567),
.Y(n_5896)
);

CKINVDCx5p33_ASAP7_75t_R g5897 ( 
.A(n_1838),
.Y(n_5897)
);

CKINVDCx5p33_ASAP7_75t_R g5898 ( 
.A(n_2180),
.Y(n_5898)
);

CKINVDCx5p33_ASAP7_75t_R g5899 ( 
.A(n_1946),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_3807),
.Y(n_5900)
);

INVx1_ASAP7_75t_SL g5901 ( 
.A(n_2136),
.Y(n_5901)
);

CKINVDCx5p33_ASAP7_75t_R g5902 ( 
.A(n_1106),
.Y(n_5902)
);

CKINVDCx5p33_ASAP7_75t_R g5903 ( 
.A(n_2873),
.Y(n_5903)
);

CKINVDCx5p33_ASAP7_75t_R g5904 ( 
.A(n_2961),
.Y(n_5904)
);

CKINVDCx5p33_ASAP7_75t_R g5905 ( 
.A(n_1173),
.Y(n_5905)
);

BUFx6f_ASAP7_75t_L g5906 ( 
.A(n_3413),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_2974),
.Y(n_5907)
);

CKINVDCx5p33_ASAP7_75t_R g5908 ( 
.A(n_2740),
.Y(n_5908)
);

CKINVDCx5p33_ASAP7_75t_R g5909 ( 
.A(n_2751),
.Y(n_5909)
);

CKINVDCx20_ASAP7_75t_R g5910 ( 
.A(n_3207),
.Y(n_5910)
);

CKINVDCx5p33_ASAP7_75t_R g5911 ( 
.A(n_3911),
.Y(n_5911)
);

CKINVDCx5p33_ASAP7_75t_R g5912 ( 
.A(n_4165),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_2316),
.Y(n_5913)
);

CKINVDCx5p33_ASAP7_75t_R g5914 ( 
.A(n_471),
.Y(n_5914)
);

INVx2_ASAP7_75t_L g5915 ( 
.A(n_2086),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_3712),
.Y(n_5916)
);

CKINVDCx5p33_ASAP7_75t_R g5917 ( 
.A(n_1610),
.Y(n_5917)
);

CKINVDCx5p33_ASAP7_75t_R g5918 ( 
.A(n_40),
.Y(n_5918)
);

CKINVDCx5p33_ASAP7_75t_R g5919 ( 
.A(n_4381),
.Y(n_5919)
);

CKINVDCx5p33_ASAP7_75t_R g5920 ( 
.A(n_2424),
.Y(n_5920)
);

CKINVDCx5p33_ASAP7_75t_R g5921 ( 
.A(n_2292),
.Y(n_5921)
);

INVx2_ASAP7_75t_L g5922 ( 
.A(n_2148),
.Y(n_5922)
);

CKINVDCx5p33_ASAP7_75t_R g5923 ( 
.A(n_1196),
.Y(n_5923)
);

CKINVDCx5p33_ASAP7_75t_R g5924 ( 
.A(n_3742),
.Y(n_5924)
);

CKINVDCx20_ASAP7_75t_R g5925 ( 
.A(n_156),
.Y(n_5925)
);

INVx2_ASAP7_75t_SL g5926 ( 
.A(n_25),
.Y(n_5926)
);

CKINVDCx5p33_ASAP7_75t_R g5927 ( 
.A(n_883),
.Y(n_5927)
);

CKINVDCx5p33_ASAP7_75t_R g5928 ( 
.A(n_4868),
.Y(n_5928)
);

INVx1_ASAP7_75t_L g5929 ( 
.A(n_179),
.Y(n_5929)
);

CKINVDCx20_ASAP7_75t_R g5930 ( 
.A(n_2265),
.Y(n_5930)
);

CKINVDCx20_ASAP7_75t_R g5931 ( 
.A(n_4729),
.Y(n_5931)
);

INVx1_ASAP7_75t_L g5932 ( 
.A(n_4702),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_1902),
.Y(n_5933)
);

CKINVDCx20_ASAP7_75t_R g5934 ( 
.A(n_4277),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_1144),
.Y(n_5935)
);

INVx1_ASAP7_75t_L g5936 ( 
.A(n_4294),
.Y(n_5936)
);

CKINVDCx5p33_ASAP7_75t_R g5937 ( 
.A(n_4564),
.Y(n_5937)
);

INVx1_ASAP7_75t_L g5938 ( 
.A(n_4098),
.Y(n_5938)
);

BUFx3_ASAP7_75t_L g5939 ( 
.A(n_838),
.Y(n_5939)
);

CKINVDCx5p33_ASAP7_75t_R g5940 ( 
.A(n_444),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_2759),
.Y(n_5941)
);

CKINVDCx5p33_ASAP7_75t_R g5942 ( 
.A(n_545),
.Y(n_5942)
);

BUFx6f_ASAP7_75t_L g5943 ( 
.A(n_4444),
.Y(n_5943)
);

CKINVDCx20_ASAP7_75t_R g5944 ( 
.A(n_57),
.Y(n_5944)
);

CKINVDCx5p33_ASAP7_75t_R g5945 ( 
.A(n_4217),
.Y(n_5945)
);

INVx1_ASAP7_75t_L g5946 ( 
.A(n_874),
.Y(n_5946)
);

INVx1_ASAP7_75t_L g5947 ( 
.A(n_2252),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_3899),
.Y(n_5948)
);

CKINVDCx5p33_ASAP7_75t_R g5949 ( 
.A(n_2738),
.Y(n_5949)
);

CKINVDCx5p33_ASAP7_75t_R g5950 ( 
.A(n_4656),
.Y(n_5950)
);

BUFx6f_ASAP7_75t_L g5951 ( 
.A(n_4068),
.Y(n_5951)
);

CKINVDCx5p33_ASAP7_75t_R g5952 ( 
.A(n_1630),
.Y(n_5952)
);

CKINVDCx5p33_ASAP7_75t_R g5953 ( 
.A(n_4666),
.Y(n_5953)
);

CKINVDCx5p33_ASAP7_75t_R g5954 ( 
.A(n_4833),
.Y(n_5954)
);

CKINVDCx5p33_ASAP7_75t_R g5955 ( 
.A(n_4295),
.Y(n_5955)
);

INVx2_ASAP7_75t_L g5956 ( 
.A(n_2173),
.Y(n_5956)
);

INVx1_ASAP7_75t_SL g5957 ( 
.A(n_4174),
.Y(n_5957)
);

CKINVDCx5p33_ASAP7_75t_R g5958 ( 
.A(n_38),
.Y(n_5958)
);

INVx1_ASAP7_75t_L g5959 ( 
.A(n_4210),
.Y(n_5959)
);

BUFx2_ASAP7_75t_R g5960 ( 
.A(n_2582),
.Y(n_5960)
);

INVxp67_ASAP7_75t_L g5961 ( 
.A(n_2019),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_4270),
.Y(n_5962)
);

CKINVDCx5p33_ASAP7_75t_R g5963 ( 
.A(n_1513),
.Y(n_5963)
);

CKINVDCx5p33_ASAP7_75t_R g5964 ( 
.A(n_3675),
.Y(n_5964)
);

CKINVDCx5p33_ASAP7_75t_R g5965 ( 
.A(n_2820),
.Y(n_5965)
);

INVx1_ASAP7_75t_L g5966 ( 
.A(n_1466),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_3406),
.Y(n_5967)
);

CKINVDCx5p33_ASAP7_75t_R g5968 ( 
.A(n_1786),
.Y(n_5968)
);

CKINVDCx5p33_ASAP7_75t_R g5969 ( 
.A(n_1930),
.Y(n_5969)
);

CKINVDCx5p33_ASAP7_75t_R g5970 ( 
.A(n_199),
.Y(n_5970)
);

CKINVDCx5p33_ASAP7_75t_R g5971 ( 
.A(n_275),
.Y(n_5971)
);

CKINVDCx20_ASAP7_75t_R g5972 ( 
.A(n_4026),
.Y(n_5972)
);

CKINVDCx20_ASAP7_75t_R g5973 ( 
.A(n_4436),
.Y(n_5973)
);

BUFx3_ASAP7_75t_L g5974 ( 
.A(n_1110),
.Y(n_5974)
);

BUFx3_ASAP7_75t_L g5975 ( 
.A(n_1122),
.Y(n_5975)
);

INVx1_ASAP7_75t_L g5976 ( 
.A(n_2635),
.Y(n_5976)
);

CKINVDCx5p33_ASAP7_75t_R g5977 ( 
.A(n_4814),
.Y(n_5977)
);

CKINVDCx5p33_ASAP7_75t_R g5978 ( 
.A(n_4604),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_4275),
.Y(n_5979)
);

CKINVDCx5p33_ASAP7_75t_R g5980 ( 
.A(n_3999),
.Y(n_5980)
);

CKINVDCx5p33_ASAP7_75t_R g5981 ( 
.A(n_1350),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_4512),
.Y(n_5982)
);

CKINVDCx5p33_ASAP7_75t_R g5983 ( 
.A(n_1045),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_4222),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_3534),
.Y(n_5985)
);

INVx2_ASAP7_75t_L g5986 ( 
.A(n_682),
.Y(n_5986)
);

CKINVDCx5p33_ASAP7_75t_R g5987 ( 
.A(n_258),
.Y(n_5987)
);

INVx1_ASAP7_75t_SL g5988 ( 
.A(n_906),
.Y(n_5988)
);

CKINVDCx5p33_ASAP7_75t_R g5989 ( 
.A(n_3107),
.Y(n_5989)
);

CKINVDCx5p33_ASAP7_75t_R g5990 ( 
.A(n_2628),
.Y(n_5990)
);

CKINVDCx5p33_ASAP7_75t_R g5991 ( 
.A(n_2776),
.Y(n_5991)
);

CKINVDCx5p33_ASAP7_75t_R g5992 ( 
.A(n_1441),
.Y(n_5992)
);

INVx2_ASAP7_75t_L g5993 ( 
.A(n_4275),
.Y(n_5993)
);

CKINVDCx5p33_ASAP7_75t_R g5994 ( 
.A(n_1874),
.Y(n_5994)
);

BUFx2_ASAP7_75t_L g5995 ( 
.A(n_2736),
.Y(n_5995)
);

CKINVDCx5p33_ASAP7_75t_R g5996 ( 
.A(n_1060),
.Y(n_5996)
);

INVx1_ASAP7_75t_L g5997 ( 
.A(n_3575),
.Y(n_5997)
);

BUFx2_ASAP7_75t_L g5998 ( 
.A(n_1309),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_2483),
.Y(n_5999)
);

CKINVDCx5p33_ASAP7_75t_R g6000 ( 
.A(n_4563),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_3775),
.Y(n_6001)
);

BUFx6f_ASAP7_75t_L g6002 ( 
.A(n_964),
.Y(n_6002)
);

CKINVDCx5p33_ASAP7_75t_R g6003 ( 
.A(n_4141),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_3674),
.Y(n_6004)
);

INVx1_ASAP7_75t_L g6005 ( 
.A(n_3829),
.Y(n_6005)
);

CKINVDCx5p33_ASAP7_75t_R g6006 ( 
.A(n_4807),
.Y(n_6006)
);

INVx1_ASAP7_75t_SL g6007 ( 
.A(n_738),
.Y(n_6007)
);

INVx2_ASAP7_75t_L g6008 ( 
.A(n_485),
.Y(n_6008)
);

CKINVDCx20_ASAP7_75t_R g6009 ( 
.A(n_3775),
.Y(n_6009)
);

CKINVDCx5p33_ASAP7_75t_R g6010 ( 
.A(n_1944),
.Y(n_6010)
);

CKINVDCx5p33_ASAP7_75t_R g6011 ( 
.A(n_4555),
.Y(n_6011)
);

CKINVDCx5p33_ASAP7_75t_R g6012 ( 
.A(n_2281),
.Y(n_6012)
);

INVx1_ASAP7_75t_L g6013 ( 
.A(n_2136),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_4284),
.Y(n_6014)
);

INVx1_ASAP7_75t_L g6015 ( 
.A(n_3819),
.Y(n_6015)
);

INVx2_ASAP7_75t_L g6016 ( 
.A(n_4267),
.Y(n_6016)
);

CKINVDCx5p33_ASAP7_75t_R g6017 ( 
.A(n_4186),
.Y(n_6017)
);

CKINVDCx5p33_ASAP7_75t_R g6018 ( 
.A(n_1190),
.Y(n_6018)
);

CKINVDCx5p33_ASAP7_75t_R g6019 ( 
.A(n_4803),
.Y(n_6019)
);

HB1xp67_ASAP7_75t_L g6020 ( 
.A(n_4383),
.Y(n_6020)
);

CKINVDCx14_ASAP7_75t_R g6021 ( 
.A(n_4266),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_3598),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_2898),
.Y(n_6023)
);

BUFx8_ASAP7_75t_SL g6024 ( 
.A(n_769),
.Y(n_6024)
);

CKINVDCx5p33_ASAP7_75t_R g6025 ( 
.A(n_4195),
.Y(n_6025)
);

CKINVDCx5p33_ASAP7_75t_R g6026 ( 
.A(n_4185),
.Y(n_6026)
);

INVx2_ASAP7_75t_L g6027 ( 
.A(n_2244),
.Y(n_6027)
);

CKINVDCx5p33_ASAP7_75t_R g6028 ( 
.A(n_830),
.Y(n_6028)
);

INVx1_ASAP7_75t_SL g6029 ( 
.A(n_91),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_2309),
.Y(n_6030)
);

CKINVDCx5p33_ASAP7_75t_R g6031 ( 
.A(n_3645),
.Y(n_6031)
);

CKINVDCx5p33_ASAP7_75t_R g6032 ( 
.A(n_4440),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_165),
.Y(n_6033)
);

CKINVDCx5p33_ASAP7_75t_R g6034 ( 
.A(n_3314),
.Y(n_6034)
);

CKINVDCx20_ASAP7_75t_R g6035 ( 
.A(n_4307),
.Y(n_6035)
);

INVx1_ASAP7_75t_L g6036 ( 
.A(n_2660),
.Y(n_6036)
);

INVx2_ASAP7_75t_SL g6037 ( 
.A(n_3804),
.Y(n_6037)
);

CKINVDCx5p33_ASAP7_75t_R g6038 ( 
.A(n_1942),
.Y(n_6038)
);

INVx1_ASAP7_75t_L g6039 ( 
.A(n_2575),
.Y(n_6039)
);

CKINVDCx5p33_ASAP7_75t_R g6040 ( 
.A(n_2589),
.Y(n_6040)
);

CKINVDCx5p33_ASAP7_75t_R g6041 ( 
.A(n_253),
.Y(n_6041)
);

BUFx3_ASAP7_75t_L g6042 ( 
.A(n_3668),
.Y(n_6042)
);

INVx1_ASAP7_75t_L g6043 ( 
.A(n_4179),
.Y(n_6043)
);

CKINVDCx5p33_ASAP7_75t_R g6044 ( 
.A(n_3343),
.Y(n_6044)
);

CKINVDCx20_ASAP7_75t_R g6045 ( 
.A(n_3909),
.Y(n_6045)
);

CKINVDCx5p33_ASAP7_75t_R g6046 ( 
.A(n_2890),
.Y(n_6046)
);

BUFx10_ASAP7_75t_L g6047 ( 
.A(n_1046),
.Y(n_6047)
);

CKINVDCx5p33_ASAP7_75t_R g6048 ( 
.A(n_2878),
.Y(n_6048)
);

CKINVDCx5p33_ASAP7_75t_R g6049 ( 
.A(n_2967),
.Y(n_6049)
);

INVx2_ASAP7_75t_L g6050 ( 
.A(n_764),
.Y(n_6050)
);

INVx1_ASAP7_75t_L g6051 ( 
.A(n_4236),
.Y(n_6051)
);

CKINVDCx5p33_ASAP7_75t_R g6052 ( 
.A(n_3175),
.Y(n_6052)
);

INVx1_ASAP7_75t_L g6053 ( 
.A(n_826),
.Y(n_6053)
);

CKINVDCx5p33_ASAP7_75t_R g6054 ( 
.A(n_4507),
.Y(n_6054)
);

INVx2_ASAP7_75t_L g6055 ( 
.A(n_3942),
.Y(n_6055)
);

INVx1_ASAP7_75t_SL g6056 ( 
.A(n_3888),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_4163),
.Y(n_6057)
);

CKINVDCx5p33_ASAP7_75t_R g6058 ( 
.A(n_1438),
.Y(n_6058)
);

INVx2_ASAP7_75t_L g6059 ( 
.A(n_1827),
.Y(n_6059)
);

CKINVDCx5p33_ASAP7_75t_R g6060 ( 
.A(n_4229),
.Y(n_6060)
);

CKINVDCx5p33_ASAP7_75t_R g6061 ( 
.A(n_1554),
.Y(n_6061)
);

CKINVDCx5p33_ASAP7_75t_R g6062 ( 
.A(n_571),
.Y(n_6062)
);

CKINVDCx5p33_ASAP7_75t_R g6063 ( 
.A(n_4206),
.Y(n_6063)
);

CKINVDCx5p33_ASAP7_75t_R g6064 ( 
.A(n_3667),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_4194),
.Y(n_6065)
);

INVx1_ASAP7_75t_L g6066 ( 
.A(n_1048),
.Y(n_6066)
);

INVx1_ASAP7_75t_L g6067 ( 
.A(n_4124),
.Y(n_6067)
);

INVxp67_ASAP7_75t_L g6068 ( 
.A(n_4296),
.Y(n_6068)
);

INVx1_ASAP7_75t_L g6069 ( 
.A(n_4745),
.Y(n_6069)
);

INVx1_ASAP7_75t_L g6070 ( 
.A(n_141),
.Y(n_6070)
);

INVx2_ASAP7_75t_SL g6071 ( 
.A(n_3176),
.Y(n_6071)
);

BUFx2_ASAP7_75t_L g6072 ( 
.A(n_295),
.Y(n_6072)
);

CKINVDCx5p33_ASAP7_75t_R g6073 ( 
.A(n_990),
.Y(n_6073)
);

CKINVDCx20_ASAP7_75t_R g6074 ( 
.A(n_2520),
.Y(n_6074)
);

BUFx5_ASAP7_75t_L g6075 ( 
.A(n_637),
.Y(n_6075)
);

CKINVDCx5p33_ASAP7_75t_R g6076 ( 
.A(n_3487),
.Y(n_6076)
);

INVx1_ASAP7_75t_L g6077 ( 
.A(n_4183),
.Y(n_6077)
);

INVx1_ASAP7_75t_L g6078 ( 
.A(n_3223),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_21),
.Y(n_6079)
);

INVx2_ASAP7_75t_L g6080 ( 
.A(n_2787),
.Y(n_6080)
);

INVx1_ASAP7_75t_SL g6081 ( 
.A(n_2938),
.Y(n_6081)
);

CKINVDCx16_ASAP7_75t_R g6082 ( 
.A(n_3490),
.Y(n_6082)
);

INVx2_ASAP7_75t_L g6083 ( 
.A(n_2586),
.Y(n_6083)
);

CKINVDCx20_ASAP7_75t_R g6084 ( 
.A(n_1314),
.Y(n_6084)
);

BUFx3_ASAP7_75t_L g6085 ( 
.A(n_4065),
.Y(n_6085)
);

CKINVDCx5p33_ASAP7_75t_R g6086 ( 
.A(n_5006),
.Y(n_6086)
);

BUFx10_ASAP7_75t_L g6087 ( 
.A(n_1108),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_904),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_1320),
.Y(n_6089)
);

CKINVDCx5p33_ASAP7_75t_R g6090 ( 
.A(n_449),
.Y(n_6090)
);

BUFx6f_ASAP7_75t_L g6091 ( 
.A(n_2165),
.Y(n_6091)
);

INVx2_ASAP7_75t_L g6092 ( 
.A(n_4749),
.Y(n_6092)
);

CKINVDCx5p33_ASAP7_75t_R g6093 ( 
.A(n_4129),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_855),
.Y(n_6094)
);

CKINVDCx5p33_ASAP7_75t_R g6095 ( 
.A(n_528),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_3087),
.Y(n_6096)
);

CKINVDCx5p33_ASAP7_75t_R g6097 ( 
.A(n_4177),
.Y(n_6097)
);

INVx2_ASAP7_75t_L g6098 ( 
.A(n_210),
.Y(n_6098)
);

INVx1_ASAP7_75t_L g6099 ( 
.A(n_3338),
.Y(n_6099)
);

BUFx3_ASAP7_75t_L g6100 ( 
.A(n_2191),
.Y(n_6100)
);

INVx1_ASAP7_75t_L g6101 ( 
.A(n_2101),
.Y(n_6101)
);

INVx1_ASAP7_75t_SL g6102 ( 
.A(n_3497),
.Y(n_6102)
);

CKINVDCx5p33_ASAP7_75t_R g6103 ( 
.A(n_4188),
.Y(n_6103)
);

CKINVDCx20_ASAP7_75t_R g6104 ( 
.A(n_1806),
.Y(n_6104)
);

INVx1_ASAP7_75t_SL g6105 ( 
.A(n_3198),
.Y(n_6105)
);

BUFx10_ASAP7_75t_L g6106 ( 
.A(n_916),
.Y(n_6106)
);

INVx1_ASAP7_75t_L g6107 ( 
.A(n_4205),
.Y(n_6107)
);

INVx1_ASAP7_75t_L g6108 ( 
.A(n_864),
.Y(n_6108)
);

CKINVDCx5p33_ASAP7_75t_R g6109 ( 
.A(n_4247),
.Y(n_6109)
);

CKINVDCx20_ASAP7_75t_R g6110 ( 
.A(n_2549),
.Y(n_6110)
);

INVx1_ASAP7_75t_SL g6111 ( 
.A(n_4647),
.Y(n_6111)
);

CKINVDCx5p33_ASAP7_75t_R g6112 ( 
.A(n_4237),
.Y(n_6112)
);

INVx1_ASAP7_75t_L g6113 ( 
.A(n_1417),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_4257),
.Y(n_6114)
);

INVx1_ASAP7_75t_SL g6115 ( 
.A(n_1470),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_2382),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_4681),
.Y(n_6117)
);

CKINVDCx5p33_ASAP7_75t_R g6118 ( 
.A(n_3122),
.Y(n_6118)
);

CKINVDCx20_ASAP7_75t_R g6119 ( 
.A(n_1702),
.Y(n_6119)
);

INVx1_ASAP7_75t_SL g6120 ( 
.A(n_3838),
.Y(n_6120)
);

INVx1_ASAP7_75t_L g6121 ( 
.A(n_639),
.Y(n_6121)
);

CKINVDCx5p33_ASAP7_75t_R g6122 ( 
.A(n_4283),
.Y(n_6122)
);

CKINVDCx5p33_ASAP7_75t_R g6123 ( 
.A(n_1821),
.Y(n_6123)
);

CKINVDCx5p33_ASAP7_75t_R g6124 ( 
.A(n_1720),
.Y(n_6124)
);

INVx1_ASAP7_75t_L g6125 ( 
.A(n_3453),
.Y(n_6125)
);

CKINVDCx5p33_ASAP7_75t_R g6126 ( 
.A(n_149),
.Y(n_6126)
);

CKINVDCx5p33_ASAP7_75t_R g6127 ( 
.A(n_4475),
.Y(n_6127)
);

CKINVDCx5p33_ASAP7_75t_R g6128 ( 
.A(n_2321),
.Y(n_6128)
);

INVx1_ASAP7_75t_L g6129 ( 
.A(n_4292),
.Y(n_6129)
);

CKINVDCx5p33_ASAP7_75t_R g6130 ( 
.A(n_4251),
.Y(n_6130)
);

CKINVDCx5p33_ASAP7_75t_R g6131 ( 
.A(n_3570),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_542),
.Y(n_6132)
);

CKINVDCx20_ASAP7_75t_R g6133 ( 
.A(n_2579),
.Y(n_6133)
);

HB1xp67_ASAP7_75t_L g6134 ( 
.A(n_4123),
.Y(n_6134)
);

INVx1_ASAP7_75t_L g6135 ( 
.A(n_4550),
.Y(n_6135)
);

CKINVDCx5p33_ASAP7_75t_R g6136 ( 
.A(n_2892),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_4248),
.Y(n_6137)
);

CKINVDCx5p33_ASAP7_75t_R g6138 ( 
.A(n_3502),
.Y(n_6138)
);

CKINVDCx5p33_ASAP7_75t_R g6139 ( 
.A(n_4071),
.Y(n_6139)
);

CKINVDCx5p33_ASAP7_75t_R g6140 ( 
.A(n_3164),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_1004),
.Y(n_6141)
);

INVx1_ASAP7_75t_SL g6142 ( 
.A(n_236),
.Y(n_6142)
);

CKINVDCx5p33_ASAP7_75t_R g6143 ( 
.A(n_4203),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_3256),
.Y(n_6144)
);

CKINVDCx5p33_ASAP7_75t_R g6145 ( 
.A(n_1105),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_1011),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_2504),
.Y(n_6147)
);

CKINVDCx5p33_ASAP7_75t_R g6148 ( 
.A(n_907),
.Y(n_6148)
);

CKINVDCx5p33_ASAP7_75t_R g6149 ( 
.A(n_921),
.Y(n_6149)
);

CKINVDCx5p33_ASAP7_75t_R g6150 ( 
.A(n_2257),
.Y(n_6150)
);

CKINVDCx16_ASAP7_75t_R g6151 ( 
.A(n_4882),
.Y(n_6151)
);

CKINVDCx5p33_ASAP7_75t_R g6152 ( 
.A(n_456),
.Y(n_6152)
);

BUFx5_ASAP7_75t_L g6153 ( 
.A(n_4285),
.Y(n_6153)
);

INVx1_ASAP7_75t_L g6154 ( 
.A(n_3118),
.Y(n_6154)
);

INVx1_ASAP7_75t_L g6155 ( 
.A(n_1159),
.Y(n_6155)
);

CKINVDCx20_ASAP7_75t_R g6156 ( 
.A(n_4991),
.Y(n_6156)
);

CKINVDCx5p33_ASAP7_75t_R g6157 ( 
.A(n_2131),
.Y(n_6157)
);

CKINVDCx5p33_ASAP7_75t_R g6158 ( 
.A(n_3388),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_4202),
.Y(n_6159)
);

CKINVDCx20_ASAP7_75t_R g6160 ( 
.A(n_1904),
.Y(n_6160)
);

BUFx8_ASAP7_75t_SL g6161 ( 
.A(n_2160),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_57),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_2253),
.Y(n_6163)
);

INVx1_ASAP7_75t_L g6164 ( 
.A(n_2124),
.Y(n_6164)
);

CKINVDCx5p33_ASAP7_75t_R g6165 ( 
.A(n_3682),
.Y(n_6165)
);

CKINVDCx5p33_ASAP7_75t_R g6166 ( 
.A(n_2583),
.Y(n_6166)
);

CKINVDCx5p33_ASAP7_75t_R g6167 ( 
.A(n_918),
.Y(n_6167)
);

CKINVDCx5p33_ASAP7_75t_R g6168 ( 
.A(n_4091),
.Y(n_6168)
);

BUFx5_ASAP7_75t_L g6169 ( 
.A(n_1978),
.Y(n_6169)
);

CKINVDCx5p33_ASAP7_75t_R g6170 ( 
.A(n_1577),
.Y(n_6170)
);

INVx1_ASAP7_75t_SL g6171 ( 
.A(n_1165),
.Y(n_6171)
);

BUFx10_ASAP7_75t_L g6172 ( 
.A(n_1607),
.Y(n_6172)
);

CKINVDCx5p33_ASAP7_75t_R g6173 ( 
.A(n_3842),
.Y(n_6173)
);

CKINVDCx5p33_ASAP7_75t_R g6174 ( 
.A(n_706),
.Y(n_6174)
);

CKINVDCx5p33_ASAP7_75t_R g6175 ( 
.A(n_2790),
.Y(n_6175)
);

CKINVDCx5p33_ASAP7_75t_R g6176 ( 
.A(n_3973),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_636),
.Y(n_6177)
);

CKINVDCx5p33_ASAP7_75t_R g6178 ( 
.A(n_4168),
.Y(n_6178)
);

BUFx2_ASAP7_75t_L g6179 ( 
.A(n_337),
.Y(n_6179)
);

CKINVDCx5p33_ASAP7_75t_R g6180 ( 
.A(n_1283),
.Y(n_6180)
);

CKINVDCx20_ASAP7_75t_R g6181 ( 
.A(n_3316),
.Y(n_6181)
);

CKINVDCx5p33_ASAP7_75t_R g6182 ( 
.A(n_1171),
.Y(n_6182)
);

CKINVDCx5p33_ASAP7_75t_R g6183 ( 
.A(n_2886),
.Y(n_6183)
);

INVx1_ASAP7_75t_L g6184 ( 
.A(n_1790),
.Y(n_6184)
);

INVx1_ASAP7_75t_L g6185 ( 
.A(n_3665),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_3752),
.Y(n_6186)
);

INVx1_ASAP7_75t_L g6187 ( 
.A(n_2269),
.Y(n_6187)
);

CKINVDCx5p33_ASAP7_75t_R g6188 ( 
.A(n_2714),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_4064),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_1634),
.Y(n_6190)
);

CKINVDCx5p33_ASAP7_75t_R g6191 ( 
.A(n_910),
.Y(n_6191)
);

INVx1_ASAP7_75t_L g6192 ( 
.A(n_3575),
.Y(n_6192)
);

CKINVDCx16_ASAP7_75t_R g6193 ( 
.A(n_2544),
.Y(n_6193)
);

INVx1_ASAP7_75t_L g6194 ( 
.A(n_3958),
.Y(n_6194)
);

CKINVDCx16_ASAP7_75t_R g6195 ( 
.A(n_3530),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_3353),
.Y(n_6196)
);

CKINVDCx5p33_ASAP7_75t_R g6197 ( 
.A(n_1172),
.Y(n_6197)
);

INVx2_ASAP7_75t_L g6198 ( 
.A(n_4184),
.Y(n_6198)
);

INVx1_ASAP7_75t_L g6199 ( 
.A(n_404),
.Y(n_6199)
);

INVx1_ASAP7_75t_L g6200 ( 
.A(n_3278),
.Y(n_6200)
);

CKINVDCx5p33_ASAP7_75t_R g6201 ( 
.A(n_2927),
.Y(n_6201)
);

CKINVDCx5p33_ASAP7_75t_R g6202 ( 
.A(n_5024),
.Y(n_6202)
);

CKINVDCx5p33_ASAP7_75t_R g6203 ( 
.A(n_3857),
.Y(n_6203)
);

INVx2_ASAP7_75t_L g6204 ( 
.A(n_4279),
.Y(n_6204)
);

CKINVDCx20_ASAP7_75t_R g6205 ( 
.A(n_623),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_600),
.Y(n_6206)
);

INVx2_ASAP7_75t_L g6207 ( 
.A(n_2613),
.Y(n_6207)
);

CKINVDCx5p33_ASAP7_75t_R g6208 ( 
.A(n_1532),
.Y(n_6208)
);

BUFx5_ASAP7_75t_L g6209 ( 
.A(n_1159),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_688),
.Y(n_6210)
);

BUFx10_ASAP7_75t_L g6211 ( 
.A(n_3572),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_4216),
.Y(n_6212)
);

INVx1_ASAP7_75t_L g6213 ( 
.A(n_1683),
.Y(n_6213)
);

INVx1_ASAP7_75t_L g6214 ( 
.A(n_4213),
.Y(n_6214)
);

CKINVDCx5p33_ASAP7_75t_R g6215 ( 
.A(n_295),
.Y(n_6215)
);

CKINVDCx5p33_ASAP7_75t_R g6216 ( 
.A(n_308),
.Y(n_6216)
);

CKINVDCx5p33_ASAP7_75t_R g6217 ( 
.A(n_2399),
.Y(n_6217)
);

BUFx3_ASAP7_75t_L g6218 ( 
.A(n_3374),
.Y(n_6218)
);

CKINVDCx5p33_ASAP7_75t_R g6219 ( 
.A(n_1499),
.Y(n_6219)
);

CKINVDCx5p33_ASAP7_75t_R g6220 ( 
.A(n_4553),
.Y(n_6220)
);

CKINVDCx5p33_ASAP7_75t_R g6221 ( 
.A(n_4252),
.Y(n_6221)
);

CKINVDCx5p33_ASAP7_75t_R g6222 ( 
.A(n_2790),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_2784),
.Y(n_6223)
);

INVx1_ASAP7_75t_L g6224 ( 
.A(n_3870),
.Y(n_6224)
);

CKINVDCx5p33_ASAP7_75t_R g6225 ( 
.A(n_4170),
.Y(n_6225)
);

CKINVDCx5p33_ASAP7_75t_R g6226 ( 
.A(n_4209),
.Y(n_6226)
);

INVx1_ASAP7_75t_L g6227 ( 
.A(n_1755),
.Y(n_6227)
);

CKINVDCx5p33_ASAP7_75t_R g6228 ( 
.A(n_4218),
.Y(n_6228)
);

INVx1_ASAP7_75t_L g6229 ( 
.A(n_3296),
.Y(n_6229)
);

CKINVDCx5p33_ASAP7_75t_R g6230 ( 
.A(n_4810),
.Y(n_6230)
);

INVx1_ASAP7_75t_L g6231 ( 
.A(n_4137),
.Y(n_6231)
);

CKINVDCx5p33_ASAP7_75t_R g6232 ( 
.A(n_3006),
.Y(n_6232)
);

CKINVDCx5p33_ASAP7_75t_R g6233 ( 
.A(n_111),
.Y(n_6233)
);

BUFx3_ASAP7_75t_L g6234 ( 
.A(n_423),
.Y(n_6234)
);

INVx1_ASAP7_75t_SL g6235 ( 
.A(n_3530),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_1476),
.Y(n_6236)
);

CKINVDCx5p33_ASAP7_75t_R g6237 ( 
.A(n_338),
.Y(n_6237)
);

INVx2_ASAP7_75t_SL g6238 ( 
.A(n_4237),
.Y(n_6238)
);

CKINVDCx20_ASAP7_75t_R g6239 ( 
.A(n_4293),
.Y(n_6239)
);

CKINVDCx5p33_ASAP7_75t_R g6240 ( 
.A(n_2273),
.Y(n_6240)
);

INVx2_ASAP7_75t_L g6241 ( 
.A(n_2933),
.Y(n_6241)
);

CKINVDCx5p33_ASAP7_75t_R g6242 ( 
.A(n_2812),
.Y(n_6242)
);

BUFx2_ASAP7_75t_L g6243 ( 
.A(n_4548),
.Y(n_6243)
);

INVx1_ASAP7_75t_L g6244 ( 
.A(n_4308),
.Y(n_6244)
);

CKINVDCx5p33_ASAP7_75t_R g6245 ( 
.A(n_2013),
.Y(n_6245)
);

CKINVDCx5p33_ASAP7_75t_R g6246 ( 
.A(n_2663),
.Y(n_6246)
);

INVx1_ASAP7_75t_L g6247 ( 
.A(n_1803),
.Y(n_6247)
);

CKINVDCx5p33_ASAP7_75t_R g6248 ( 
.A(n_1123),
.Y(n_6248)
);

CKINVDCx5p33_ASAP7_75t_R g6249 ( 
.A(n_812),
.Y(n_6249)
);

CKINVDCx16_ASAP7_75t_R g6250 ( 
.A(n_3068),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_3963),
.Y(n_6251)
);

CKINVDCx5p33_ASAP7_75t_R g6252 ( 
.A(n_3350),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_3262),
.Y(n_6253)
);

CKINVDCx5p33_ASAP7_75t_R g6254 ( 
.A(n_1747),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_2542),
.Y(n_6255)
);

CKINVDCx5p33_ASAP7_75t_R g6256 ( 
.A(n_222),
.Y(n_6256)
);

BUFx2_ASAP7_75t_L g6257 ( 
.A(n_3045),
.Y(n_6257)
);

CKINVDCx5p33_ASAP7_75t_R g6258 ( 
.A(n_1605),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_2180),
.Y(n_6259)
);

INVx1_ASAP7_75t_L g6260 ( 
.A(n_4999),
.Y(n_6260)
);

BUFx3_ASAP7_75t_L g6261 ( 
.A(n_4264),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_2185),
.Y(n_6262)
);

CKINVDCx5p33_ASAP7_75t_R g6263 ( 
.A(n_4994),
.Y(n_6263)
);

CKINVDCx16_ASAP7_75t_R g6264 ( 
.A(n_3679),
.Y(n_6264)
);

CKINVDCx5p33_ASAP7_75t_R g6265 ( 
.A(n_1055),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_872),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_4135),
.Y(n_6267)
);

INVx1_ASAP7_75t_L g6268 ( 
.A(n_278),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_3797),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_4823),
.Y(n_6270)
);

CKINVDCx5p33_ASAP7_75t_R g6271 ( 
.A(n_796),
.Y(n_6271)
);

CKINVDCx5p33_ASAP7_75t_R g6272 ( 
.A(n_1198),
.Y(n_6272)
);

CKINVDCx5p33_ASAP7_75t_R g6273 ( 
.A(n_4207),
.Y(n_6273)
);

CKINVDCx5p33_ASAP7_75t_R g6274 ( 
.A(n_1223),
.Y(n_6274)
);

CKINVDCx20_ASAP7_75t_R g6275 ( 
.A(n_3130),
.Y(n_6275)
);

CKINVDCx5p33_ASAP7_75t_R g6276 ( 
.A(n_4172),
.Y(n_6276)
);

CKINVDCx5p33_ASAP7_75t_R g6277 ( 
.A(n_1414),
.Y(n_6277)
);

CKINVDCx5p33_ASAP7_75t_R g6278 ( 
.A(n_1568),
.Y(n_6278)
);

CKINVDCx5p33_ASAP7_75t_R g6279 ( 
.A(n_3082),
.Y(n_6279)
);

BUFx6f_ASAP7_75t_L g6280 ( 
.A(n_54),
.Y(n_6280)
);

BUFx6f_ASAP7_75t_L g6281 ( 
.A(n_4718),
.Y(n_6281)
);

BUFx6f_ASAP7_75t_L g6282 ( 
.A(n_4225),
.Y(n_6282)
);

INVx1_ASAP7_75t_SL g6283 ( 
.A(n_2000),
.Y(n_6283)
);

INVx1_ASAP7_75t_L g6284 ( 
.A(n_3637),
.Y(n_6284)
);

CKINVDCx5p33_ASAP7_75t_R g6285 ( 
.A(n_2629),
.Y(n_6285)
);

CKINVDCx5p33_ASAP7_75t_R g6286 ( 
.A(n_2299),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_1462),
.Y(n_6287)
);

INVx2_ASAP7_75t_L g6288 ( 
.A(n_3738),
.Y(n_6288)
);

CKINVDCx5p33_ASAP7_75t_R g6289 ( 
.A(n_3168),
.Y(n_6289)
);

CKINVDCx5p33_ASAP7_75t_R g6290 ( 
.A(n_264),
.Y(n_6290)
);

INVx1_ASAP7_75t_L g6291 ( 
.A(n_5009),
.Y(n_6291)
);

CKINVDCx5p33_ASAP7_75t_R g6292 ( 
.A(n_1792),
.Y(n_6292)
);

CKINVDCx5p33_ASAP7_75t_R g6293 ( 
.A(n_2376),
.Y(n_6293)
);

CKINVDCx5p33_ASAP7_75t_R g6294 ( 
.A(n_3202),
.Y(n_6294)
);

BUFx3_ASAP7_75t_L g6295 ( 
.A(n_4989),
.Y(n_6295)
);

CKINVDCx5p33_ASAP7_75t_R g6296 ( 
.A(n_2511),
.Y(n_6296)
);

INVx2_ASAP7_75t_L g6297 ( 
.A(n_1714),
.Y(n_6297)
);

CKINVDCx20_ASAP7_75t_R g6298 ( 
.A(n_1724),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_4899),
.Y(n_6299)
);

CKINVDCx5p33_ASAP7_75t_R g6300 ( 
.A(n_736),
.Y(n_6300)
);

CKINVDCx20_ASAP7_75t_R g6301 ( 
.A(n_4265),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_2633),
.Y(n_6302)
);

CKINVDCx5p33_ASAP7_75t_R g6303 ( 
.A(n_3801),
.Y(n_6303)
);

CKINVDCx5p33_ASAP7_75t_R g6304 ( 
.A(n_3954),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_2677),
.Y(n_6305)
);

BUFx2_ASAP7_75t_L g6306 ( 
.A(n_773),
.Y(n_6306)
);

CKINVDCx20_ASAP7_75t_R g6307 ( 
.A(n_114),
.Y(n_6307)
);

CKINVDCx5p33_ASAP7_75t_R g6308 ( 
.A(n_5019),
.Y(n_6308)
);

CKINVDCx5p33_ASAP7_75t_R g6309 ( 
.A(n_200),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_933),
.Y(n_6310)
);

CKINVDCx5p33_ASAP7_75t_R g6311 ( 
.A(n_1911),
.Y(n_6311)
);

CKINVDCx5p33_ASAP7_75t_R g6312 ( 
.A(n_3687),
.Y(n_6312)
);

CKINVDCx16_ASAP7_75t_R g6313 ( 
.A(n_35),
.Y(n_6313)
);

CKINVDCx5p33_ASAP7_75t_R g6314 ( 
.A(n_4676),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_2257),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_1392),
.Y(n_6316)
);

CKINVDCx5p33_ASAP7_75t_R g6317 ( 
.A(n_2523),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_4137),
.Y(n_6318)
);

INVx1_ASAP7_75t_L g6319 ( 
.A(n_4829),
.Y(n_6319)
);

HB1xp67_ASAP7_75t_L g6320 ( 
.A(n_3217),
.Y(n_6320)
);

CKINVDCx5p33_ASAP7_75t_R g6321 ( 
.A(n_3549),
.Y(n_6321)
);

CKINVDCx5p33_ASAP7_75t_R g6322 ( 
.A(n_1505),
.Y(n_6322)
);

CKINVDCx5p33_ASAP7_75t_R g6323 ( 
.A(n_4593),
.Y(n_6323)
);

CKINVDCx5p33_ASAP7_75t_R g6324 ( 
.A(n_4130),
.Y(n_6324)
);

INVx2_ASAP7_75t_L g6325 ( 
.A(n_3126),
.Y(n_6325)
);

CKINVDCx5p33_ASAP7_75t_R g6326 ( 
.A(n_1506),
.Y(n_6326)
);

CKINVDCx5p33_ASAP7_75t_R g6327 ( 
.A(n_1777),
.Y(n_6327)
);

BUFx2_ASAP7_75t_L g6328 ( 
.A(n_4111),
.Y(n_6328)
);

BUFx2_ASAP7_75t_L g6329 ( 
.A(n_2942),
.Y(n_6329)
);

CKINVDCx14_ASAP7_75t_R g6330 ( 
.A(n_3063),
.Y(n_6330)
);

CKINVDCx5p33_ASAP7_75t_R g6331 ( 
.A(n_1979),
.Y(n_6331)
);

CKINVDCx5p33_ASAP7_75t_R g6332 ( 
.A(n_3619),
.Y(n_6332)
);

INVx1_ASAP7_75t_L g6333 ( 
.A(n_254),
.Y(n_6333)
);

INVx4_ASAP7_75t_R g6334 ( 
.A(n_336),
.Y(n_6334)
);

BUFx3_ASAP7_75t_L g6335 ( 
.A(n_4700),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_4772),
.Y(n_6336)
);

INVx1_ASAP7_75t_L g6337 ( 
.A(n_2924),
.Y(n_6337)
);

INVx2_ASAP7_75t_L g6338 ( 
.A(n_4108),
.Y(n_6338)
);

CKINVDCx5p33_ASAP7_75t_R g6339 ( 
.A(n_1768),
.Y(n_6339)
);

CKINVDCx5p33_ASAP7_75t_R g6340 ( 
.A(n_3904),
.Y(n_6340)
);

CKINVDCx20_ASAP7_75t_R g6341 ( 
.A(n_4157),
.Y(n_6341)
);

CKINVDCx5p33_ASAP7_75t_R g6342 ( 
.A(n_2099),
.Y(n_6342)
);

CKINVDCx5p33_ASAP7_75t_R g6343 ( 
.A(n_4250),
.Y(n_6343)
);

BUFx10_ASAP7_75t_L g6344 ( 
.A(n_848),
.Y(n_6344)
);

BUFx3_ASAP7_75t_L g6345 ( 
.A(n_969),
.Y(n_6345)
);

BUFx3_ASAP7_75t_L g6346 ( 
.A(n_437),
.Y(n_6346)
);

HB1xp67_ASAP7_75t_L g6347 ( 
.A(n_2569),
.Y(n_6347)
);

INVx1_ASAP7_75t_L g6348 ( 
.A(n_3660),
.Y(n_6348)
);

CKINVDCx5p33_ASAP7_75t_R g6349 ( 
.A(n_4246),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_1306),
.Y(n_6350)
);

CKINVDCx5p33_ASAP7_75t_R g6351 ( 
.A(n_744),
.Y(n_6351)
);

CKINVDCx5p33_ASAP7_75t_R g6352 ( 
.A(n_741),
.Y(n_6352)
);

BUFx2_ASAP7_75t_L g6353 ( 
.A(n_3488),
.Y(n_6353)
);

INVx1_ASAP7_75t_SL g6354 ( 
.A(n_283),
.Y(n_6354)
);

INVx1_ASAP7_75t_L g6355 ( 
.A(n_1976),
.Y(n_6355)
);

CKINVDCx5p33_ASAP7_75t_R g6356 ( 
.A(n_4496),
.Y(n_6356)
);

INVx1_ASAP7_75t_SL g6357 ( 
.A(n_4121),
.Y(n_6357)
);

CKINVDCx5p33_ASAP7_75t_R g6358 ( 
.A(n_4641),
.Y(n_6358)
);

CKINVDCx5p33_ASAP7_75t_R g6359 ( 
.A(n_2),
.Y(n_6359)
);

INVx1_ASAP7_75t_L g6360 ( 
.A(n_3508),
.Y(n_6360)
);

INVx1_ASAP7_75t_SL g6361 ( 
.A(n_4158),
.Y(n_6361)
);

CKINVDCx16_ASAP7_75t_R g6362 ( 
.A(n_348),
.Y(n_6362)
);

CKINVDCx5p33_ASAP7_75t_R g6363 ( 
.A(n_4208),
.Y(n_6363)
);

INVx1_ASAP7_75t_L g6364 ( 
.A(n_2473),
.Y(n_6364)
);

CKINVDCx20_ASAP7_75t_R g6365 ( 
.A(n_3337),
.Y(n_6365)
);

CKINVDCx5p33_ASAP7_75t_R g6366 ( 
.A(n_2006),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_845),
.Y(n_6367)
);

INVx2_ASAP7_75t_L g6368 ( 
.A(n_3406),
.Y(n_6368)
);

BUFx3_ASAP7_75t_L g6369 ( 
.A(n_4200),
.Y(n_6369)
);

CKINVDCx5p33_ASAP7_75t_R g6370 ( 
.A(n_4097),
.Y(n_6370)
);

INVx1_ASAP7_75t_L g6371 ( 
.A(n_191),
.Y(n_6371)
);

INVx1_ASAP7_75t_L g6372 ( 
.A(n_4268),
.Y(n_6372)
);

INVx1_ASAP7_75t_L g6373 ( 
.A(n_3945),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_1639),
.Y(n_6374)
);

INVx1_ASAP7_75t_SL g6375 ( 
.A(n_4974),
.Y(n_6375)
);

CKINVDCx5p33_ASAP7_75t_R g6376 ( 
.A(n_1479),
.Y(n_6376)
);

CKINVDCx5p33_ASAP7_75t_R g6377 ( 
.A(n_3101),
.Y(n_6377)
);

CKINVDCx5p33_ASAP7_75t_R g6378 ( 
.A(n_482),
.Y(n_6378)
);

CKINVDCx5p33_ASAP7_75t_R g6379 ( 
.A(n_1445),
.Y(n_6379)
);

BUFx3_ASAP7_75t_L g6380 ( 
.A(n_2425),
.Y(n_6380)
);

INVx1_ASAP7_75t_L g6381 ( 
.A(n_1510),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_3839),
.Y(n_6382)
);

BUFx5_ASAP7_75t_L g6383 ( 
.A(n_96),
.Y(n_6383)
);

CKINVDCx20_ASAP7_75t_R g6384 ( 
.A(n_2356),
.Y(n_6384)
);

CKINVDCx5p33_ASAP7_75t_R g6385 ( 
.A(n_4244),
.Y(n_6385)
);

CKINVDCx5p33_ASAP7_75t_R g6386 ( 
.A(n_4409),
.Y(n_6386)
);

CKINVDCx5p33_ASAP7_75t_R g6387 ( 
.A(n_1126),
.Y(n_6387)
);

CKINVDCx5p33_ASAP7_75t_R g6388 ( 
.A(n_3979),
.Y(n_6388)
);

CKINVDCx5p33_ASAP7_75t_R g6389 ( 
.A(n_3672),
.Y(n_6389)
);

INVx1_ASAP7_75t_L g6390 ( 
.A(n_2072),
.Y(n_6390)
);

CKINVDCx5p33_ASAP7_75t_R g6391 ( 
.A(n_1890),
.Y(n_6391)
);

CKINVDCx5p33_ASAP7_75t_R g6392 ( 
.A(n_3317),
.Y(n_6392)
);

CKINVDCx5p33_ASAP7_75t_R g6393 ( 
.A(n_3035),
.Y(n_6393)
);

CKINVDCx5p33_ASAP7_75t_R g6394 ( 
.A(n_689),
.Y(n_6394)
);

CKINVDCx5p33_ASAP7_75t_R g6395 ( 
.A(n_1999),
.Y(n_6395)
);

INVx1_ASAP7_75t_SL g6396 ( 
.A(n_4305),
.Y(n_6396)
);

CKINVDCx5p33_ASAP7_75t_R g6397 ( 
.A(n_4120),
.Y(n_6397)
);

CKINVDCx5p33_ASAP7_75t_R g6398 ( 
.A(n_2191),
.Y(n_6398)
);

CKINVDCx16_ASAP7_75t_R g6399 ( 
.A(n_3967),
.Y(n_6399)
);

CKINVDCx20_ASAP7_75t_R g6400 ( 
.A(n_3560),
.Y(n_6400)
);

CKINVDCx5p33_ASAP7_75t_R g6401 ( 
.A(n_800),
.Y(n_6401)
);

CKINVDCx5p33_ASAP7_75t_R g6402 ( 
.A(n_1173),
.Y(n_6402)
);

CKINVDCx20_ASAP7_75t_R g6403 ( 
.A(n_4198),
.Y(n_6403)
);

CKINVDCx5p33_ASAP7_75t_R g6404 ( 
.A(n_3566),
.Y(n_6404)
);

INVx1_ASAP7_75t_L g6405 ( 
.A(n_538),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_4240),
.Y(n_6406)
);

INVx2_ASAP7_75t_L g6407 ( 
.A(n_3367),
.Y(n_6407)
);

CKINVDCx20_ASAP7_75t_R g6408 ( 
.A(n_3771),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_2517),
.Y(n_6409)
);

BUFx3_ASAP7_75t_L g6410 ( 
.A(n_1043),
.Y(n_6410)
);

CKINVDCx5p33_ASAP7_75t_R g6411 ( 
.A(n_2934),
.Y(n_6411)
);

CKINVDCx5p33_ASAP7_75t_R g6412 ( 
.A(n_3807),
.Y(n_6412)
);

INVx1_ASAP7_75t_SL g6413 ( 
.A(n_2259),
.Y(n_6413)
);

CKINVDCx5p33_ASAP7_75t_R g6414 ( 
.A(n_4399),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_4146),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_3435),
.Y(n_6416)
);

CKINVDCx20_ASAP7_75t_R g6417 ( 
.A(n_734),
.Y(n_6417)
);

CKINVDCx5p33_ASAP7_75t_R g6418 ( 
.A(n_1122),
.Y(n_6418)
);

INVxp33_ASAP7_75t_SL g6419 ( 
.A(n_3316),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_1342),
.Y(n_6420)
);

CKINVDCx20_ASAP7_75t_R g6421 ( 
.A(n_4258),
.Y(n_6421)
);

INVx2_ASAP7_75t_SL g6422 ( 
.A(n_91),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_1927),
.Y(n_6423)
);

CKINVDCx5p33_ASAP7_75t_R g6424 ( 
.A(n_3227),
.Y(n_6424)
);

CKINVDCx5p33_ASAP7_75t_R g6425 ( 
.A(n_1088),
.Y(n_6425)
);

CKINVDCx5p33_ASAP7_75t_R g6426 ( 
.A(n_3749),
.Y(n_6426)
);

BUFx3_ASAP7_75t_L g6427 ( 
.A(n_4280),
.Y(n_6427)
);

CKINVDCx5p33_ASAP7_75t_R g6428 ( 
.A(n_4150),
.Y(n_6428)
);

INVx1_ASAP7_75t_L g6429 ( 
.A(n_2423),
.Y(n_6429)
);

CKINVDCx16_ASAP7_75t_R g6430 ( 
.A(n_2495),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_4026),
.Y(n_6431)
);

CKINVDCx5p33_ASAP7_75t_R g6432 ( 
.A(n_4196),
.Y(n_6432)
);

INVx1_ASAP7_75t_L g6433 ( 
.A(n_703),
.Y(n_6433)
);

CKINVDCx20_ASAP7_75t_R g6434 ( 
.A(n_4147),
.Y(n_6434)
);

CKINVDCx5p33_ASAP7_75t_R g6435 ( 
.A(n_3420),
.Y(n_6435)
);

CKINVDCx5p33_ASAP7_75t_R g6436 ( 
.A(n_4495),
.Y(n_6436)
);

CKINVDCx5p33_ASAP7_75t_R g6437 ( 
.A(n_3043),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_2628),
.Y(n_6438)
);

CKINVDCx5p33_ASAP7_75t_R g6439 ( 
.A(n_73),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_235),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_3141),
.Y(n_6441)
);

INVx1_ASAP7_75t_L g6442 ( 
.A(n_2976),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_4178),
.Y(n_6443)
);

CKINVDCx5p33_ASAP7_75t_R g6444 ( 
.A(n_4352),
.Y(n_6444)
);

CKINVDCx5p33_ASAP7_75t_R g6445 ( 
.A(n_296),
.Y(n_6445)
);

CKINVDCx5p33_ASAP7_75t_R g6446 ( 
.A(n_2591),
.Y(n_6446)
);

INVx1_ASAP7_75t_L g6447 ( 
.A(n_4146),
.Y(n_6447)
);

CKINVDCx5p33_ASAP7_75t_R g6448 ( 
.A(n_3590),
.Y(n_6448)
);

INVx2_ASAP7_75t_SL g6449 ( 
.A(n_4230),
.Y(n_6449)
);

CKINVDCx5p33_ASAP7_75t_R g6450 ( 
.A(n_4180),
.Y(n_6450)
);

CKINVDCx5p33_ASAP7_75t_R g6451 ( 
.A(n_3975),
.Y(n_6451)
);

CKINVDCx5p33_ASAP7_75t_R g6452 ( 
.A(n_4022),
.Y(n_6452)
);

CKINVDCx5p33_ASAP7_75t_R g6453 ( 
.A(n_3368),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_375),
.Y(n_6454)
);

INVx1_ASAP7_75t_L g6455 ( 
.A(n_4162),
.Y(n_6455)
);

BUFx10_ASAP7_75t_L g6456 ( 
.A(n_790),
.Y(n_6456)
);

INVx1_ASAP7_75t_L g6457 ( 
.A(n_4101),
.Y(n_6457)
);

CKINVDCx5p33_ASAP7_75t_R g6458 ( 
.A(n_2160),
.Y(n_6458)
);

CKINVDCx20_ASAP7_75t_R g6459 ( 
.A(n_4262),
.Y(n_6459)
);

INVx2_ASAP7_75t_SL g6460 ( 
.A(n_139),
.Y(n_6460)
);

CKINVDCx5p33_ASAP7_75t_R g6461 ( 
.A(n_4204),
.Y(n_6461)
);

INVx1_ASAP7_75t_L g6462 ( 
.A(n_1467),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_2650),
.Y(n_6463)
);

CKINVDCx5p33_ASAP7_75t_R g6464 ( 
.A(n_1375),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_4233),
.Y(n_6465)
);

BUFx3_ASAP7_75t_L g6466 ( 
.A(n_3698),
.Y(n_6466)
);

CKINVDCx16_ASAP7_75t_R g6467 ( 
.A(n_614),
.Y(n_6467)
);

INVxp67_ASAP7_75t_L g6468 ( 
.A(n_1520),
.Y(n_6468)
);

BUFx2_ASAP7_75t_L g6469 ( 
.A(n_3409),
.Y(n_6469)
);

CKINVDCx20_ASAP7_75t_R g6470 ( 
.A(n_3094),
.Y(n_6470)
);

CKINVDCx5p33_ASAP7_75t_R g6471 ( 
.A(n_4302),
.Y(n_6471)
);

INVx1_ASAP7_75t_L g6472 ( 
.A(n_1961),
.Y(n_6472)
);

CKINVDCx5p33_ASAP7_75t_R g6473 ( 
.A(n_2652),
.Y(n_6473)
);

INVx1_ASAP7_75t_L g6474 ( 
.A(n_2687),
.Y(n_6474)
);

CKINVDCx5p33_ASAP7_75t_R g6475 ( 
.A(n_4322),
.Y(n_6475)
);

CKINVDCx5p33_ASAP7_75t_R g6476 ( 
.A(n_3093),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_2793),
.Y(n_6477)
);

BUFx3_ASAP7_75t_L g6478 ( 
.A(n_3215),
.Y(n_6478)
);

CKINVDCx5p33_ASAP7_75t_R g6479 ( 
.A(n_343),
.Y(n_6479)
);

CKINVDCx5p33_ASAP7_75t_R g6480 ( 
.A(n_252),
.Y(n_6480)
);

CKINVDCx5p33_ASAP7_75t_R g6481 ( 
.A(n_3971),
.Y(n_6481)
);

INVx2_ASAP7_75t_L g6482 ( 
.A(n_4282),
.Y(n_6482)
);

CKINVDCx5p33_ASAP7_75t_R g6483 ( 
.A(n_1979),
.Y(n_6483)
);

INVx1_ASAP7_75t_L g6484 ( 
.A(n_4245),
.Y(n_6484)
);

INVx1_ASAP7_75t_SL g6485 ( 
.A(n_4049),
.Y(n_6485)
);

BUFx6f_ASAP7_75t_L g6486 ( 
.A(n_3382),
.Y(n_6486)
);

BUFx8_ASAP7_75t_SL g6487 ( 
.A(n_3097),
.Y(n_6487)
);

CKINVDCx5p33_ASAP7_75t_R g6488 ( 
.A(n_1743),
.Y(n_6488)
);

CKINVDCx5p33_ASAP7_75t_R g6489 ( 
.A(n_4182),
.Y(n_6489)
);

INVx2_ASAP7_75t_L g6490 ( 
.A(n_5175),
.Y(n_6490)
);

CKINVDCx5p33_ASAP7_75t_R g6491 ( 
.A(n_5333),
.Y(n_6491)
);

INVx2_ASAP7_75t_L g6492 ( 
.A(n_5175),
.Y(n_6492)
);

INVx1_ASAP7_75t_L g6493 ( 
.A(n_5175),
.Y(n_6493)
);

CKINVDCx5p33_ASAP7_75t_R g6494 ( 
.A(n_5596),
.Y(n_6494)
);

NOR2xp33_ASAP7_75t_L g6495 ( 
.A(n_6243),
.B(n_5136),
.Y(n_6495)
);

BUFx3_ASAP7_75t_L g6496 ( 
.A(n_5312),
.Y(n_6496)
);

INVxp67_ASAP7_75t_L g6497 ( 
.A(n_5041),
.Y(n_6497)
);

BUFx3_ASAP7_75t_L g6498 ( 
.A(n_5312),
.Y(n_6498)
);

CKINVDCx5p33_ASAP7_75t_R g6499 ( 
.A(n_6024),
.Y(n_6499)
);

CKINVDCx5p33_ASAP7_75t_R g6500 ( 
.A(n_6161),
.Y(n_6500)
);

CKINVDCx5p33_ASAP7_75t_R g6501 ( 
.A(n_6487),
.Y(n_6501)
);

INVx1_ASAP7_75t_L g6502 ( 
.A(n_5175),
.Y(n_6502)
);

INVx1_ASAP7_75t_L g6503 ( 
.A(n_5175),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_5457),
.Y(n_6504)
);

INVxp67_ASAP7_75t_SL g6505 ( 
.A(n_6020),
.Y(n_6505)
);

CKINVDCx5p33_ASAP7_75t_R g6506 ( 
.A(n_5044),
.Y(n_6506)
);

INVx1_ASAP7_75t_L g6507 ( 
.A(n_5457),
.Y(n_6507)
);

BUFx2_ASAP7_75t_L g6508 ( 
.A(n_5043),
.Y(n_6508)
);

INVxp67_ASAP7_75t_L g6509 ( 
.A(n_5087),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_5457),
.Y(n_6510)
);

CKINVDCx20_ASAP7_75t_R g6511 ( 
.A(n_5688),
.Y(n_6511)
);

BUFx3_ASAP7_75t_L g6512 ( 
.A(n_5133),
.Y(n_6512)
);

INVx2_ASAP7_75t_L g6513 ( 
.A(n_5457),
.Y(n_6513)
);

CKINVDCx5p33_ASAP7_75t_R g6514 ( 
.A(n_5051),
.Y(n_6514)
);

CKINVDCx5p33_ASAP7_75t_R g6515 ( 
.A(n_5058),
.Y(n_6515)
);

INVx1_ASAP7_75t_L g6516 ( 
.A(n_5457),
.Y(n_6516)
);

CKINVDCx5p33_ASAP7_75t_R g6517 ( 
.A(n_5065),
.Y(n_6517)
);

INVx1_ASAP7_75t_L g6518 ( 
.A(n_5698),
.Y(n_6518)
);

CKINVDCx5p33_ASAP7_75t_R g6519 ( 
.A(n_5077),
.Y(n_6519)
);

INVx2_ASAP7_75t_SL g6520 ( 
.A(n_5073),
.Y(n_6520)
);

CKINVDCx5p33_ASAP7_75t_R g6521 ( 
.A(n_5101),
.Y(n_6521)
);

INVx1_ASAP7_75t_L g6522 ( 
.A(n_5698),
.Y(n_6522)
);

INVx1_ASAP7_75t_L g6523 ( 
.A(n_5698),
.Y(n_6523)
);

BUFx2_ASAP7_75t_SL g6524 ( 
.A(n_5771),
.Y(n_6524)
);

HB1xp67_ASAP7_75t_L g6525 ( 
.A(n_5151),
.Y(n_6525)
);

BUFx6f_ASAP7_75t_L g6526 ( 
.A(n_5057),
.Y(n_6526)
);

INVx2_ASAP7_75t_SL g6527 ( 
.A(n_5073),
.Y(n_6527)
);

CKINVDCx5p33_ASAP7_75t_R g6528 ( 
.A(n_5104),
.Y(n_6528)
);

INVx2_ASAP7_75t_L g6529 ( 
.A(n_5698),
.Y(n_6529)
);

INVx1_ASAP7_75t_L g6530 ( 
.A(n_5698),
.Y(n_6530)
);

INVx1_ASAP7_75t_L g6531 ( 
.A(n_6075),
.Y(n_6531)
);

INVx1_ASAP7_75t_L g6532 ( 
.A(n_6075),
.Y(n_6532)
);

CKINVDCx5p33_ASAP7_75t_R g6533 ( 
.A(n_5156),
.Y(n_6533)
);

CKINVDCx5p33_ASAP7_75t_R g6534 ( 
.A(n_5167),
.Y(n_6534)
);

CKINVDCx5p33_ASAP7_75t_R g6535 ( 
.A(n_5189),
.Y(n_6535)
);

INVx1_ASAP7_75t_L g6536 ( 
.A(n_6075),
.Y(n_6536)
);

CKINVDCx20_ASAP7_75t_R g6537 ( 
.A(n_5931),
.Y(n_6537)
);

CKINVDCx5p33_ASAP7_75t_R g6538 ( 
.A(n_5240),
.Y(n_6538)
);

INVx1_ASAP7_75t_L g6539 ( 
.A(n_6075),
.Y(n_6539)
);

INVx1_ASAP7_75t_L g6540 ( 
.A(n_6075),
.Y(n_6540)
);

BUFx3_ASAP7_75t_L g6541 ( 
.A(n_5374),
.Y(n_6541)
);

INVxp67_ASAP7_75t_L g6542 ( 
.A(n_5134),
.Y(n_6542)
);

INVx2_ASAP7_75t_L g6543 ( 
.A(n_6153),
.Y(n_6543)
);

CKINVDCx5p33_ASAP7_75t_R g6544 ( 
.A(n_5315),
.Y(n_6544)
);

CKINVDCx5p33_ASAP7_75t_R g6545 ( 
.A(n_5334),
.Y(n_6545)
);

CKINVDCx20_ASAP7_75t_R g6546 ( 
.A(n_5973),
.Y(n_6546)
);

CKINVDCx5p33_ASAP7_75t_R g6547 ( 
.A(n_5364),
.Y(n_6547)
);

INVx1_ASAP7_75t_L g6548 ( 
.A(n_6153),
.Y(n_6548)
);

INVx2_ASAP7_75t_L g6549 ( 
.A(n_6153),
.Y(n_6549)
);

CKINVDCx5p33_ASAP7_75t_R g6550 ( 
.A(n_5430),
.Y(n_6550)
);

INVx1_ASAP7_75t_L g6551 ( 
.A(n_6153),
.Y(n_6551)
);

CKINVDCx5p33_ASAP7_75t_R g6552 ( 
.A(n_5458),
.Y(n_6552)
);

BUFx2_ASAP7_75t_L g6553 ( 
.A(n_5194),
.Y(n_6553)
);

BUFx6f_ASAP7_75t_L g6554 ( 
.A(n_5057),
.Y(n_6554)
);

INVx2_ASAP7_75t_L g6555 ( 
.A(n_6153),
.Y(n_6555)
);

CKINVDCx5p33_ASAP7_75t_R g6556 ( 
.A(n_5463),
.Y(n_6556)
);

INVx1_ASAP7_75t_L g6557 ( 
.A(n_6169),
.Y(n_6557)
);

INVx2_ASAP7_75t_SL g6558 ( 
.A(n_5210),
.Y(n_6558)
);

INVx1_ASAP7_75t_L g6559 ( 
.A(n_6169),
.Y(n_6559)
);

INVx1_ASAP7_75t_L g6560 ( 
.A(n_6169),
.Y(n_6560)
);

INVx1_ASAP7_75t_L g6561 ( 
.A(n_6169),
.Y(n_6561)
);

CKINVDCx5p33_ASAP7_75t_R g6562 ( 
.A(n_5474),
.Y(n_6562)
);

CKINVDCx5p33_ASAP7_75t_R g6563 ( 
.A(n_5477),
.Y(n_6563)
);

CKINVDCx5p33_ASAP7_75t_R g6564 ( 
.A(n_5488),
.Y(n_6564)
);

BUFx6f_ASAP7_75t_L g6565 ( 
.A(n_5057),
.Y(n_6565)
);

INVx2_ASAP7_75t_L g6566 ( 
.A(n_6169),
.Y(n_6566)
);

INVx1_ASAP7_75t_L g6567 ( 
.A(n_6209),
.Y(n_6567)
);

CKINVDCx5p33_ASAP7_75t_R g6568 ( 
.A(n_5503),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_6209),
.Y(n_6569)
);

INVx1_ASAP7_75t_L g6570 ( 
.A(n_6209),
.Y(n_6570)
);

INVx1_ASAP7_75t_L g6571 ( 
.A(n_6209),
.Y(n_6571)
);

INVx1_ASAP7_75t_L g6572 ( 
.A(n_6209),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_6383),
.Y(n_6573)
);

CKINVDCx5p33_ASAP7_75t_R g6574 ( 
.A(n_5506),
.Y(n_6574)
);

INVx1_ASAP7_75t_L g6575 ( 
.A(n_6383),
.Y(n_6575)
);

CKINVDCx5p33_ASAP7_75t_R g6576 ( 
.A(n_5547),
.Y(n_6576)
);

CKINVDCx5p33_ASAP7_75t_R g6577 ( 
.A(n_5555),
.Y(n_6577)
);

CKINVDCx5p33_ASAP7_75t_R g6578 ( 
.A(n_5590),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_6383),
.Y(n_6579)
);

CKINVDCx5p33_ASAP7_75t_R g6580 ( 
.A(n_5604),
.Y(n_6580)
);

HB1xp67_ASAP7_75t_L g6581 ( 
.A(n_5264),
.Y(n_6581)
);

INVx2_ASAP7_75t_SL g6582 ( 
.A(n_5210),
.Y(n_6582)
);

CKINVDCx5p33_ASAP7_75t_R g6583 ( 
.A(n_5605),
.Y(n_6583)
);

CKINVDCx5p33_ASAP7_75t_R g6584 ( 
.A(n_5622),
.Y(n_6584)
);

BUFx2_ASAP7_75t_L g6585 ( 
.A(n_5269),
.Y(n_6585)
);

INVx2_ASAP7_75t_L g6586 ( 
.A(n_6383),
.Y(n_6586)
);

CKINVDCx5p33_ASAP7_75t_R g6587 ( 
.A(n_5656),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_6383),
.Y(n_6588)
);

INVx2_ASAP7_75t_L g6589 ( 
.A(n_6486),
.Y(n_6589)
);

CKINVDCx5p33_ASAP7_75t_R g6590 ( 
.A(n_5665),
.Y(n_6590)
);

CKINVDCx5p33_ASAP7_75t_R g6591 ( 
.A(n_5668),
.Y(n_6591)
);

BUFx5_ASAP7_75t_L g6592 ( 
.A(n_5055),
.Y(n_6592)
);

CKINVDCx5p33_ASAP7_75t_R g6593 ( 
.A(n_5679),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_5176),
.Y(n_6594)
);

CKINVDCx5p33_ASAP7_75t_R g6595 ( 
.A(n_5681),
.Y(n_6595)
);

INVx2_ASAP7_75t_L g6596 ( 
.A(n_6486),
.Y(n_6596)
);

CKINVDCx16_ASAP7_75t_R g6597 ( 
.A(n_5302),
.Y(n_6597)
);

CKINVDCx5p33_ASAP7_75t_R g6598 ( 
.A(n_5693),
.Y(n_6598)
);

INVx1_ASAP7_75t_L g6599 ( 
.A(n_5176),
.Y(n_6599)
);

CKINVDCx20_ASAP7_75t_R g6600 ( 
.A(n_6156),
.Y(n_6600)
);

NOR2xp67_ASAP7_75t_L g6601 ( 
.A(n_5308),
.B(n_0),
.Y(n_6601)
);

INVx2_ASAP7_75t_L g6602 ( 
.A(n_6486),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_5308),
.Y(n_6603)
);

CKINVDCx20_ASAP7_75t_R g6604 ( 
.A(n_6151),
.Y(n_6604)
);

BUFx8_ASAP7_75t_SL g6605 ( 
.A(n_5287),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_5170),
.Y(n_6606)
);

BUFx2_ASAP7_75t_L g6607 ( 
.A(n_5330),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_5170),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_5170),
.Y(n_6609)
);

CKINVDCx5p33_ASAP7_75t_R g6610 ( 
.A(n_5701),
.Y(n_6610)
);

CKINVDCx5p33_ASAP7_75t_R g6611 ( 
.A(n_5711),
.Y(n_6611)
);

INVx1_ASAP7_75t_L g6612 ( 
.A(n_5177),
.Y(n_6612)
);

INVx1_ASAP7_75t_L g6613 ( 
.A(n_5177),
.Y(n_6613)
);

BUFx10_ASAP7_75t_L g6614 ( 
.A(n_5099),
.Y(n_6614)
);

CKINVDCx5p33_ASAP7_75t_R g6615 ( 
.A(n_5714),
.Y(n_6615)
);

HB1xp67_ASAP7_75t_L g6616 ( 
.A(n_5318),
.Y(n_6616)
);

CKINVDCx5p33_ASAP7_75t_R g6617 ( 
.A(n_5738),
.Y(n_6617)
);

CKINVDCx5p33_ASAP7_75t_R g6618 ( 
.A(n_5743),
.Y(n_6618)
);

CKINVDCx5p33_ASAP7_75t_R g6619 ( 
.A(n_5764),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_5177),
.Y(n_6620)
);

CKINVDCx5p33_ASAP7_75t_R g6621 ( 
.A(n_5768),
.Y(n_6621)
);

BUFx3_ASAP7_75t_L g6622 ( 
.A(n_5707),
.Y(n_6622)
);

CKINVDCx5p33_ASAP7_75t_R g6623 ( 
.A(n_5854),
.Y(n_6623)
);

INVx1_ASAP7_75t_L g6624 ( 
.A(n_5221),
.Y(n_6624)
);

CKINVDCx5p33_ASAP7_75t_R g6625 ( 
.A(n_5865),
.Y(n_6625)
);

CKINVDCx20_ASAP7_75t_R g6626 ( 
.A(n_5080),
.Y(n_6626)
);

NOR2xp67_ASAP7_75t_L g6627 ( 
.A(n_5256),
.B(n_0),
.Y(n_6627)
);

INVx2_ASAP7_75t_L g6628 ( 
.A(n_5221),
.Y(n_6628)
);

CKINVDCx5p33_ASAP7_75t_R g6629 ( 
.A(n_5877),
.Y(n_6629)
);

INVx1_ASAP7_75t_L g6630 ( 
.A(n_5221),
.Y(n_6630)
);

CKINVDCx20_ASAP7_75t_R g6631 ( 
.A(n_5184),
.Y(n_6631)
);

INVx1_ASAP7_75t_L g6632 ( 
.A(n_5224),
.Y(n_6632)
);

BUFx2_ASAP7_75t_L g6633 ( 
.A(n_5342),
.Y(n_6633)
);

NOR2xp67_ASAP7_75t_L g6634 ( 
.A(n_5376),
.B(n_1),
.Y(n_6634)
);

BUFx3_ASAP7_75t_L g6635 ( 
.A(n_6295),
.Y(n_6635)
);

CKINVDCx5p33_ASAP7_75t_R g6636 ( 
.A(n_5919),
.Y(n_6636)
);

NOR2xp67_ASAP7_75t_L g6637 ( 
.A(n_5539),
.B(n_1),
.Y(n_6637)
);

INVx1_ASAP7_75t_L g6638 ( 
.A(n_5224),
.Y(n_6638)
);

INVx1_ASAP7_75t_L g6639 ( 
.A(n_5224),
.Y(n_6639)
);

CKINVDCx20_ASAP7_75t_R g6640 ( 
.A(n_5252),
.Y(n_6640)
);

CKINVDCx5p33_ASAP7_75t_R g6641 ( 
.A(n_5928),
.Y(n_6641)
);

CKINVDCx5p33_ASAP7_75t_R g6642 ( 
.A(n_5937),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_5676),
.Y(n_6643)
);

CKINVDCx5p33_ASAP7_75t_R g6644 ( 
.A(n_5950),
.Y(n_6644)
);

INVx1_ASAP7_75t_L g6645 ( 
.A(n_5676),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_5676),
.Y(n_6646)
);

CKINVDCx5p33_ASAP7_75t_R g6647 ( 
.A(n_5953),
.Y(n_6647)
);

CKINVDCx5p33_ASAP7_75t_R g6648 ( 
.A(n_5954),
.Y(n_6648)
);

CKINVDCx5p33_ASAP7_75t_R g6649 ( 
.A(n_5977),
.Y(n_6649)
);

CKINVDCx5p33_ASAP7_75t_R g6650 ( 
.A(n_5978),
.Y(n_6650)
);

BUFx6f_ASAP7_75t_L g6651 ( 
.A(n_5690),
.Y(n_6651)
);

CKINVDCx20_ASAP7_75t_R g6652 ( 
.A(n_5762),
.Y(n_6652)
);

INVx1_ASAP7_75t_L g6653 ( 
.A(n_5690),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_5690),
.Y(n_6654)
);

HB1xp67_ASAP7_75t_L g6655 ( 
.A(n_5356),
.Y(n_6655)
);

INVx1_ASAP7_75t_L g6656 ( 
.A(n_5821),
.Y(n_6656)
);

BUFx3_ASAP7_75t_L g6657 ( 
.A(n_6335),
.Y(n_6657)
);

CKINVDCx5p33_ASAP7_75t_R g6658 ( 
.A(n_6000),
.Y(n_6658)
);

INVx2_ASAP7_75t_L g6659 ( 
.A(n_5821),
.Y(n_6659)
);

CKINVDCx5p33_ASAP7_75t_R g6660 ( 
.A(n_6006),
.Y(n_6660)
);

HB1xp67_ASAP7_75t_L g6661 ( 
.A(n_5434),
.Y(n_6661)
);

CKINVDCx5p33_ASAP7_75t_R g6662 ( 
.A(n_6011),
.Y(n_6662)
);

INVx2_ASAP7_75t_L g6663 ( 
.A(n_5821),
.Y(n_6663)
);

INVx2_ASAP7_75t_SL g6664 ( 
.A(n_5216),
.Y(n_6664)
);

BUFx5_ASAP7_75t_L g6665 ( 
.A(n_5067),
.Y(n_6665)
);

CKINVDCx5p33_ASAP7_75t_R g6666 ( 
.A(n_6019),
.Y(n_6666)
);

CKINVDCx5p33_ASAP7_75t_R g6667 ( 
.A(n_6032),
.Y(n_6667)
);

INVxp33_ASAP7_75t_SL g6668 ( 
.A(n_5214),
.Y(n_6668)
);

CKINVDCx5p33_ASAP7_75t_R g6669 ( 
.A(n_6054),
.Y(n_6669)
);

CKINVDCx5p33_ASAP7_75t_R g6670 ( 
.A(n_6086),
.Y(n_6670)
);

BUFx3_ASAP7_75t_L g6671 ( 
.A(n_5054),
.Y(n_6671)
);

INVx1_ASAP7_75t_SL g6672 ( 
.A(n_5476),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_5906),
.Y(n_6673)
);

CKINVDCx5p33_ASAP7_75t_R g6674 ( 
.A(n_6127),
.Y(n_6674)
);

INVx1_ASAP7_75t_SL g6675 ( 
.A(n_5640),
.Y(n_6675)
);

INVx1_ASAP7_75t_L g6676 ( 
.A(n_5906),
.Y(n_6676)
);

INVx1_ASAP7_75t_L g6677 ( 
.A(n_5906),
.Y(n_6677)
);

CKINVDCx5p33_ASAP7_75t_R g6678 ( 
.A(n_6202),
.Y(n_6678)
);

CKINVDCx5p33_ASAP7_75t_R g6679 ( 
.A(n_6220),
.Y(n_6679)
);

CKINVDCx5p33_ASAP7_75t_R g6680 ( 
.A(n_6230),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_5951),
.Y(n_6681)
);

CKINVDCx5p33_ASAP7_75t_R g6682 ( 
.A(n_6263),
.Y(n_6682)
);

INVx1_ASAP7_75t_L g6683 ( 
.A(n_5951),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_5951),
.Y(n_6684)
);

CKINVDCx5p33_ASAP7_75t_R g6685 ( 
.A(n_6308),
.Y(n_6685)
);

INVxp67_ASAP7_75t_SL g6686 ( 
.A(n_5814),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_6002),
.Y(n_6687)
);

INVx1_ASAP7_75t_SL g6688 ( 
.A(n_5773),
.Y(n_6688)
);

INVx1_ASAP7_75t_L g6689 ( 
.A(n_6002),
.Y(n_6689)
);

CKINVDCx5p33_ASAP7_75t_R g6690 ( 
.A(n_6314),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6002),
.Y(n_6691)
);

INVx1_ASAP7_75t_SL g6692 ( 
.A(n_5820),
.Y(n_6692)
);

INVx1_ASAP7_75t_L g6693 ( 
.A(n_6091),
.Y(n_6693)
);

CKINVDCx20_ASAP7_75t_R g6694 ( 
.A(n_5789),
.Y(n_6694)
);

INVx1_ASAP7_75t_L g6695 ( 
.A(n_6091),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_6091),
.Y(n_6696)
);

CKINVDCx5p33_ASAP7_75t_R g6697 ( 
.A(n_6323),
.Y(n_6697)
);

CKINVDCx5p33_ASAP7_75t_R g6698 ( 
.A(n_6356),
.Y(n_6698)
);

INVx1_ASAP7_75t_L g6699 ( 
.A(n_6280),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_6280),
.Y(n_6700)
);

INVxp67_ASAP7_75t_SL g6701 ( 
.A(n_5382),
.Y(n_6701)
);

INVx2_ASAP7_75t_L g6702 ( 
.A(n_6280),
.Y(n_6702)
);

CKINVDCx5p33_ASAP7_75t_R g6703 ( 
.A(n_6358),
.Y(n_6703)
);

INVx1_ASAP7_75t_L g6704 ( 
.A(n_6282),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_6282),
.Y(n_6705)
);

INVx2_ASAP7_75t_L g6706 ( 
.A(n_6282),
.Y(n_6706)
);

CKINVDCx5p33_ASAP7_75t_R g6707 ( 
.A(n_6386),
.Y(n_6707)
);

CKINVDCx5p33_ASAP7_75t_R g6708 ( 
.A(n_6414),
.Y(n_6708)
);

NAND2xp5_ASAP7_75t_L g6709 ( 
.A(n_5830),
.B(n_6021),
.Y(n_6709)
);

INVx1_ASAP7_75t_L g6710 ( 
.A(n_5089),
.Y(n_6710)
);

CKINVDCx5p33_ASAP7_75t_R g6711 ( 
.A(n_6436),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_5105),
.Y(n_6712)
);

INVx1_ASAP7_75t_L g6713 ( 
.A(n_5150),
.Y(n_6713)
);

INVx1_ASAP7_75t_L g6714 ( 
.A(n_5206),
.Y(n_6714)
);

CKINVDCx5p33_ASAP7_75t_R g6715 ( 
.A(n_6444),
.Y(n_6715)
);

CKINVDCx5p33_ASAP7_75t_R g6716 ( 
.A(n_6330),
.Y(n_6716)
);

CKINVDCx5p33_ASAP7_75t_R g6717 ( 
.A(n_5523),
.Y(n_6717)
);

INVx1_ASAP7_75t_L g6718 ( 
.A(n_5286),
.Y(n_6718)
);

CKINVDCx5p33_ASAP7_75t_R g6719 ( 
.A(n_5741),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_5327),
.Y(n_6720)
);

CKINVDCx20_ASAP7_75t_R g6721 ( 
.A(n_6082),
.Y(n_6721)
);

INVx1_ASAP7_75t_SL g6722 ( 
.A(n_5995),
.Y(n_6722)
);

BUFx3_ASAP7_75t_L g6723 ( 
.A(n_5328),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_5409),
.Y(n_6724)
);

CKINVDCx5p33_ASAP7_75t_R g6725 ( 
.A(n_6193),
.Y(n_6725)
);

CKINVDCx5p33_ASAP7_75t_R g6726 ( 
.A(n_6195),
.Y(n_6726)
);

CKINVDCx5p33_ASAP7_75t_R g6727 ( 
.A(n_6250),
.Y(n_6727)
);

INVxp33_ASAP7_75t_L g6728 ( 
.A(n_5467),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_5426),
.Y(n_6729)
);

INVx1_ASAP7_75t_L g6730 ( 
.A(n_5536),
.Y(n_6730)
);

CKINVDCx5p33_ASAP7_75t_R g6731 ( 
.A(n_6264),
.Y(n_6731)
);

CKINVDCx5p33_ASAP7_75t_R g6732 ( 
.A(n_6313),
.Y(n_6732)
);

BUFx6f_ASAP7_75t_L g6733 ( 
.A(n_5621),
.Y(n_6733)
);

INVx1_ASAP7_75t_L g6734 ( 
.A(n_5816),
.Y(n_6734)
);

CKINVDCx5p33_ASAP7_75t_R g6735 ( 
.A(n_6362),
.Y(n_6735)
);

CKINVDCx5p33_ASAP7_75t_R g6736 ( 
.A(n_6399),
.Y(n_6736)
);

INVx1_ASAP7_75t_L g6737 ( 
.A(n_5829),
.Y(n_6737)
);

INVxp67_ASAP7_75t_L g6738 ( 
.A(n_5998),
.Y(n_6738)
);

BUFx3_ASAP7_75t_L g6739 ( 
.A(n_5849),
.Y(n_6739)
);

CKINVDCx5p33_ASAP7_75t_R g6740 ( 
.A(n_6430),
.Y(n_6740)
);

INVx1_ASAP7_75t_L g6741 ( 
.A(n_5939),
.Y(n_6741)
);

INVx1_ASAP7_75t_L g6742 ( 
.A(n_5974),
.Y(n_6742)
);

HB1xp67_ASAP7_75t_L g6743 ( 
.A(n_6467),
.Y(n_6743)
);

INVx1_ASAP7_75t_L g6744 ( 
.A(n_5975),
.Y(n_6744)
);

INVx1_ASAP7_75t_L g6745 ( 
.A(n_6042),
.Y(n_6745)
);

INVx1_ASAP7_75t_L g6746 ( 
.A(n_6085),
.Y(n_6746)
);

CKINVDCx5p33_ASAP7_75t_R g6747 ( 
.A(n_6476),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_5273),
.Y(n_6748)
);

CKINVDCx5p33_ASAP7_75t_R g6749 ( 
.A(n_6479),
.Y(n_6749)
);

CKINVDCx5p33_ASAP7_75t_R g6750 ( 
.A(n_6480),
.Y(n_6750)
);

INVx1_ASAP7_75t_L g6751 ( 
.A(n_6100),
.Y(n_6751)
);

CKINVDCx20_ASAP7_75t_R g6752 ( 
.A(n_5140),
.Y(n_6752)
);

INVx1_ASAP7_75t_L g6753 ( 
.A(n_6218),
.Y(n_6753)
);

INVx1_ASAP7_75t_L g6754 ( 
.A(n_6234),
.Y(n_6754)
);

INVx1_ASAP7_75t_L g6755 ( 
.A(n_6261),
.Y(n_6755)
);

INVx1_ASAP7_75t_L g6756 ( 
.A(n_6345),
.Y(n_6756)
);

CKINVDCx5p33_ASAP7_75t_R g6757 ( 
.A(n_6488),
.Y(n_6757)
);

CKINVDCx5p33_ASAP7_75t_R g6758 ( 
.A(n_6489),
.Y(n_6758)
);

CKINVDCx5p33_ASAP7_75t_R g6759 ( 
.A(n_5039),
.Y(n_6759)
);

CKINVDCx5p33_ASAP7_75t_R g6760 ( 
.A(n_5040),
.Y(n_6760)
);

CKINVDCx5p33_ASAP7_75t_R g6761 ( 
.A(n_6471),
.Y(n_6761)
);

CKINVDCx5p33_ASAP7_75t_R g6762 ( 
.A(n_6473),
.Y(n_6762)
);

INVx1_ASAP7_75t_L g6763 ( 
.A(n_6346),
.Y(n_6763)
);

INVx1_ASAP7_75t_L g6764 ( 
.A(n_6369),
.Y(n_6764)
);

BUFx2_ASAP7_75t_L g6765 ( 
.A(n_6072),
.Y(n_6765)
);

CKINVDCx5p33_ASAP7_75t_R g6766 ( 
.A(n_6475),
.Y(n_6766)
);

INVx1_ASAP7_75t_L g6767 ( 
.A(n_6380),
.Y(n_6767)
);

CKINVDCx16_ASAP7_75t_R g6768 ( 
.A(n_5216),
.Y(n_6768)
);

CKINVDCx5p33_ASAP7_75t_R g6769 ( 
.A(n_6481),
.Y(n_6769)
);

INVx1_ASAP7_75t_L g6770 ( 
.A(n_6410),
.Y(n_6770)
);

INVx1_ASAP7_75t_L g6771 ( 
.A(n_6427),
.Y(n_6771)
);

INVx1_ASAP7_75t_SL g6772 ( 
.A(n_6179),
.Y(n_6772)
);

BUFx3_ASAP7_75t_L g6773 ( 
.A(n_6466),
.Y(n_6773)
);

CKINVDCx5p33_ASAP7_75t_R g6774 ( 
.A(n_5042),
.Y(n_6774)
);

CKINVDCx20_ASAP7_75t_R g6775 ( 
.A(n_5155),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_6478),
.Y(n_6776)
);

INVx2_ASAP7_75t_L g6777 ( 
.A(n_5273),
.Y(n_6777)
);

CKINVDCx5p33_ASAP7_75t_R g6778 ( 
.A(n_6461),
.Y(n_6778)
);

CKINVDCx5p33_ASAP7_75t_R g6779 ( 
.A(n_6464),
.Y(n_6779)
);

INVx1_ASAP7_75t_L g6780 ( 
.A(n_6462),
.Y(n_6780)
);

CKINVDCx20_ASAP7_75t_R g6781 ( 
.A(n_5162),
.Y(n_6781)
);

CKINVDCx5p33_ASAP7_75t_R g6782 ( 
.A(n_6483),
.Y(n_6782)
);

INVx1_ASAP7_75t_L g6783 ( 
.A(n_6465),
.Y(n_6783)
);

INVx1_ASAP7_75t_L g6784 ( 
.A(n_6472),
.Y(n_6784)
);

INVx2_ASAP7_75t_L g6785 ( 
.A(n_5273),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_6474),
.Y(n_6786)
);

CKINVDCx16_ASAP7_75t_R g6787 ( 
.A(n_5290),
.Y(n_6787)
);

NOR2xp67_ASAP7_75t_L g6788 ( 
.A(n_6468),
.B(n_2),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_6477),
.Y(n_6789)
);

CKINVDCx5p33_ASAP7_75t_R g6790 ( 
.A(n_5046),
.Y(n_6790)
);

INVx1_ASAP7_75t_L g6791 ( 
.A(n_6484),
.Y(n_6791)
);

INVx1_ASAP7_75t_L g6792 ( 
.A(n_5045),
.Y(n_6792)
);

INVx2_ASAP7_75t_L g6793 ( 
.A(n_5273),
.Y(n_6793)
);

BUFx2_ASAP7_75t_L g6794 ( 
.A(n_6257),
.Y(n_6794)
);

INVx1_ASAP7_75t_L g6795 ( 
.A(n_5049),
.Y(n_6795)
);

INVx2_ASAP7_75t_L g6796 ( 
.A(n_5273),
.Y(n_6796)
);

CKINVDCx5p33_ASAP7_75t_R g6797 ( 
.A(n_6451),
.Y(n_6797)
);

BUFx3_ASAP7_75t_L g6798 ( 
.A(n_5290),
.Y(n_6798)
);

INVx1_ASAP7_75t_L g6799 ( 
.A(n_6454),
.Y(n_6799)
);

CKINVDCx5p33_ASAP7_75t_R g6800 ( 
.A(n_6453),
.Y(n_6800)
);

CKINVDCx5p33_ASAP7_75t_R g6801 ( 
.A(n_6458),
.Y(n_6801)
);

INVx1_ASAP7_75t_L g6802 ( 
.A(n_6455),
.Y(n_6802)
);

BUFx2_ASAP7_75t_SL g6803 ( 
.A(n_5797),
.Y(n_6803)
);

INVx2_ASAP7_75t_L g6804 ( 
.A(n_5053),
.Y(n_6804)
);

INVxp67_ASAP7_75t_SL g6805 ( 
.A(n_5577),
.Y(n_6805)
);

CKINVDCx20_ASAP7_75t_R g6806 ( 
.A(n_5185),
.Y(n_6806)
);

CKINVDCx5p33_ASAP7_75t_R g6807 ( 
.A(n_5047),
.Y(n_6807)
);

CKINVDCx5p33_ASAP7_75t_R g6808 ( 
.A(n_5050),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_5060),
.Y(n_6809)
);

BUFx3_ASAP7_75t_L g6810 ( 
.A(n_5363),
.Y(n_6810)
);

INVx1_ASAP7_75t_SL g6811 ( 
.A(n_6306),
.Y(n_6811)
);

INVxp67_ASAP7_75t_L g6812 ( 
.A(n_6328),
.Y(n_6812)
);

INVx2_ASAP7_75t_L g6813 ( 
.A(n_5061),
.Y(n_6813)
);

BUFx3_ASAP7_75t_L g6814 ( 
.A(n_5363),
.Y(n_6814)
);

INVx1_ASAP7_75t_L g6815 ( 
.A(n_6447),
.Y(n_6815)
);

INVx1_ASAP7_75t_L g6816 ( 
.A(n_6457),
.Y(n_6816)
);

INVx1_ASAP7_75t_L g6817 ( 
.A(n_6463),
.Y(n_6817)
);

CKINVDCx5p33_ASAP7_75t_R g6818 ( 
.A(n_6448),
.Y(n_6818)
);

CKINVDCx5p33_ASAP7_75t_R g6819 ( 
.A(n_6450),
.Y(n_6819)
);

CKINVDCx5p33_ASAP7_75t_R g6820 ( 
.A(n_6452),
.Y(n_6820)
);

INVx1_ASAP7_75t_L g6821 ( 
.A(n_5063),
.Y(n_6821)
);

INVx1_ASAP7_75t_L g6822 ( 
.A(n_5071),
.Y(n_6822)
);

CKINVDCx16_ASAP7_75t_R g6823 ( 
.A(n_5405),
.Y(n_6823)
);

INVx1_ASAP7_75t_L g6824 ( 
.A(n_5072),
.Y(n_6824)
);

INVx1_ASAP7_75t_L g6825 ( 
.A(n_5075),
.Y(n_6825)
);

INVx2_ASAP7_75t_L g6826 ( 
.A(n_5078),
.Y(n_6826)
);

INVx1_ASAP7_75t_SL g6827 ( 
.A(n_6329),
.Y(n_6827)
);

INVx1_ASAP7_75t_L g6828 ( 
.A(n_5082),
.Y(n_6828)
);

INVx1_ASAP7_75t_L g6829 ( 
.A(n_5084),
.Y(n_6829)
);

CKINVDCx14_ASAP7_75t_R g6830 ( 
.A(n_6353),
.Y(n_6830)
);

INVx1_ASAP7_75t_L g6831 ( 
.A(n_6441),
.Y(n_6831)
);

INVx1_ASAP7_75t_L g6832 ( 
.A(n_6442),
.Y(n_6832)
);

INVxp67_ASAP7_75t_SL g6833 ( 
.A(n_5742),
.Y(n_6833)
);

INVxp67_ASAP7_75t_L g6834 ( 
.A(n_6469),
.Y(n_6834)
);

CKINVDCx5p33_ASAP7_75t_R g6835 ( 
.A(n_6445),
.Y(n_6835)
);

CKINVDCx5p33_ASAP7_75t_R g6836 ( 
.A(n_6446),
.Y(n_6836)
);

NOR2xp67_ASAP7_75t_L g6837 ( 
.A(n_5709),
.B(n_3),
.Y(n_6837)
);

CKINVDCx20_ASAP7_75t_R g6838 ( 
.A(n_5192),
.Y(n_6838)
);

CKINVDCx5p33_ASAP7_75t_R g6839 ( 
.A(n_5056),
.Y(n_6839)
);

CKINVDCx5p33_ASAP7_75t_R g6840 ( 
.A(n_5059),
.Y(n_6840)
);

CKINVDCx5p33_ASAP7_75t_R g6841 ( 
.A(n_5062),
.Y(n_6841)
);

INVx1_ASAP7_75t_L g6842 ( 
.A(n_5086),
.Y(n_6842)
);

CKINVDCx5p33_ASAP7_75t_R g6843 ( 
.A(n_5064),
.Y(n_6843)
);

CKINVDCx20_ASAP7_75t_R g6844 ( 
.A(n_5235),
.Y(n_6844)
);

INVx2_ASAP7_75t_L g6845 ( 
.A(n_5088),
.Y(n_6845)
);

INVx1_ASAP7_75t_L g6846 ( 
.A(n_5093),
.Y(n_6846)
);

CKINVDCx5p33_ASAP7_75t_R g6847 ( 
.A(n_6435),
.Y(n_6847)
);

BUFx6f_ASAP7_75t_L g6848 ( 
.A(n_5613),
.Y(n_6848)
);

CKINVDCx5p33_ASAP7_75t_R g6849 ( 
.A(n_6437),
.Y(n_6849)
);

CKINVDCx5p33_ASAP7_75t_R g6850 ( 
.A(n_6439),
.Y(n_6850)
);

BUFx5_ASAP7_75t_L g6851 ( 
.A(n_5111),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_6438),
.Y(n_6852)
);

CKINVDCx5p33_ASAP7_75t_R g6853 ( 
.A(n_5066),
.Y(n_6853)
);

INVx1_ASAP7_75t_L g6854 ( 
.A(n_6443),
.Y(n_6854)
);

INVx2_ASAP7_75t_L g6855 ( 
.A(n_5098),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_5106),
.Y(n_6856)
);

INVx1_ASAP7_75t_SL g6857 ( 
.A(n_5279),
.Y(n_6857)
);

INVx1_ASAP7_75t_L g6858 ( 
.A(n_5107),
.Y(n_6858)
);

INVx1_ASAP7_75t_L g6859 ( 
.A(n_5109),
.Y(n_6859)
);

INVx1_ASAP7_75t_L g6860 ( 
.A(n_5114),
.Y(n_6860)
);

BUFx10_ASAP7_75t_L g6861 ( 
.A(n_5842),
.Y(n_6861)
);

CKINVDCx20_ASAP7_75t_R g6862 ( 
.A(n_5258),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_5116),
.Y(n_6863)
);

CKINVDCx5p33_ASAP7_75t_R g6864 ( 
.A(n_6426),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_6429),
.Y(n_6865)
);

INVx2_ASAP7_75t_L g6866 ( 
.A(n_5118),
.Y(n_6866)
);

CKINVDCx5p33_ASAP7_75t_R g6867 ( 
.A(n_6432),
.Y(n_6867)
);

CKINVDCx5p33_ASAP7_75t_R g6868 ( 
.A(n_5069),
.Y(n_6868)
);

INVx2_ASAP7_75t_L g6869 ( 
.A(n_5122),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_5125),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_5138),
.Y(n_6871)
);

CKINVDCx20_ASAP7_75t_R g6872 ( 
.A(n_5272),
.Y(n_6872)
);

INVx1_ASAP7_75t_L g6873 ( 
.A(n_5144),
.Y(n_6873)
);

BUFx2_ASAP7_75t_L g6874 ( 
.A(n_6134),
.Y(n_6874)
);

CKINVDCx5p33_ASAP7_75t_R g6875 ( 
.A(n_5070),
.Y(n_6875)
);

INVx1_ASAP7_75t_L g6876 ( 
.A(n_5145),
.Y(n_6876)
);

INVx1_ASAP7_75t_L g6877 ( 
.A(n_5147),
.Y(n_6877)
);

CKINVDCx5p33_ASAP7_75t_R g6878 ( 
.A(n_5074),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_5149),
.Y(n_6879)
);

INVx1_ASAP7_75t_SL g6880 ( 
.A(n_5551),
.Y(n_6880)
);

CKINVDCx5p33_ASAP7_75t_R g6881 ( 
.A(n_6424),
.Y(n_6881)
);

BUFx6f_ASAP7_75t_L g6882 ( 
.A(n_5613),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_6431),
.Y(n_6883)
);

INVx1_ASAP7_75t_L g6884 ( 
.A(n_6433),
.Y(n_6884)
);

NOR2xp67_ASAP7_75t_L g6885 ( 
.A(n_5833),
.B(n_3),
.Y(n_6885)
);

CKINVDCx5p33_ASAP7_75t_R g6886 ( 
.A(n_6428),
.Y(n_6886)
);

CKINVDCx5p33_ASAP7_75t_R g6887 ( 
.A(n_5076),
.Y(n_6887)
);

CKINVDCx5p33_ASAP7_75t_R g6888 ( 
.A(n_5079),
.Y(n_6888)
);

CKINVDCx14_ASAP7_75t_R g6889 ( 
.A(n_5405),
.Y(n_6889)
);

BUFx5_ASAP7_75t_L g6890 ( 
.A(n_5112),
.Y(n_6890)
);

CKINVDCx5p33_ASAP7_75t_R g6891 ( 
.A(n_5081),
.Y(n_6891)
);

CKINVDCx5p33_ASAP7_75t_R g6892 ( 
.A(n_5083),
.Y(n_6892)
);

CKINVDCx5p33_ASAP7_75t_R g6893 ( 
.A(n_5090),
.Y(n_6893)
);

CKINVDCx5p33_ASAP7_75t_R g6894 ( 
.A(n_5091),
.Y(n_6894)
);

CKINVDCx5p33_ASAP7_75t_R g6895 ( 
.A(n_5092),
.Y(n_6895)
);

INVx1_ASAP7_75t_L g6896 ( 
.A(n_5153),
.Y(n_6896)
);

CKINVDCx5p33_ASAP7_75t_R g6897 ( 
.A(n_6425),
.Y(n_6897)
);

CKINVDCx5p33_ASAP7_75t_R g6898 ( 
.A(n_5094),
.Y(n_6898)
);

INVx1_ASAP7_75t_L g6899 ( 
.A(n_6420),
.Y(n_6899)
);

INVx2_ASAP7_75t_L g6900 ( 
.A(n_5159),
.Y(n_6900)
);

CKINVDCx5p33_ASAP7_75t_R g6901 ( 
.A(n_5095),
.Y(n_6901)
);

CKINVDCx5p33_ASAP7_75t_R g6902 ( 
.A(n_5096),
.Y(n_6902)
);

INVx2_ASAP7_75t_SL g6903 ( 
.A(n_5439),
.Y(n_6903)
);

INVx2_ASAP7_75t_L g6904 ( 
.A(n_5163),
.Y(n_6904)
);

BUFx6f_ASAP7_75t_L g6905 ( 
.A(n_5613),
.Y(n_6905)
);

CKINVDCx5p33_ASAP7_75t_R g6906 ( 
.A(n_5097),
.Y(n_6906)
);

INVx1_ASAP7_75t_L g6907 ( 
.A(n_5164),
.Y(n_6907)
);

BUFx6f_ASAP7_75t_L g6908 ( 
.A(n_5943),
.Y(n_6908)
);

CKINVDCx5p33_ASAP7_75t_R g6909 ( 
.A(n_5100),
.Y(n_6909)
);

CKINVDCx5p33_ASAP7_75t_R g6910 ( 
.A(n_5102),
.Y(n_6910)
);

BUFx6f_ASAP7_75t_L g6911 ( 
.A(n_5943),
.Y(n_6911)
);

INVx1_ASAP7_75t_L g6912 ( 
.A(n_5168),
.Y(n_6912)
);

BUFx2_ASAP7_75t_L g6913 ( 
.A(n_6320),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_5171),
.Y(n_6914)
);

CKINVDCx20_ASAP7_75t_R g6915 ( 
.A(n_5289),
.Y(n_6915)
);

BUFx3_ASAP7_75t_L g6916 ( 
.A(n_5439),
.Y(n_6916)
);

INVx1_ASAP7_75t_L g6917 ( 
.A(n_6423),
.Y(n_6917)
);

BUFx6f_ASAP7_75t_L g6918 ( 
.A(n_5943),
.Y(n_6918)
);

CKINVDCx16_ASAP7_75t_R g6919 ( 
.A(n_6456),
.Y(n_6919)
);

INVx2_ASAP7_75t_SL g6920 ( 
.A(n_5515),
.Y(n_6920)
);

CKINVDCx5p33_ASAP7_75t_R g6921 ( 
.A(n_5108),
.Y(n_6921)
);

CKINVDCx5p33_ASAP7_75t_R g6922 ( 
.A(n_5110),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_5174),
.Y(n_6923)
);

INVx1_ASAP7_75t_L g6924 ( 
.A(n_5180),
.Y(n_6924)
);

INVx1_ASAP7_75t_SL g6925 ( 
.A(n_5483),
.Y(n_6925)
);

CKINVDCx5p33_ASAP7_75t_R g6926 ( 
.A(n_5113),
.Y(n_6926)
);

BUFx5_ASAP7_75t_L g6927 ( 
.A(n_5146),
.Y(n_6927)
);

CKINVDCx5p33_ASAP7_75t_R g6928 ( 
.A(n_5115),
.Y(n_6928)
);

CKINVDCx5p33_ASAP7_75t_R g6929 ( 
.A(n_5117),
.Y(n_6929)
);

INVxp67_ASAP7_75t_L g6930 ( 
.A(n_6347),
.Y(n_6930)
);

CKINVDCx5p33_ASAP7_75t_R g6931 ( 
.A(n_5119),
.Y(n_6931)
);

INVx1_ASAP7_75t_L g6932 ( 
.A(n_5183),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_5186),
.Y(n_6933)
);

CKINVDCx20_ASAP7_75t_R g6934 ( 
.A(n_5305),
.Y(n_6934)
);

CKINVDCx5p33_ASAP7_75t_R g6935 ( 
.A(n_6418),
.Y(n_6935)
);

CKINVDCx5p33_ASAP7_75t_R g6936 ( 
.A(n_5123),
.Y(n_6936)
);

CKINVDCx20_ASAP7_75t_R g6937 ( 
.A(n_5314),
.Y(n_6937)
);

CKINVDCx20_ASAP7_75t_R g6938 ( 
.A(n_5317),
.Y(n_6938)
);

BUFx6f_ASAP7_75t_L g6939 ( 
.A(n_6281),
.Y(n_6939)
);

CKINVDCx5p33_ASAP7_75t_R g6940 ( 
.A(n_5124),
.Y(n_6940)
);

BUFx3_ASAP7_75t_L g6941 ( 
.A(n_5515),
.Y(n_6941)
);

INVx1_ASAP7_75t_L g6942 ( 
.A(n_5195),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_5198),
.Y(n_6943)
);

CKINVDCx5p33_ASAP7_75t_R g6944 ( 
.A(n_5126),
.Y(n_6944)
);

CKINVDCx5p33_ASAP7_75t_R g6945 ( 
.A(n_5127),
.Y(n_6945)
);

CKINVDCx5p33_ASAP7_75t_R g6946 ( 
.A(n_5128),
.Y(n_6946)
);

INVx2_ASAP7_75t_L g6947 ( 
.A(n_5203),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_6848),
.Y(n_6948)
);

CKINVDCx5p33_ASAP7_75t_R g6949 ( 
.A(n_6506),
.Y(n_6949)
);

INVxp33_ASAP7_75t_L g6950 ( 
.A(n_6525),
.Y(n_6950)
);

INVxp67_ASAP7_75t_SL g6951 ( 
.A(n_6512),
.Y(n_6951)
);

INVx1_ASAP7_75t_L g6952 ( 
.A(n_6848),
.Y(n_6952)
);

INVxp33_ASAP7_75t_SL g6953 ( 
.A(n_6491),
.Y(n_6953)
);

INVx1_ASAP7_75t_L g6954 ( 
.A(n_6882),
.Y(n_6954)
);

CKINVDCx20_ASAP7_75t_R g6955 ( 
.A(n_6511),
.Y(n_6955)
);

INVx1_ASAP7_75t_L g6956 ( 
.A(n_6882),
.Y(n_6956)
);

NOR2xp33_ASAP7_75t_L g6957 ( 
.A(n_6495),
.B(n_6419),
.Y(n_6957)
);

INVx1_ASAP7_75t_L g6958 ( 
.A(n_6905),
.Y(n_6958)
);

CKINVDCx5p33_ASAP7_75t_R g6959 ( 
.A(n_6514),
.Y(n_6959)
);

INVx1_ASAP7_75t_L g6960 ( 
.A(n_6905),
.Y(n_6960)
);

INVx1_ASAP7_75t_L g6961 ( 
.A(n_6908),
.Y(n_6961)
);

INVxp67_ASAP7_75t_SL g6962 ( 
.A(n_6541),
.Y(n_6962)
);

CKINVDCx5p33_ASAP7_75t_R g6963 ( 
.A(n_6515),
.Y(n_6963)
);

INVx1_ASAP7_75t_L g6964 ( 
.A(n_6908),
.Y(n_6964)
);

CKINVDCx5p33_ASAP7_75t_R g6965 ( 
.A(n_6517),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6911),
.Y(n_6966)
);

CKINVDCx5p33_ASAP7_75t_R g6967 ( 
.A(n_6519),
.Y(n_6967)
);

INVx1_ASAP7_75t_L g6968 ( 
.A(n_6911),
.Y(n_6968)
);

INVxp33_ASAP7_75t_L g6969 ( 
.A(n_6581),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6918),
.Y(n_6970)
);

INVx1_ASAP7_75t_L g6971 ( 
.A(n_6918),
.Y(n_6971)
);

CKINVDCx5p33_ASAP7_75t_R g6972 ( 
.A(n_6521),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_6939),
.Y(n_6973)
);

CKINVDCx5p33_ASAP7_75t_R g6974 ( 
.A(n_6528),
.Y(n_6974)
);

INVx1_ASAP7_75t_L g6975 ( 
.A(n_6939),
.Y(n_6975)
);

INVxp67_ASAP7_75t_SL g6976 ( 
.A(n_6622),
.Y(n_6976)
);

CKINVDCx5p33_ASAP7_75t_R g6977 ( 
.A(n_6533),
.Y(n_6977)
);

INVxp67_ASAP7_75t_SL g6978 ( 
.A(n_6635),
.Y(n_6978)
);

HB1xp67_ASAP7_75t_L g6979 ( 
.A(n_6717),
.Y(n_6979)
);

CKINVDCx14_ASAP7_75t_R g6980 ( 
.A(n_6889),
.Y(n_6980)
);

INVx1_ASAP7_75t_L g6981 ( 
.A(n_6526),
.Y(n_6981)
);

INVx1_ASAP7_75t_L g6982 ( 
.A(n_6526),
.Y(n_6982)
);

INVx1_ASAP7_75t_L g6983 ( 
.A(n_6554),
.Y(n_6983)
);

INVx1_ASAP7_75t_L g6984 ( 
.A(n_6554),
.Y(n_6984)
);

INVx1_ASAP7_75t_L g6985 ( 
.A(n_6565),
.Y(n_6985)
);

CKINVDCx16_ASAP7_75t_R g6986 ( 
.A(n_6626),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_6565),
.Y(n_6987)
);

INVx1_ASAP7_75t_L g6988 ( 
.A(n_6651),
.Y(n_6988)
);

INVx1_ASAP7_75t_L g6989 ( 
.A(n_6651),
.Y(n_6989)
);

INVx1_ASAP7_75t_L g6990 ( 
.A(n_6589),
.Y(n_6990)
);

INVx2_ASAP7_75t_L g6991 ( 
.A(n_6596),
.Y(n_6991)
);

INVx1_ASAP7_75t_L g6992 ( 
.A(n_6602),
.Y(n_6992)
);

INVx1_ASAP7_75t_L g6993 ( 
.A(n_6628),
.Y(n_6993)
);

CKINVDCx5p33_ASAP7_75t_R g6994 ( 
.A(n_6534),
.Y(n_6994)
);

INVxp33_ASAP7_75t_L g6995 ( 
.A(n_6616),
.Y(n_6995)
);

INVx1_ASAP7_75t_L g6996 ( 
.A(n_6659),
.Y(n_6996)
);

INVx1_ASAP7_75t_L g6997 ( 
.A(n_6663),
.Y(n_6997)
);

INVx2_ASAP7_75t_L g6998 ( 
.A(n_6673),
.Y(n_6998)
);

INVx1_ASAP7_75t_L g6999 ( 
.A(n_6702),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6706),
.Y(n_7000)
);

BUFx2_ASAP7_75t_SL g7001 ( 
.A(n_6604),
.Y(n_7001)
);

INVxp67_ASAP7_75t_SL g7002 ( 
.A(n_6657),
.Y(n_7002)
);

INVx1_ASAP7_75t_L g7003 ( 
.A(n_6606),
.Y(n_7003)
);

INVx1_ASAP7_75t_L g7004 ( 
.A(n_6608),
.Y(n_7004)
);

CKINVDCx5p33_ASAP7_75t_R g7005 ( 
.A(n_6535),
.Y(n_7005)
);

INVxp33_ASAP7_75t_L g7006 ( 
.A(n_6655),
.Y(n_7006)
);

CKINVDCx5p33_ASAP7_75t_R g7007 ( 
.A(n_6538),
.Y(n_7007)
);

INVx1_ASAP7_75t_L g7008 ( 
.A(n_6609),
.Y(n_7008)
);

INVx1_ASAP7_75t_L g7009 ( 
.A(n_6612),
.Y(n_7009)
);

INVx1_ASAP7_75t_L g7010 ( 
.A(n_6613),
.Y(n_7010)
);

INVx1_ASAP7_75t_L g7011 ( 
.A(n_6620),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6624),
.Y(n_7012)
);

CKINVDCx5p33_ASAP7_75t_R g7013 ( 
.A(n_6544),
.Y(n_7013)
);

INVxp67_ASAP7_75t_SL g7014 ( 
.A(n_6709),
.Y(n_7014)
);

INVx1_ASAP7_75t_L g7015 ( 
.A(n_6630),
.Y(n_7015)
);

CKINVDCx16_ASAP7_75t_R g7016 ( 
.A(n_6631),
.Y(n_7016)
);

INVxp67_ASAP7_75t_SL g7017 ( 
.A(n_6671),
.Y(n_7017)
);

INVx1_ASAP7_75t_L g7018 ( 
.A(n_6632),
.Y(n_7018)
);

INVx1_ASAP7_75t_L g7019 ( 
.A(n_6638),
.Y(n_7019)
);

BUFx3_ASAP7_75t_L g7020 ( 
.A(n_6723),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6639),
.Y(n_7021)
);

INVx2_ASAP7_75t_L g7022 ( 
.A(n_6643),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_6645),
.Y(n_7023)
);

BUFx2_ASAP7_75t_L g7024 ( 
.A(n_6721),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6646),
.Y(n_7025)
);

INVx1_ASAP7_75t_L g7026 ( 
.A(n_6653),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_6654),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6656),
.Y(n_7028)
);

HB1xp67_ASAP7_75t_L g7029 ( 
.A(n_6719),
.Y(n_7029)
);

BUFx3_ASAP7_75t_L g7030 ( 
.A(n_6739),
.Y(n_7030)
);

INVxp67_ASAP7_75t_SL g7031 ( 
.A(n_6773),
.Y(n_7031)
);

INVx2_ASAP7_75t_L g7032 ( 
.A(n_6676),
.Y(n_7032)
);

INVx2_ASAP7_75t_L g7033 ( 
.A(n_6677),
.Y(n_7033)
);

INVx1_ASAP7_75t_L g7034 ( 
.A(n_6681),
.Y(n_7034)
);

CKINVDCx20_ASAP7_75t_R g7035 ( 
.A(n_6537),
.Y(n_7035)
);

INVx1_ASAP7_75t_L g7036 ( 
.A(n_6683),
.Y(n_7036)
);

INVx2_ASAP7_75t_L g7037 ( 
.A(n_6684),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6687),
.Y(n_7038)
);

CKINVDCx5p33_ASAP7_75t_R g7039 ( 
.A(n_6545),
.Y(n_7039)
);

CKINVDCx16_ASAP7_75t_R g7040 ( 
.A(n_6640),
.Y(n_7040)
);

CKINVDCx5p33_ASAP7_75t_R g7041 ( 
.A(n_6547),
.Y(n_7041)
);

INVx1_ASAP7_75t_L g7042 ( 
.A(n_6689),
.Y(n_7042)
);

INVx1_ASAP7_75t_L g7043 ( 
.A(n_6691),
.Y(n_7043)
);

BUFx3_ASAP7_75t_L g7044 ( 
.A(n_6733),
.Y(n_7044)
);

INVxp33_ASAP7_75t_SL g7045 ( 
.A(n_6494),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_6693),
.Y(n_7046)
);

INVx2_ASAP7_75t_L g7047 ( 
.A(n_6695),
.Y(n_7047)
);

INVx1_ASAP7_75t_L g7048 ( 
.A(n_6696),
.Y(n_7048)
);

INVx2_ASAP7_75t_L g7049 ( 
.A(n_6699),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_6700),
.Y(n_7050)
);

CKINVDCx20_ASAP7_75t_R g7051 ( 
.A(n_6546),
.Y(n_7051)
);

CKINVDCx5p33_ASAP7_75t_R g7052 ( 
.A(n_6550),
.Y(n_7052)
);

CKINVDCx5p33_ASAP7_75t_R g7053 ( 
.A(n_6552),
.Y(n_7053)
);

NOR2xp33_ASAP7_75t_L g7054 ( 
.A(n_6803),
.B(n_5760),
.Y(n_7054)
);

INVxp67_ASAP7_75t_L g7055 ( 
.A(n_6661),
.Y(n_7055)
);

NOR2xp67_ASAP7_75t_L g7056 ( 
.A(n_6556),
.B(n_5161),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_6704),
.Y(n_7057)
);

BUFx3_ASAP7_75t_L g7058 ( 
.A(n_6733),
.Y(n_7058)
);

INVx1_ASAP7_75t_L g7059 ( 
.A(n_6705),
.Y(n_7059)
);

INVx1_ASAP7_75t_L g7060 ( 
.A(n_6493),
.Y(n_7060)
);

INVx1_ASAP7_75t_L g7061 ( 
.A(n_6502),
.Y(n_7061)
);

INVx1_ASAP7_75t_L g7062 ( 
.A(n_6503),
.Y(n_7062)
);

INVx1_ASAP7_75t_L g7063 ( 
.A(n_6504),
.Y(n_7063)
);

BUFx3_ASAP7_75t_L g7064 ( 
.A(n_6710),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_6507),
.Y(n_7065)
);

BUFx3_ASAP7_75t_L g7066 ( 
.A(n_6712),
.Y(n_7066)
);

INVx2_ASAP7_75t_L g7067 ( 
.A(n_6490),
.Y(n_7067)
);

INVx1_ASAP7_75t_L g7068 ( 
.A(n_6510),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_6516),
.Y(n_7069)
);

CKINVDCx5p33_ASAP7_75t_R g7070 ( 
.A(n_6562),
.Y(n_7070)
);

INVx1_ASAP7_75t_L g7071 ( 
.A(n_6518),
.Y(n_7071)
);

CKINVDCx20_ASAP7_75t_R g7072 ( 
.A(n_6600),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_6522),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_6523),
.Y(n_7074)
);

INVx1_ASAP7_75t_L g7075 ( 
.A(n_6530),
.Y(n_7075)
);

INVx1_ASAP7_75t_L g7076 ( 
.A(n_6531),
.Y(n_7076)
);

INVx1_ASAP7_75t_L g7077 ( 
.A(n_6532),
.Y(n_7077)
);

INVx3_ASAP7_75t_L g7078 ( 
.A(n_6804),
.Y(n_7078)
);

INVxp67_ASAP7_75t_SL g7079 ( 
.A(n_6686),
.Y(n_7079)
);

INVx1_ASAP7_75t_L g7080 ( 
.A(n_6536),
.Y(n_7080)
);

BUFx6f_ASAP7_75t_L g7081 ( 
.A(n_6492),
.Y(n_7081)
);

INVx1_ASAP7_75t_L g7082 ( 
.A(n_6539),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6540),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_6548),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_6551),
.Y(n_7085)
);

INVx1_ASAP7_75t_L g7086 ( 
.A(n_6557),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_6559),
.Y(n_7087)
);

INVxp67_ASAP7_75t_SL g7088 ( 
.A(n_6798),
.Y(n_7088)
);

INVx1_ASAP7_75t_L g7089 ( 
.A(n_6560),
.Y(n_7089)
);

INVx1_ASAP7_75t_L g7090 ( 
.A(n_6561),
.Y(n_7090)
);

INVx1_ASAP7_75t_L g7091 ( 
.A(n_6567),
.Y(n_7091)
);

INVx1_ASAP7_75t_L g7092 ( 
.A(n_6569),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6570),
.Y(n_7093)
);

INVx1_ASAP7_75t_L g7094 ( 
.A(n_6571),
.Y(n_7094)
);

INVx1_ASAP7_75t_L g7095 ( 
.A(n_6572),
.Y(n_7095)
);

INVx2_ASAP7_75t_L g7096 ( 
.A(n_6513),
.Y(n_7096)
);

INVx1_ASAP7_75t_L g7097 ( 
.A(n_6573),
.Y(n_7097)
);

INVx1_ASAP7_75t_L g7098 ( 
.A(n_6575),
.Y(n_7098)
);

INVxp67_ASAP7_75t_SL g7099 ( 
.A(n_6810),
.Y(n_7099)
);

CKINVDCx20_ASAP7_75t_R g7100 ( 
.A(n_6752),
.Y(n_7100)
);

INVxp67_ASAP7_75t_L g7101 ( 
.A(n_6743),
.Y(n_7101)
);

INVxp67_ASAP7_75t_SL g7102 ( 
.A(n_6814),
.Y(n_7102)
);

CKINVDCx20_ASAP7_75t_R g7103 ( 
.A(n_6775),
.Y(n_7103)
);

INVxp67_ASAP7_75t_SL g7104 ( 
.A(n_6916),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_6579),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_6588),
.Y(n_7106)
);

INVx1_ASAP7_75t_L g7107 ( 
.A(n_6594),
.Y(n_7107)
);

INVx1_ASAP7_75t_L g7108 ( 
.A(n_6599),
.Y(n_7108)
);

CKINVDCx20_ASAP7_75t_R g7109 ( 
.A(n_6781),
.Y(n_7109)
);

CKINVDCx20_ASAP7_75t_R g7110 ( 
.A(n_6806),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6603),
.Y(n_7111)
);

CKINVDCx5p33_ASAP7_75t_R g7112 ( 
.A(n_6563),
.Y(n_7112)
);

INVxp67_ASAP7_75t_SL g7113 ( 
.A(n_6941),
.Y(n_7113)
);

CKINVDCx20_ASAP7_75t_R g7114 ( 
.A(n_6838),
.Y(n_7114)
);

INVx2_ASAP7_75t_L g7115 ( 
.A(n_6529),
.Y(n_7115)
);

INVxp33_ASAP7_75t_L g7116 ( 
.A(n_6728),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_6780),
.Y(n_7117)
);

INVx1_ASAP7_75t_L g7118 ( 
.A(n_6783),
.Y(n_7118)
);

INVxp33_ASAP7_75t_SL g7119 ( 
.A(n_6499),
.Y(n_7119)
);

INVx1_ASAP7_75t_L g7120 ( 
.A(n_6784),
.Y(n_7120)
);

INVxp67_ASAP7_75t_SL g7121 ( 
.A(n_6713),
.Y(n_7121)
);

INVx2_ASAP7_75t_L g7122 ( 
.A(n_6543),
.Y(n_7122)
);

INVxp67_ASAP7_75t_SL g7123 ( 
.A(n_6714),
.Y(n_7123)
);

INVx2_ASAP7_75t_L g7124 ( 
.A(n_6549),
.Y(n_7124)
);

BUFx3_ASAP7_75t_L g7125 ( 
.A(n_6718),
.Y(n_7125)
);

INVx1_ASAP7_75t_L g7126 ( 
.A(n_6786),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6789),
.Y(n_7127)
);

INVxp67_ASAP7_75t_SL g7128 ( 
.A(n_6720),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_6791),
.Y(n_7129)
);

INVx1_ASAP7_75t_L g7130 ( 
.A(n_6792),
.Y(n_7130)
);

INVxp67_ASAP7_75t_SL g7131 ( 
.A(n_6724),
.Y(n_7131)
);

INVx1_ASAP7_75t_L g7132 ( 
.A(n_6795),
.Y(n_7132)
);

INVx1_ASAP7_75t_L g7133 ( 
.A(n_6799),
.Y(n_7133)
);

INVxp67_ASAP7_75t_SL g7134 ( 
.A(n_6729),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_6802),
.Y(n_7135)
);

INVxp67_ASAP7_75t_L g7136 ( 
.A(n_6496),
.Y(n_7136)
);

INVx1_ASAP7_75t_L g7137 ( 
.A(n_6809),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_6815),
.Y(n_7138)
);

CKINVDCx20_ASAP7_75t_R g7139 ( 
.A(n_6844),
.Y(n_7139)
);

INVxp67_ASAP7_75t_SL g7140 ( 
.A(n_6730),
.Y(n_7140)
);

INVx1_ASAP7_75t_L g7141 ( 
.A(n_6816),
.Y(n_7141)
);

BUFx2_ASAP7_75t_L g7142 ( 
.A(n_6652),
.Y(n_7142)
);

INVxp33_ASAP7_75t_L g7143 ( 
.A(n_6508),
.Y(n_7143)
);

INVx1_ASAP7_75t_L g7144 ( 
.A(n_6817),
.Y(n_7144)
);

CKINVDCx20_ASAP7_75t_R g7145 ( 
.A(n_6862),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_6821),
.Y(n_7146)
);

CKINVDCx20_ASAP7_75t_R g7147 ( 
.A(n_6872),
.Y(n_7147)
);

CKINVDCx5p33_ASAP7_75t_R g7148 ( 
.A(n_6564),
.Y(n_7148)
);

CKINVDCx5p33_ASAP7_75t_R g7149 ( 
.A(n_6568),
.Y(n_7149)
);

CKINVDCx20_ASAP7_75t_R g7150 ( 
.A(n_6915),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_6822),
.Y(n_7151)
);

BUFx2_ASAP7_75t_L g7152 ( 
.A(n_6694),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_6824),
.Y(n_7153)
);

CKINVDCx5p33_ASAP7_75t_R g7154 ( 
.A(n_6574),
.Y(n_7154)
);

INVx1_ASAP7_75t_L g7155 ( 
.A(n_6825),
.Y(n_7155)
);

CKINVDCx5p33_ASAP7_75t_R g7156 ( 
.A(n_6576),
.Y(n_7156)
);

CKINVDCx5p33_ASAP7_75t_R g7157 ( 
.A(n_6577),
.Y(n_7157)
);

CKINVDCx5p33_ASAP7_75t_R g7158 ( 
.A(n_6578),
.Y(n_7158)
);

CKINVDCx5p33_ASAP7_75t_R g7159 ( 
.A(n_6580),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_6828),
.Y(n_7160)
);

INVx1_ASAP7_75t_L g7161 ( 
.A(n_6829),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_6831),
.Y(n_7162)
);

CKINVDCx5p33_ASAP7_75t_R g7163 ( 
.A(n_6583),
.Y(n_7163)
);

INVx1_ASAP7_75t_L g7164 ( 
.A(n_6832),
.Y(n_7164)
);

INVx1_ASAP7_75t_L g7165 ( 
.A(n_6842),
.Y(n_7165)
);

INVx1_ASAP7_75t_L g7166 ( 
.A(n_6846),
.Y(n_7166)
);

INVx1_ASAP7_75t_L g7167 ( 
.A(n_6852),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_6854),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_6856),
.Y(n_7169)
);

CKINVDCx20_ASAP7_75t_R g7170 ( 
.A(n_6934),
.Y(n_7170)
);

INVx1_ASAP7_75t_L g7171 ( 
.A(n_6858),
.Y(n_7171)
);

INVx1_ASAP7_75t_L g7172 ( 
.A(n_6859),
.Y(n_7172)
);

CKINVDCx20_ASAP7_75t_R g7173 ( 
.A(n_6937),
.Y(n_7173)
);

CKINVDCx5p33_ASAP7_75t_R g7174 ( 
.A(n_6584),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_6860),
.Y(n_7175)
);

INVxp33_ASAP7_75t_L g7176 ( 
.A(n_6553),
.Y(n_7176)
);

INVxp67_ASAP7_75t_SL g7177 ( 
.A(n_6734),
.Y(n_7177)
);

INVx1_ASAP7_75t_L g7178 ( 
.A(n_6863),
.Y(n_7178)
);

CKINVDCx20_ASAP7_75t_R g7179 ( 
.A(n_6938),
.Y(n_7179)
);

CKINVDCx20_ASAP7_75t_R g7180 ( 
.A(n_6597),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_6865),
.Y(n_7181)
);

CKINVDCx5p33_ASAP7_75t_R g7182 ( 
.A(n_6587),
.Y(n_7182)
);

INVx1_ASAP7_75t_L g7183 ( 
.A(n_6870),
.Y(n_7183)
);

BUFx6f_ASAP7_75t_L g7184 ( 
.A(n_6555),
.Y(n_7184)
);

INVx1_ASAP7_75t_L g7185 ( 
.A(n_6871),
.Y(n_7185)
);

CKINVDCx14_ASAP7_75t_R g7186 ( 
.A(n_6830),
.Y(n_7186)
);

INVxp67_ASAP7_75t_L g7187 ( 
.A(n_6498),
.Y(n_7187)
);

INVxp67_ASAP7_75t_L g7188 ( 
.A(n_6520),
.Y(n_7188)
);

CKINVDCx5p33_ASAP7_75t_R g7189 ( 
.A(n_6590),
.Y(n_7189)
);

INVx1_ASAP7_75t_L g7190 ( 
.A(n_6873),
.Y(n_7190)
);

CKINVDCx20_ASAP7_75t_R g7191 ( 
.A(n_6591),
.Y(n_7191)
);

INVx1_ASAP7_75t_L g7192 ( 
.A(n_6876),
.Y(n_7192)
);

INVxp67_ASAP7_75t_SL g7193 ( 
.A(n_6737),
.Y(n_7193)
);

HB1xp67_ASAP7_75t_L g7194 ( 
.A(n_6725),
.Y(n_7194)
);

CKINVDCx5p33_ASAP7_75t_R g7195 ( 
.A(n_6593),
.Y(n_7195)
);

INVx1_ASAP7_75t_L g7196 ( 
.A(n_6877),
.Y(n_7196)
);

CKINVDCx5p33_ASAP7_75t_R g7197 ( 
.A(n_6595),
.Y(n_7197)
);

INVx1_ASAP7_75t_L g7198 ( 
.A(n_6879),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_6883),
.Y(n_7199)
);

INVx1_ASAP7_75t_L g7200 ( 
.A(n_6884),
.Y(n_7200)
);

INVx1_ASAP7_75t_L g7201 ( 
.A(n_6896),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_6899),
.Y(n_7202)
);

INVxp33_ASAP7_75t_SL g7203 ( 
.A(n_6500),
.Y(n_7203)
);

CKINVDCx5p33_ASAP7_75t_R g7204 ( 
.A(n_6598),
.Y(n_7204)
);

INVxp33_ASAP7_75t_L g7205 ( 
.A(n_6585),
.Y(n_7205)
);

INVx1_ASAP7_75t_L g7206 ( 
.A(n_6907),
.Y(n_7206)
);

INVxp67_ASAP7_75t_SL g7207 ( 
.A(n_6741),
.Y(n_7207)
);

CKINVDCx5p33_ASAP7_75t_R g7208 ( 
.A(n_6610),
.Y(n_7208)
);

INVxp33_ASAP7_75t_L g7209 ( 
.A(n_6607),
.Y(n_7209)
);

INVx1_ASAP7_75t_SL g7210 ( 
.A(n_6857),
.Y(n_7210)
);

CKINVDCx20_ASAP7_75t_R g7211 ( 
.A(n_6611),
.Y(n_7211)
);

INVxp67_ASAP7_75t_SL g7212 ( 
.A(n_6742),
.Y(n_7212)
);

CKINVDCx20_ASAP7_75t_R g7213 ( 
.A(n_6615),
.Y(n_7213)
);

INVx1_ASAP7_75t_L g7214 ( 
.A(n_6912),
.Y(n_7214)
);

INVx1_ASAP7_75t_L g7215 ( 
.A(n_6914),
.Y(n_7215)
);

CKINVDCx20_ASAP7_75t_R g7216 ( 
.A(n_6617),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_6917),
.Y(n_7217)
);

CKINVDCx5p33_ASAP7_75t_R g7218 ( 
.A(n_6618),
.Y(n_7218)
);

INVx1_ASAP7_75t_L g7219 ( 
.A(n_6923),
.Y(n_7219)
);

INVxp33_ASAP7_75t_SL g7220 ( 
.A(n_6501),
.Y(n_7220)
);

INVx1_ASAP7_75t_L g7221 ( 
.A(n_6924),
.Y(n_7221)
);

INVx1_ASAP7_75t_L g7222 ( 
.A(n_6932),
.Y(n_7222)
);

INVx1_ASAP7_75t_L g7223 ( 
.A(n_6933),
.Y(n_7223)
);

BUFx3_ASAP7_75t_L g7224 ( 
.A(n_6744),
.Y(n_7224)
);

INVx1_ASAP7_75t_L g7225 ( 
.A(n_6942),
.Y(n_7225)
);

INVxp67_ASAP7_75t_L g7226 ( 
.A(n_6527),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_6943),
.Y(n_7227)
);

INVx1_ASAP7_75t_L g7228 ( 
.A(n_6566),
.Y(n_7228)
);

INVx1_ASAP7_75t_L g7229 ( 
.A(n_6586),
.Y(n_7229)
);

INVx1_ASAP7_75t_L g7230 ( 
.A(n_6813),
.Y(n_7230)
);

BUFx5_ASAP7_75t_L g7231 ( 
.A(n_6745),
.Y(n_7231)
);

CKINVDCx20_ASAP7_75t_R g7232 ( 
.A(n_6619),
.Y(n_7232)
);

CKINVDCx5p33_ASAP7_75t_R g7233 ( 
.A(n_6621),
.Y(n_7233)
);

CKINVDCx20_ASAP7_75t_R g7234 ( 
.A(n_6623),
.Y(n_7234)
);

INVx1_ASAP7_75t_L g7235 ( 
.A(n_6826),
.Y(n_7235)
);

INVx1_ASAP7_75t_L g7236 ( 
.A(n_6845),
.Y(n_7236)
);

CKINVDCx5p33_ASAP7_75t_R g7237 ( 
.A(n_6625),
.Y(n_7237)
);

CKINVDCx20_ASAP7_75t_R g7238 ( 
.A(n_6629),
.Y(n_7238)
);

INVx1_ASAP7_75t_L g7239 ( 
.A(n_6855),
.Y(n_7239)
);

INVx1_ASAP7_75t_L g7240 ( 
.A(n_6866),
.Y(n_7240)
);

INVx1_ASAP7_75t_L g7241 ( 
.A(n_6869),
.Y(n_7241)
);

INVx1_ASAP7_75t_L g7242 ( 
.A(n_6900),
.Y(n_7242)
);

CKINVDCx5p33_ASAP7_75t_R g7243 ( 
.A(n_6636),
.Y(n_7243)
);

INVx1_ASAP7_75t_L g7244 ( 
.A(n_6904),
.Y(n_7244)
);

INVx1_ASAP7_75t_L g7245 ( 
.A(n_6947),
.Y(n_7245)
);

HB1xp67_ASAP7_75t_L g7246 ( 
.A(n_6726),
.Y(n_7246)
);

CKINVDCx20_ASAP7_75t_R g7247 ( 
.A(n_6641),
.Y(n_7247)
);

INVx1_ASAP7_75t_L g7248 ( 
.A(n_6746),
.Y(n_7248)
);

BUFx2_ASAP7_75t_L g7249 ( 
.A(n_6727),
.Y(n_7249)
);

INVx1_ASAP7_75t_L g7250 ( 
.A(n_6751),
.Y(n_7250)
);

INVxp33_ASAP7_75t_L g7251 ( 
.A(n_6633),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_6753),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_6754),
.Y(n_7253)
);

INVx1_ASAP7_75t_L g7254 ( 
.A(n_6755),
.Y(n_7254)
);

INVx1_ASAP7_75t_L g7255 ( 
.A(n_6756),
.Y(n_7255)
);

INVx1_ASAP7_75t_L g7256 ( 
.A(n_6763),
.Y(n_7256)
);

HB1xp67_ASAP7_75t_L g7257 ( 
.A(n_6731),
.Y(n_7257)
);

CKINVDCx5p33_ASAP7_75t_R g7258 ( 
.A(n_6642),
.Y(n_7258)
);

INVx1_ASAP7_75t_L g7259 ( 
.A(n_6764),
.Y(n_7259)
);

INVxp33_ASAP7_75t_SL g7260 ( 
.A(n_6732),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_6767),
.Y(n_7261)
);

CKINVDCx16_ASAP7_75t_R g7262 ( 
.A(n_6768),
.Y(n_7262)
);

INVxp33_ASAP7_75t_SL g7263 ( 
.A(n_6735),
.Y(n_7263)
);

INVx1_ASAP7_75t_SL g7264 ( 
.A(n_6880),
.Y(n_7264)
);

INVxp67_ASAP7_75t_L g7265 ( 
.A(n_6558),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_6770),
.Y(n_7266)
);

CKINVDCx5p33_ASAP7_75t_R g7267 ( 
.A(n_6644),
.Y(n_7267)
);

INVx1_ASAP7_75t_L g7268 ( 
.A(n_6771),
.Y(n_7268)
);

CKINVDCx5p33_ASAP7_75t_R g7269 ( 
.A(n_6647),
.Y(n_7269)
);

INVxp67_ASAP7_75t_SL g7270 ( 
.A(n_6776),
.Y(n_7270)
);

INVx1_ASAP7_75t_L g7271 ( 
.A(n_6748),
.Y(n_7271)
);

CKINVDCx5p33_ASAP7_75t_R g7272 ( 
.A(n_6648),
.Y(n_7272)
);

INVx1_ASAP7_75t_L g7273 ( 
.A(n_6777),
.Y(n_7273)
);

INVx1_ASAP7_75t_L g7274 ( 
.A(n_6785),
.Y(n_7274)
);

INVx1_ASAP7_75t_L g7275 ( 
.A(n_6793),
.Y(n_7275)
);

INVx1_ASAP7_75t_L g7276 ( 
.A(n_6796),
.Y(n_7276)
);

INVx2_ASAP7_75t_L g7277 ( 
.A(n_6592),
.Y(n_7277)
);

CKINVDCx20_ASAP7_75t_R g7278 ( 
.A(n_6649),
.Y(n_7278)
);

BUFx2_ASAP7_75t_L g7279 ( 
.A(n_6736),
.Y(n_7279)
);

CKINVDCx5p33_ASAP7_75t_R g7280 ( 
.A(n_6650),
.Y(n_7280)
);

HB1xp67_ASAP7_75t_L g7281 ( 
.A(n_6740),
.Y(n_7281)
);

CKINVDCx5p33_ASAP7_75t_R g7282 ( 
.A(n_6658),
.Y(n_7282)
);

INVxp67_ASAP7_75t_SL g7283 ( 
.A(n_6601),
.Y(n_7283)
);

INVx1_ASAP7_75t_L g7284 ( 
.A(n_6592),
.Y(n_7284)
);

INVx2_ASAP7_75t_L g7285 ( 
.A(n_6592),
.Y(n_7285)
);

CKINVDCx5p33_ASAP7_75t_R g7286 ( 
.A(n_6660),
.Y(n_7286)
);

INVx1_ASAP7_75t_L g7287 ( 
.A(n_6592),
.Y(n_7287)
);

BUFx2_ASAP7_75t_L g7288 ( 
.A(n_6946),
.Y(n_7288)
);

INVx1_ASAP7_75t_L g7289 ( 
.A(n_6665),
.Y(n_7289)
);

INVx1_ASAP7_75t_L g7290 ( 
.A(n_6665),
.Y(n_7290)
);

CKINVDCx5p33_ASAP7_75t_R g7291 ( 
.A(n_6662),
.Y(n_7291)
);

INVx2_ASAP7_75t_L g7292 ( 
.A(n_6665),
.Y(n_7292)
);

BUFx3_ASAP7_75t_L g7293 ( 
.A(n_6666),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_6665),
.Y(n_7294)
);

INVx2_ASAP7_75t_L g7295 ( 
.A(n_6851),
.Y(n_7295)
);

INVx1_ASAP7_75t_L g7296 ( 
.A(n_6851),
.Y(n_7296)
);

CKINVDCx5p33_ASAP7_75t_R g7297 ( 
.A(n_6667),
.Y(n_7297)
);

INVx1_ASAP7_75t_L g7298 ( 
.A(n_6851),
.Y(n_7298)
);

BUFx6f_ASAP7_75t_L g7299 ( 
.A(n_6747),
.Y(n_7299)
);

CKINVDCx16_ASAP7_75t_R g7300 ( 
.A(n_6787),
.Y(n_7300)
);

INVx1_ASAP7_75t_L g7301 ( 
.A(n_6851),
.Y(n_7301)
);

INVx1_ASAP7_75t_L g7302 ( 
.A(n_6890),
.Y(n_7302)
);

CKINVDCx5p33_ASAP7_75t_R g7303 ( 
.A(n_6669),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_6890),
.Y(n_7304)
);

INVxp67_ASAP7_75t_SL g7305 ( 
.A(n_6930),
.Y(n_7305)
);

CKINVDCx5p33_ASAP7_75t_R g7306 ( 
.A(n_6670),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_6890),
.Y(n_7307)
);

HB1xp67_ASAP7_75t_L g7308 ( 
.A(n_6749),
.Y(n_7308)
);

CKINVDCx5p33_ASAP7_75t_R g7309 ( 
.A(n_6674),
.Y(n_7309)
);

INVx1_ASAP7_75t_L g7310 ( 
.A(n_6890),
.Y(n_7310)
);

INVxp33_ASAP7_75t_SL g7311 ( 
.A(n_6678),
.Y(n_7311)
);

INVx1_ASAP7_75t_L g7312 ( 
.A(n_6927),
.Y(n_7312)
);

INVxp33_ASAP7_75t_SL g7313 ( 
.A(n_6679),
.Y(n_7313)
);

INVx2_ASAP7_75t_L g7314 ( 
.A(n_6927),
.Y(n_7314)
);

BUFx3_ASAP7_75t_L g7315 ( 
.A(n_6680),
.Y(n_7315)
);

INVx1_ASAP7_75t_L g7316 ( 
.A(n_6927),
.Y(n_7316)
);

CKINVDCx20_ASAP7_75t_R g7317 ( 
.A(n_6682),
.Y(n_7317)
);

INVx1_ASAP7_75t_L g7318 ( 
.A(n_6927),
.Y(n_7318)
);

BUFx6f_ASAP7_75t_L g7319 ( 
.A(n_6750),
.Y(n_7319)
);

INVx1_ASAP7_75t_L g7320 ( 
.A(n_6701),
.Y(n_7320)
);

INVx1_ASAP7_75t_L g7321 ( 
.A(n_6805),
.Y(n_7321)
);

HB1xp67_ASAP7_75t_L g7322 ( 
.A(n_6757),
.Y(n_7322)
);

BUFx2_ASAP7_75t_L g7323 ( 
.A(n_6758),
.Y(n_7323)
);

HB1xp67_ASAP7_75t_L g7324 ( 
.A(n_6759),
.Y(n_7324)
);

CKINVDCx20_ASAP7_75t_R g7325 ( 
.A(n_6685),
.Y(n_7325)
);

INVxp67_ASAP7_75t_SL g7326 ( 
.A(n_6833),
.Y(n_7326)
);

CKINVDCx5p33_ASAP7_75t_R g7327 ( 
.A(n_6690),
.Y(n_7327)
);

INVx1_ASAP7_75t_L g7328 ( 
.A(n_6945),
.Y(n_7328)
);

INVx1_ASAP7_75t_L g7329 ( 
.A(n_6760),
.Y(n_7329)
);

CKINVDCx5p33_ASAP7_75t_R g7330 ( 
.A(n_6697),
.Y(n_7330)
);

INVx1_ASAP7_75t_L g7331 ( 
.A(n_6761),
.Y(n_7331)
);

INVx1_ASAP7_75t_L g7332 ( 
.A(n_6944),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_6762),
.Y(n_7333)
);

INVx1_ASAP7_75t_L g7334 ( 
.A(n_6940),
.Y(n_7334)
);

CKINVDCx20_ASAP7_75t_R g7335 ( 
.A(n_6698),
.Y(n_7335)
);

CKINVDCx20_ASAP7_75t_R g7336 ( 
.A(n_6703),
.Y(n_7336)
);

INVxp33_ASAP7_75t_SL g7337 ( 
.A(n_6707),
.Y(n_7337)
);

CKINVDCx5p33_ASAP7_75t_R g7338 ( 
.A(n_6708),
.Y(n_7338)
);

INVx1_ASAP7_75t_L g7339 ( 
.A(n_6766),
.Y(n_7339)
);

INVxp67_ASAP7_75t_SL g7340 ( 
.A(n_6505),
.Y(n_7340)
);

INVxp67_ASAP7_75t_SL g7341 ( 
.A(n_6497),
.Y(n_7341)
);

CKINVDCx5p33_ASAP7_75t_R g7342 ( 
.A(n_6711),
.Y(n_7342)
);

INVx1_ASAP7_75t_L g7343 ( 
.A(n_6769),
.Y(n_7343)
);

INVxp67_ASAP7_75t_L g7344 ( 
.A(n_6582),
.Y(n_7344)
);

INVxp67_ASAP7_75t_SL g7345 ( 
.A(n_6509),
.Y(n_7345)
);

INVx1_ASAP7_75t_L g7346 ( 
.A(n_6936),
.Y(n_7346)
);

INVx1_ASAP7_75t_L g7347 ( 
.A(n_6774),
.Y(n_7347)
);

INVx1_ASAP7_75t_L g7348 ( 
.A(n_6935),
.Y(n_7348)
);

INVx1_ASAP7_75t_L g7349 ( 
.A(n_6778),
.Y(n_7349)
);

CKINVDCx5p33_ASAP7_75t_R g7350 ( 
.A(n_6715),
.Y(n_7350)
);

INVxp33_ASAP7_75t_SL g7351 ( 
.A(n_6716),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_6931),
.Y(n_7352)
);

INVx2_ASAP7_75t_L g7353 ( 
.A(n_6779),
.Y(n_7353)
);

INVxp67_ASAP7_75t_SL g7354 ( 
.A(n_6542),
.Y(n_7354)
);

INVx1_ASAP7_75t_L g7355 ( 
.A(n_6782),
.Y(n_7355)
);

INVx1_ASAP7_75t_L g7356 ( 
.A(n_6929),
.Y(n_7356)
);

INVx2_ASAP7_75t_L g7357 ( 
.A(n_6790),
.Y(n_7357)
);

HB1xp67_ASAP7_75t_L g7358 ( 
.A(n_6797),
.Y(n_7358)
);

INVxp67_ASAP7_75t_SL g7359 ( 
.A(n_6738),
.Y(n_7359)
);

CKINVDCx5p33_ASAP7_75t_R g7360 ( 
.A(n_6800),
.Y(n_7360)
);

INVx1_ASAP7_75t_L g7361 ( 
.A(n_6801),
.Y(n_7361)
);

INVx1_ASAP7_75t_L g7362 ( 
.A(n_6928),
.Y(n_7362)
);

INVx1_ASAP7_75t_L g7363 ( 
.A(n_6807),
.Y(n_7363)
);

INVxp67_ASAP7_75t_SL g7364 ( 
.A(n_6812),
.Y(n_7364)
);

INVx1_ASAP7_75t_L g7365 ( 
.A(n_6808),
.Y(n_7365)
);

BUFx3_ASAP7_75t_L g7366 ( 
.A(n_6818),
.Y(n_7366)
);

CKINVDCx20_ASAP7_75t_R g7367 ( 
.A(n_6524),
.Y(n_7367)
);

INVxp33_ASAP7_75t_SL g7368 ( 
.A(n_6819),
.Y(n_7368)
);

INVx1_ASAP7_75t_L g7369 ( 
.A(n_6820),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_6926),
.Y(n_7370)
);

INVx1_ASAP7_75t_L g7371 ( 
.A(n_6835),
.Y(n_7371)
);

BUFx3_ASAP7_75t_L g7372 ( 
.A(n_6836),
.Y(n_7372)
);

CKINVDCx20_ASAP7_75t_R g7373 ( 
.A(n_6925),
.Y(n_7373)
);

BUFx5_ASAP7_75t_L g7374 ( 
.A(n_6614),
.Y(n_7374)
);

INVx1_ASAP7_75t_L g7375 ( 
.A(n_6839),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_6922),
.Y(n_7376)
);

INVxp67_ASAP7_75t_L g7377 ( 
.A(n_6664),
.Y(n_7377)
);

CKINVDCx5p33_ASAP7_75t_R g7378 ( 
.A(n_6840),
.Y(n_7378)
);

INVx1_ASAP7_75t_L g7379 ( 
.A(n_6841),
.Y(n_7379)
);

INVxp67_ASAP7_75t_SL g7380 ( 
.A(n_6834),
.Y(n_7380)
);

INVx1_ASAP7_75t_L g7381 ( 
.A(n_6843),
.Y(n_7381)
);

BUFx3_ASAP7_75t_L g7382 ( 
.A(n_6847),
.Y(n_7382)
);

INVx1_ASAP7_75t_L g7383 ( 
.A(n_6849),
.Y(n_7383)
);

INVx1_ASAP7_75t_L g7384 ( 
.A(n_6921),
.Y(n_7384)
);

CKINVDCx20_ASAP7_75t_R g7385 ( 
.A(n_6850),
.Y(n_7385)
);

CKINVDCx20_ASAP7_75t_R g7386 ( 
.A(n_6853),
.Y(n_7386)
);

INVx1_ASAP7_75t_L g7387 ( 
.A(n_6864),
.Y(n_7387)
);

INVxp67_ASAP7_75t_SL g7388 ( 
.A(n_6627),
.Y(n_7388)
);

INVx1_ASAP7_75t_L g7389 ( 
.A(n_6867),
.Y(n_7389)
);

INVx1_ASAP7_75t_L g7390 ( 
.A(n_6868),
.Y(n_7390)
);

CKINVDCx5p33_ASAP7_75t_R g7391 ( 
.A(n_6875),
.Y(n_7391)
);

INVx1_ASAP7_75t_L g7392 ( 
.A(n_6878),
.Y(n_7392)
);

INVxp67_ASAP7_75t_SL g7393 ( 
.A(n_6634),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_6881),
.Y(n_7394)
);

INVxp67_ASAP7_75t_L g7395 ( 
.A(n_6903),
.Y(n_7395)
);

INVx1_ASAP7_75t_L g7396 ( 
.A(n_6886),
.Y(n_7396)
);

INVx2_ASAP7_75t_L g7397 ( 
.A(n_6887),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_6888),
.Y(n_7398)
);

CKINVDCx5p33_ASAP7_75t_R g7399 ( 
.A(n_6891),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_6892),
.Y(n_7400)
);

INVx1_ASAP7_75t_L g7401 ( 
.A(n_6893),
.Y(n_7401)
);

CKINVDCx20_ASAP7_75t_R g7402 ( 
.A(n_6894),
.Y(n_7402)
);

INVx1_ASAP7_75t_L g7403 ( 
.A(n_6895),
.Y(n_7403)
);

HB1xp67_ASAP7_75t_L g7404 ( 
.A(n_6897),
.Y(n_7404)
);

CKINVDCx5p33_ASAP7_75t_R g7405 ( 
.A(n_6898),
.Y(n_7405)
);

INVx1_ASAP7_75t_SL g7406 ( 
.A(n_6672),
.Y(n_7406)
);

CKINVDCx5p33_ASAP7_75t_R g7407 ( 
.A(n_6901),
.Y(n_7407)
);

CKINVDCx20_ASAP7_75t_R g7408 ( 
.A(n_6902),
.Y(n_7408)
);

INVx1_ASAP7_75t_L g7409 ( 
.A(n_6906),
.Y(n_7409)
);

INVxp33_ASAP7_75t_L g7410 ( 
.A(n_6765),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_6909),
.Y(n_7411)
);

INVx1_ASAP7_75t_L g7412 ( 
.A(n_6910),
.Y(n_7412)
);

INVx1_ASAP7_75t_L g7413 ( 
.A(n_6637),
.Y(n_7413)
);

INVx1_ASAP7_75t_L g7414 ( 
.A(n_6788),
.Y(n_7414)
);

CKINVDCx5p33_ASAP7_75t_R g7415 ( 
.A(n_6605),
.Y(n_7415)
);

INVx1_ASAP7_75t_L g7416 ( 
.A(n_6837),
.Y(n_7416)
);

INVxp67_ASAP7_75t_SL g7417 ( 
.A(n_6885),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_6920),
.Y(n_7418)
);

INVx1_ASAP7_75t_L g7419 ( 
.A(n_6874),
.Y(n_7419)
);

HB1xp67_ASAP7_75t_L g7420 ( 
.A(n_6675),
.Y(n_7420)
);

INVxp67_ASAP7_75t_L g7421 ( 
.A(n_6794),
.Y(n_7421)
);

INVx3_ASAP7_75t_L g7422 ( 
.A(n_6861),
.Y(n_7422)
);

INVx1_ASAP7_75t_L g7423 ( 
.A(n_6913),
.Y(n_7423)
);

INVx1_ASAP7_75t_L g7424 ( 
.A(n_6668),
.Y(n_7424)
);

CKINVDCx20_ASAP7_75t_R g7425 ( 
.A(n_6823),
.Y(n_7425)
);

CKINVDCx5p33_ASAP7_75t_R g7426 ( 
.A(n_6919),
.Y(n_7426)
);

INVx2_ASAP7_75t_L g7427 ( 
.A(n_6688),
.Y(n_7427)
);

INVx2_ASAP7_75t_SL g7428 ( 
.A(n_6692),
.Y(n_7428)
);

INVx2_ASAP7_75t_L g7429 ( 
.A(n_6722),
.Y(n_7429)
);

INVx1_ASAP7_75t_L g7430 ( 
.A(n_6772),
.Y(n_7430)
);

CKINVDCx5p33_ASAP7_75t_R g7431 ( 
.A(n_6811),
.Y(n_7431)
);

CKINVDCx20_ASAP7_75t_R g7432 ( 
.A(n_6827),
.Y(n_7432)
);

INVx1_ASAP7_75t_L g7433 ( 
.A(n_6848),
.Y(n_7433)
);

BUFx3_ASAP7_75t_L g7434 ( 
.A(n_6512),
.Y(n_7434)
);

CKINVDCx5p33_ASAP7_75t_R g7435 ( 
.A(n_6506),
.Y(n_7435)
);

INVx2_ASAP7_75t_L g7436 ( 
.A(n_6589),
.Y(n_7436)
);

CKINVDCx20_ASAP7_75t_R g7437 ( 
.A(n_6511),
.Y(n_7437)
);

INVxp33_ASAP7_75t_L g7438 ( 
.A(n_6525),
.Y(n_7438)
);

INVxp33_ASAP7_75t_L g7439 ( 
.A(n_6525),
.Y(n_7439)
);

BUFx6f_ASAP7_75t_L g7440 ( 
.A(n_6526),
.Y(n_7440)
);

INVxp67_ASAP7_75t_L g7441 ( 
.A(n_6525),
.Y(n_7441)
);

INVx1_ASAP7_75t_L g7442 ( 
.A(n_6848),
.Y(n_7442)
);

INVx1_ASAP7_75t_L g7443 ( 
.A(n_6848),
.Y(n_7443)
);

INVxp67_ASAP7_75t_SL g7444 ( 
.A(n_6512),
.Y(n_7444)
);

CKINVDCx20_ASAP7_75t_R g7445 ( 
.A(n_6511),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_6848),
.Y(n_7446)
);

INVx1_ASAP7_75t_L g7447 ( 
.A(n_6848),
.Y(n_7447)
);

INVx1_ASAP7_75t_L g7448 ( 
.A(n_6848),
.Y(n_7448)
);

NOR2xp33_ASAP7_75t_L g7449 ( 
.A(n_6495),
.B(n_5260),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_6848),
.Y(n_7450)
);

BUFx6f_ASAP7_75t_L g7451 ( 
.A(n_6526),
.Y(n_7451)
);

CKINVDCx16_ASAP7_75t_R g7452 ( 
.A(n_6626),
.Y(n_7452)
);

CKINVDCx20_ASAP7_75t_R g7453 ( 
.A(n_6511),
.Y(n_7453)
);

INVx2_ASAP7_75t_L g7454 ( 
.A(n_6589),
.Y(n_7454)
);

CKINVDCx5p33_ASAP7_75t_R g7455 ( 
.A(n_6506),
.Y(n_7455)
);

INVx1_ASAP7_75t_L g7456 ( 
.A(n_6848),
.Y(n_7456)
);

CKINVDCx5p33_ASAP7_75t_R g7457 ( 
.A(n_6506),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_6848),
.Y(n_7458)
);

INVx1_ASAP7_75t_L g7459 ( 
.A(n_6848),
.Y(n_7459)
);

INVxp67_ASAP7_75t_SL g7460 ( 
.A(n_6512),
.Y(n_7460)
);

INVx1_ASAP7_75t_L g7461 ( 
.A(n_6848),
.Y(n_7461)
);

INVx2_ASAP7_75t_L g7462 ( 
.A(n_6589),
.Y(n_7462)
);

INVx1_ASAP7_75t_L g7463 ( 
.A(n_6848),
.Y(n_7463)
);

INVxp67_ASAP7_75t_L g7464 ( 
.A(n_6525),
.Y(n_7464)
);

CKINVDCx5p33_ASAP7_75t_R g7465 ( 
.A(n_6506),
.Y(n_7465)
);

INVx1_ASAP7_75t_L g7466 ( 
.A(n_6848),
.Y(n_7466)
);

INVx1_ASAP7_75t_L g7467 ( 
.A(n_6848),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_6848),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_6848),
.Y(n_7469)
);

INVx1_ASAP7_75t_L g7470 ( 
.A(n_6848),
.Y(n_7470)
);

BUFx6f_ASAP7_75t_SL g7471 ( 
.A(n_6496),
.Y(n_7471)
);

INVx1_ASAP7_75t_L g7472 ( 
.A(n_6848),
.Y(n_7472)
);

BUFx2_ASAP7_75t_L g7473 ( 
.A(n_7432),
.Y(n_7473)
);

AND2x4_ASAP7_75t_L g7474 ( 
.A(n_7434),
.B(n_5052),
.Y(n_7474)
);

INVx2_ASAP7_75t_L g7475 ( 
.A(n_7081),
.Y(n_7475)
);

INVxp67_ASAP7_75t_L g7476 ( 
.A(n_7420),
.Y(n_7476)
);

NAND2xp5_ASAP7_75t_L g7477 ( 
.A(n_7014),
.B(n_5323),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_7117),
.Y(n_7478)
);

AND2x2_ASAP7_75t_L g7479 ( 
.A(n_7427),
.B(n_5538),
.Y(n_7479)
);

INVx2_ASAP7_75t_L g7480 ( 
.A(n_7081),
.Y(n_7480)
);

INVx2_ASAP7_75t_L g7481 ( 
.A(n_7081),
.Y(n_7481)
);

NAND2xp5_ASAP7_75t_L g7482 ( 
.A(n_7283),
.B(n_5765),
.Y(n_7482)
);

BUFx3_ASAP7_75t_L g7483 ( 
.A(n_7020),
.Y(n_7483)
);

NAND2xp5_ASAP7_75t_L g7484 ( 
.A(n_7388),
.B(n_6111),
.Y(n_7484)
);

BUFx2_ASAP7_75t_L g7485 ( 
.A(n_7431),
.Y(n_7485)
);

BUFx2_ASAP7_75t_L g7486 ( 
.A(n_7406),
.Y(n_7486)
);

INVx5_ASAP7_75t_L g7487 ( 
.A(n_7422),
.Y(n_7487)
);

BUFx6f_ASAP7_75t_L g7488 ( 
.A(n_7440),
.Y(n_7488)
);

AOI22xp5_ASAP7_75t_L g7489 ( 
.A1(n_6957),
.A2(n_5262),
.B1(n_6375),
.B2(n_5085),
.Y(n_7489)
);

BUFx6f_ASAP7_75t_L g7490 ( 
.A(n_7440),
.Y(n_7490)
);

AND2x4_ASAP7_75t_L g7491 ( 
.A(n_6951),
.B(n_5148),
.Y(n_7491)
);

INVx1_ASAP7_75t_L g7492 ( 
.A(n_7118),
.Y(n_7492)
);

NAND2xp5_ASAP7_75t_L g7493 ( 
.A(n_7393),
.B(n_5233),
.Y(n_7493)
);

AOI22xp5_ASAP7_75t_L g7494 ( 
.A1(n_7449),
.A2(n_5103),
.B1(n_5121),
.B2(n_5048),
.Y(n_7494)
);

INVx3_ASAP7_75t_L g7495 ( 
.A(n_7044),
.Y(n_7495)
);

OAI22xp5_ASAP7_75t_L g7496 ( 
.A1(n_7079),
.A2(n_7328),
.B1(n_7331),
.B2(n_7329),
.Y(n_7496)
);

OAI22xp5_ASAP7_75t_SL g7497 ( 
.A1(n_7373),
.A2(n_5329),
.B1(n_5384),
.B2(n_5368),
.Y(n_7497)
);

INVx2_ASAP7_75t_L g7498 ( 
.A(n_7184),
.Y(n_7498)
);

BUFx6f_ASAP7_75t_L g7499 ( 
.A(n_7440),
.Y(n_7499)
);

INVx1_ASAP7_75t_L g7500 ( 
.A(n_7120),
.Y(n_7500)
);

HB1xp67_ASAP7_75t_L g7501 ( 
.A(n_7428),
.Y(n_7501)
);

BUFx6f_ASAP7_75t_L g7502 ( 
.A(n_7451),
.Y(n_7502)
);

BUFx6f_ASAP7_75t_L g7503 ( 
.A(n_7451),
.Y(n_7503)
);

INVx3_ASAP7_75t_L g7504 ( 
.A(n_7058),
.Y(n_7504)
);

NAND2xp5_ASAP7_75t_L g7505 ( 
.A(n_7417),
.B(n_5243),
.Y(n_7505)
);

BUFx6f_ASAP7_75t_L g7506 ( 
.A(n_7451),
.Y(n_7506)
);

AND2x6_ASAP7_75t_L g7507 ( 
.A(n_7299),
.B(n_5297),
.Y(n_7507)
);

CKINVDCx5p33_ASAP7_75t_R g7508 ( 
.A(n_6949),
.Y(n_7508)
);

INVx1_ASAP7_75t_L g7509 ( 
.A(n_7126),
.Y(n_7509)
);

AND2x4_ASAP7_75t_L g7510 ( 
.A(n_6962),
.B(n_5172),
.Y(n_7510)
);

BUFx8_ASAP7_75t_L g7511 ( 
.A(n_7471),
.Y(n_7511)
);

INVx2_ASAP7_75t_L g7512 ( 
.A(n_7184),
.Y(n_7512)
);

INVx3_ASAP7_75t_L g7513 ( 
.A(n_7030),
.Y(n_7513)
);

OAI22xp5_ASAP7_75t_L g7514 ( 
.A1(n_7332),
.A2(n_6068),
.B1(n_5961),
.B2(n_5130),
.Y(n_7514)
);

INVx2_ASAP7_75t_L g7515 ( 
.A(n_7184),
.Y(n_7515)
);

OAI21x1_ASAP7_75t_L g7516 ( 
.A1(n_7277),
.A2(n_5542),
.B(n_5416),
.Y(n_7516)
);

BUFx6f_ASAP7_75t_L g7517 ( 
.A(n_7064),
.Y(n_7517)
);

INVx3_ASAP7_75t_L g7518 ( 
.A(n_7066),
.Y(n_7518)
);

INVx2_ASAP7_75t_L g7519 ( 
.A(n_6991),
.Y(n_7519)
);

BUFx2_ASAP7_75t_L g7520 ( 
.A(n_7429),
.Y(n_7520)
);

NAND2xp5_ASAP7_75t_L g7521 ( 
.A(n_7056),
.B(n_5251),
.Y(n_7521)
);

BUFx6f_ASAP7_75t_L g7522 ( 
.A(n_7125),
.Y(n_7522)
);

BUFx6f_ASAP7_75t_L g7523 ( 
.A(n_7224),
.Y(n_7523)
);

INVx2_ASAP7_75t_L g7524 ( 
.A(n_6998),
.Y(n_7524)
);

INVx3_ASAP7_75t_L g7525 ( 
.A(n_7067),
.Y(n_7525)
);

INVx3_ASAP7_75t_L g7526 ( 
.A(n_7096),
.Y(n_7526)
);

INVx2_ASAP7_75t_L g7527 ( 
.A(n_7436),
.Y(n_7527)
);

AND2x2_ASAP7_75t_L g7528 ( 
.A(n_7116),
.B(n_5538),
.Y(n_7528)
);

NOR2xp33_ASAP7_75t_SL g7529 ( 
.A(n_7368),
.B(n_5960),
.Y(n_7529)
);

NAND2xp33_ASAP7_75t_L g7530 ( 
.A(n_7353),
.B(n_6281),
.Y(n_7530)
);

BUFx8_ASAP7_75t_L g7531 ( 
.A(n_7471),
.Y(n_7531)
);

INVx6_ASAP7_75t_L g7532 ( 
.A(n_7262),
.Y(n_7532)
);

OAI22xp5_ASAP7_75t_L g7533 ( 
.A1(n_7333),
.A2(n_5131),
.B1(n_5132),
.B2(n_5129),
.Y(n_7533)
);

BUFx2_ASAP7_75t_L g7534 ( 
.A(n_7210),
.Y(n_7534)
);

INVx3_ASAP7_75t_L g7535 ( 
.A(n_7115),
.Y(n_7535)
);

HB1xp67_ASAP7_75t_L g7536 ( 
.A(n_7264),
.Y(n_7536)
);

INVx2_ASAP7_75t_L g7537 ( 
.A(n_7454),
.Y(n_7537)
);

INVx2_ASAP7_75t_L g7538 ( 
.A(n_7462),
.Y(n_7538)
);

INVx1_ASAP7_75t_L g7539 ( 
.A(n_7127),
.Y(n_7539)
);

INVx3_ASAP7_75t_L g7540 ( 
.A(n_7122),
.Y(n_7540)
);

BUFx2_ASAP7_75t_L g7541 ( 
.A(n_7430),
.Y(n_7541)
);

INVx5_ASAP7_75t_L g7542 ( 
.A(n_7422),
.Y(n_7542)
);

NAND2xp5_ASAP7_75t_L g7543 ( 
.A(n_7340),
.B(n_5267),
.Y(n_7543)
);

OA21x2_ASAP7_75t_L g7544 ( 
.A1(n_7285),
.A2(n_6092),
.B(n_5338),
.Y(n_7544)
);

INVx1_ASAP7_75t_L g7545 ( 
.A(n_7129),
.Y(n_7545)
);

AND2x2_ASAP7_75t_L g7546 ( 
.A(n_7054),
.B(n_5587),
.Y(n_7546)
);

CKINVDCx5p33_ASAP7_75t_R g7547 ( 
.A(n_6959),
.Y(n_7547)
);

INVx2_ASAP7_75t_L g7548 ( 
.A(n_7124),
.Y(n_7548)
);

INVx1_ASAP7_75t_L g7549 ( 
.A(n_7130),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7132),
.Y(n_7550)
);

OAI21x1_ASAP7_75t_L g7551 ( 
.A1(n_7292),
.A2(n_5358),
.B(n_5271),
.Y(n_7551)
);

BUFx6f_ASAP7_75t_L g7552 ( 
.A(n_6948),
.Y(n_7552)
);

INVx2_ASAP7_75t_L g7553 ( 
.A(n_7022),
.Y(n_7553)
);

INVx2_ASAP7_75t_L g7554 ( 
.A(n_7032),
.Y(n_7554)
);

BUFx2_ASAP7_75t_L g7555 ( 
.A(n_7180),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_7133),
.Y(n_7556)
);

BUFx6f_ASAP7_75t_L g7557 ( 
.A(n_7472),
.Y(n_7557)
);

BUFx2_ASAP7_75t_L g7558 ( 
.A(n_7425),
.Y(n_7558)
);

INVx3_ASAP7_75t_L g7559 ( 
.A(n_6952),
.Y(n_7559)
);

INVx3_ASAP7_75t_L g7560 ( 
.A(n_6954),
.Y(n_7560)
);

INVx1_ASAP7_75t_L g7561 ( 
.A(n_7135),
.Y(n_7561)
);

INVx1_ASAP7_75t_L g7562 ( 
.A(n_7137),
.Y(n_7562)
);

OAI21x1_ASAP7_75t_L g7563 ( 
.A1(n_7295),
.A2(n_7314),
.B(n_7287),
.Y(n_7563)
);

BUFx8_ASAP7_75t_SL g7564 ( 
.A(n_7415),
.Y(n_7564)
);

INVx2_ASAP7_75t_L g7565 ( 
.A(n_7033),
.Y(n_7565)
);

NAND2xp5_ASAP7_75t_L g7566 ( 
.A(n_7231),
.B(n_5361),
.Y(n_7566)
);

INVx2_ASAP7_75t_L g7567 ( 
.A(n_7037),
.Y(n_7567)
);

HB1xp67_ASAP7_75t_L g7568 ( 
.A(n_7421),
.Y(n_7568)
);

CKINVDCx5p33_ASAP7_75t_R g7569 ( 
.A(n_6963),
.Y(n_7569)
);

HB1xp67_ASAP7_75t_L g7570 ( 
.A(n_7055),
.Y(n_7570)
);

INVx2_ASAP7_75t_L g7571 ( 
.A(n_7047),
.Y(n_7571)
);

OAI21x1_ASAP7_75t_L g7572 ( 
.A1(n_7284),
.A2(n_5549),
.B(n_5400),
.Y(n_7572)
);

AOI22xp5_ASAP7_75t_L g7573 ( 
.A1(n_7326),
.A2(n_5352),
.B1(n_5398),
.B2(n_5339),
.Y(n_7573)
);

NAND2xp5_ASAP7_75t_L g7574 ( 
.A(n_7231),
.B(n_7060),
.Y(n_7574)
);

INVx2_ASAP7_75t_L g7575 ( 
.A(n_7049),
.Y(n_7575)
);

INVx2_ASAP7_75t_L g7576 ( 
.A(n_7228),
.Y(n_7576)
);

INVx2_ASAP7_75t_L g7577 ( 
.A(n_7229),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_7138),
.Y(n_7578)
);

INVxp67_ASAP7_75t_L g7579 ( 
.A(n_7424),
.Y(n_7579)
);

NAND2xp5_ASAP7_75t_L g7580 ( 
.A(n_7231),
.B(n_5580),
.Y(n_7580)
);

INVx2_ASAP7_75t_L g7581 ( 
.A(n_7003),
.Y(n_7581)
);

BUFx6f_ASAP7_75t_L g7582 ( 
.A(n_6956),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_7141),
.Y(n_7583)
);

BUFx6f_ASAP7_75t_L g7584 ( 
.A(n_6958),
.Y(n_7584)
);

OAI21x1_ASAP7_75t_L g7585 ( 
.A1(n_7289),
.A2(n_5641),
.B(n_5598),
.Y(n_7585)
);

CKINVDCx20_ASAP7_75t_R g7586 ( 
.A(n_6955),
.Y(n_7586)
);

HB1xp67_ASAP7_75t_L g7587 ( 
.A(n_7101),
.Y(n_7587)
);

BUFx3_ASAP7_75t_L g7588 ( 
.A(n_7367),
.Y(n_7588)
);

AND2x2_ASAP7_75t_L g7589 ( 
.A(n_7305),
.B(n_5587),
.Y(n_7589)
);

INVx2_ASAP7_75t_L g7590 ( 
.A(n_7004),
.Y(n_7590)
);

OAI22xp5_ASAP7_75t_L g7591 ( 
.A1(n_7334),
.A2(n_5137),
.B1(n_5139),
.B2(n_5135),
.Y(n_7591)
);

AND2x2_ASAP7_75t_L g7592 ( 
.A(n_7341),
.B(n_5595),
.Y(n_7592)
);

INVx1_ASAP7_75t_L g7593 ( 
.A(n_7144),
.Y(n_7593)
);

INVx2_ASAP7_75t_L g7594 ( 
.A(n_7008),
.Y(n_7594)
);

INVx2_ASAP7_75t_L g7595 ( 
.A(n_7009),
.Y(n_7595)
);

AND2x2_ASAP7_75t_L g7596 ( 
.A(n_7345),
.B(n_5595),
.Y(n_7596)
);

AOI22xp5_ASAP7_75t_L g7597 ( 
.A1(n_7354),
.A2(n_5450),
.B1(n_5479),
.B2(n_5440),
.Y(n_7597)
);

INVx2_ASAP7_75t_L g7598 ( 
.A(n_7010),
.Y(n_7598)
);

HB1xp67_ASAP7_75t_L g7599 ( 
.A(n_7441),
.Y(n_7599)
);

BUFx8_ASAP7_75t_L g7600 ( 
.A(n_7024),
.Y(n_7600)
);

INVx5_ASAP7_75t_L g7601 ( 
.A(n_7299),
.Y(n_7601)
);

OA21x2_ASAP7_75t_L g7602 ( 
.A1(n_7290),
.A2(n_5748),
.B(n_5744),
.Y(n_7602)
);

INVx2_ASAP7_75t_SL g7603 ( 
.A(n_7419),
.Y(n_7603)
);

NOR2xp33_ASAP7_75t_SL g7604 ( 
.A(n_7260),
.B(n_5387),
.Y(n_7604)
);

NAND2xp5_ASAP7_75t_L g7605 ( 
.A(n_7231),
.B(n_5750),
.Y(n_7605)
);

BUFx6f_ASAP7_75t_L g7606 ( 
.A(n_6960),
.Y(n_7606)
);

INVx2_ASAP7_75t_L g7607 ( 
.A(n_7011),
.Y(n_7607)
);

AOI22x1_ASAP7_75t_SL g7608 ( 
.A1(n_7035),
.A2(n_5420),
.B1(n_5455),
.B2(n_5388),
.Y(n_7608)
);

INVx1_ASAP7_75t_L g7609 ( 
.A(n_7146),
.Y(n_7609)
);

AND2x6_ASAP7_75t_L g7610 ( 
.A(n_7299),
.B(n_5501),
.Y(n_7610)
);

BUFx3_ASAP7_75t_L g7611 ( 
.A(n_7293),
.Y(n_7611)
);

BUFx3_ASAP7_75t_L g7612 ( 
.A(n_7315),
.Y(n_7612)
);

BUFx6f_ASAP7_75t_L g7613 ( 
.A(n_7470),
.Y(n_7613)
);

INVx1_ASAP7_75t_L g7614 ( 
.A(n_7151),
.Y(n_7614)
);

HB1xp67_ASAP7_75t_L g7615 ( 
.A(n_7464),
.Y(n_7615)
);

INVx1_ASAP7_75t_L g7616 ( 
.A(n_7153),
.Y(n_7616)
);

INVx1_ASAP7_75t_L g7617 ( 
.A(n_7155),
.Y(n_7617)
);

INVx2_ASAP7_75t_L g7618 ( 
.A(n_7012),
.Y(n_7618)
);

INVx4_ASAP7_75t_L g7619 ( 
.A(n_7319),
.Y(n_7619)
);

INVx3_ASAP7_75t_L g7620 ( 
.A(n_6961),
.Y(n_7620)
);

BUFx6f_ASAP7_75t_L g7621 ( 
.A(n_6964),
.Y(n_7621)
);

NAND2xp5_ASAP7_75t_L g7622 ( 
.A(n_7231),
.B(n_5759),
.Y(n_7622)
);

INVx3_ASAP7_75t_L g7623 ( 
.A(n_6966),
.Y(n_7623)
);

INVx2_ASAP7_75t_L g7624 ( 
.A(n_7015),
.Y(n_7624)
);

HB1xp67_ASAP7_75t_L g7625 ( 
.A(n_7188),
.Y(n_7625)
);

AND2x6_ASAP7_75t_L g7626 ( 
.A(n_7319),
.B(n_5516),
.Y(n_7626)
);

INVx2_ASAP7_75t_L g7627 ( 
.A(n_7018),
.Y(n_7627)
);

BUFx8_ASAP7_75t_L g7628 ( 
.A(n_7142),
.Y(n_7628)
);

INVxp67_ASAP7_75t_L g7629 ( 
.A(n_7359),
.Y(n_7629)
);

BUFx6f_ASAP7_75t_L g7630 ( 
.A(n_6968),
.Y(n_7630)
);

OAI22x1_ASAP7_75t_SL g7631 ( 
.A1(n_7100),
.A2(n_5491),
.B1(n_5499),
.B2(n_5468),
.Y(n_7631)
);

INVx1_ASAP7_75t_L g7632 ( 
.A(n_7160),
.Y(n_7632)
);

OAI22xp5_ASAP7_75t_L g7633 ( 
.A1(n_7339),
.A2(n_5142),
.B1(n_5143),
.B2(n_5141),
.Y(n_7633)
);

NOR2xp33_ASAP7_75t_L g7634 ( 
.A(n_7343),
.B(n_5373),
.Y(n_7634)
);

NAND2xp5_ASAP7_75t_L g7635 ( 
.A(n_7061),
.B(n_5810),
.Y(n_7635)
);

INVx2_ASAP7_75t_L g7636 ( 
.A(n_7019),
.Y(n_7636)
);

BUFx6f_ASAP7_75t_L g7637 ( 
.A(n_7469),
.Y(n_7637)
);

INVx1_ASAP7_75t_L g7638 ( 
.A(n_7161),
.Y(n_7638)
);

INVx3_ASAP7_75t_L g7639 ( 
.A(n_6970),
.Y(n_7639)
);

BUFx6f_ASAP7_75t_L g7640 ( 
.A(n_6971),
.Y(n_7640)
);

CKINVDCx6p67_ASAP7_75t_R g7641 ( 
.A(n_7300),
.Y(n_7641)
);

AND2x4_ASAP7_75t_L g7642 ( 
.A(n_6976),
.B(n_5413),
.Y(n_7642)
);

INVx6_ASAP7_75t_L g7643 ( 
.A(n_7319),
.Y(n_7643)
);

INVx2_ASAP7_75t_L g7644 ( 
.A(n_7021),
.Y(n_7644)
);

INVx2_ASAP7_75t_L g7645 ( 
.A(n_7023),
.Y(n_7645)
);

NAND2xp5_ASAP7_75t_L g7646 ( 
.A(n_7062),
.B(n_5848),
.Y(n_7646)
);

INVx2_ASAP7_75t_L g7647 ( 
.A(n_7025),
.Y(n_7647)
);

CKINVDCx11_ASAP7_75t_R g7648 ( 
.A(n_7103),
.Y(n_7648)
);

BUFx6f_ASAP7_75t_L g7649 ( 
.A(n_7468),
.Y(n_7649)
);

BUFx3_ASAP7_75t_L g7650 ( 
.A(n_7191),
.Y(n_7650)
);

INVx1_ASAP7_75t_L g7651 ( 
.A(n_7162),
.Y(n_7651)
);

OA21x2_ASAP7_75t_L g7652 ( 
.A1(n_7294),
.A2(n_5856),
.B(n_5853),
.Y(n_7652)
);

INVx2_ASAP7_75t_L g7653 ( 
.A(n_7026),
.Y(n_7653)
);

INVx1_ASAP7_75t_L g7654 ( 
.A(n_7164),
.Y(n_7654)
);

INVx1_ASAP7_75t_L g7655 ( 
.A(n_7165),
.Y(n_7655)
);

INVx3_ASAP7_75t_L g7656 ( 
.A(n_6973),
.Y(n_7656)
);

INVx2_ASAP7_75t_L g7657 ( 
.A(n_7027),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_7166),
.Y(n_7658)
);

BUFx6f_ASAP7_75t_L g7659 ( 
.A(n_7467),
.Y(n_7659)
);

NAND2xp5_ASAP7_75t_L g7660 ( 
.A(n_7063),
.B(n_5875),
.Y(n_7660)
);

INVx4_ASAP7_75t_L g7661 ( 
.A(n_6965),
.Y(n_7661)
);

BUFx6f_ASAP7_75t_L g7662 ( 
.A(n_6975),
.Y(n_7662)
);

BUFx6f_ASAP7_75t_L g7663 ( 
.A(n_7466),
.Y(n_7663)
);

AND2x4_ASAP7_75t_L g7664 ( 
.A(n_6978),
.B(n_5461),
.Y(n_7664)
);

BUFx12f_ASAP7_75t_L g7665 ( 
.A(n_7426),
.Y(n_7665)
);

HB1xp67_ASAP7_75t_L g7666 ( 
.A(n_7226),
.Y(n_7666)
);

INVx3_ASAP7_75t_L g7667 ( 
.A(n_7433),
.Y(n_7667)
);

BUFx6f_ASAP7_75t_L g7668 ( 
.A(n_7442),
.Y(n_7668)
);

OA21x2_ASAP7_75t_L g7669 ( 
.A1(n_7296),
.A2(n_7301),
.B(n_7298),
.Y(n_7669)
);

INVx1_ASAP7_75t_L g7670 ( 
.A(n_7167),
.Y(n_7670)
);

NAND2xp5_ASAP7_75t_L g7671 ( 
.A(n_7065),
.B(n_5883),
.Y(n_7671)
);

BUFx8_ASAP7_75t_SL g7672 ( 
.A(n_7109),
.Y(n_7672)
);

BUFx3_ASAP7_75t_L g7673 ( 
.A(n_7211),
.Y(n_7673)
);

NAND2xp5_ASAP7_75t_L g7674 ( 
.A(n_7068),
.B(n_5887),
.Y(n_7674)
);

AND2x6_ASAP7_75t_L g7675 ( 
.A(n_7346),
.B(n_5527),
.Y(n_7675)
);

INVx1_ASAP7_75t_L g7676 ( 
.A(n_7168),
.Y(n_7676)
);

NOR2xp33_ASAP7_75t_L g7677 ( 
.A(n_7347),
.B(n_5521),
.Y(n_7677)
);

BUFx6f_ASAP7_75t_L g7678 ( 
.A(n_7443),
.Y(n_7678)
);

INVx1_ASAP7_75t_L g7679 ( 
.A(n_7169),
.Y(n_7679)
);

BUFx8_ASAP7_75t_L g7680 ( 
.A(n_7152),
.Y(n_7680)
);

INVx1_ASAP7_75t_L g7681 ( 
.A(n_7171),
.Y(n_7681)
);

BUFx6f_ASAP7_75t_L g7682 ( 
.A(n_7446),
.Y(n_7682)
);

HB1xp67_ASAP7_75t_L g7683 ( 
.A(n_7265),
.Y(n_7683)
);

INVx1_ASAP7_75t_L g7684 ( 
.A(n_7172),
.Y(n_7684)
);

BUFx12f_ASAP7_75t_L g7685 ( 
.A(n_7360),
.Y(n_7685)
);

BUFx6f_ASAP7_75t_L g7686 ( 
.A(n_7447),
.Y(n_7686)
);

AND2x2_ASAP7_75t_L g7687 ( 
.A(n_7364),
.B(n_5627),
.Y(n_7687)
);

BUFx6f_ASAP7_75t_L g7688 ( 
.A(n_7448),
.Y(n_7688)
);

AND2x2_ASAP7_75t_SL g7689 ( 
.A(n_7249),
.B(n_5068),
.Y(n_7689)
);

BUFx6f_ASAP7_75t_L g7690 ( 
.A(n_7450),
.Y(n_7690)
);

INVxp33_ASAP7_75t_SL g7691 ( 
.A(n_7378),
.Y(n_7691)
);

AND2x4_ASAP7_75t_L g7692 ( 
.A(n_7002),
.B(n_7444),
.Y(n_7692)
);

CKINVDCx5p33_ASAP7_75t_R g7693 ( 
.A(n_6967),
.Y(n_7693)
);

BUFx6f_ASAP7_75t_L g7694 ( 
.A(n_7456),
.Y(n_7694)
);

INVx2_ASAP7_75t_L g7695 ( 
.A(n_7028),
.Y(n_7695)
);

INVx1_ASAP7_75t_L g7696 ( 
.A(n_7175),
.Y(n_7696)
);

AOI22xp5_ASAP7_75t_L g7697 ( 
.A1(n_7380),
.A2(n_5597),
.B1(n_5616),
.B2(n_5529),
.Y(n_7697)
);

NAND2xp5_ASAP7_75t_L g7698 ( 
.A(n_7069),
.B(n_7071),
.Y(n_7698)
);

NAND2xp5_ASAP7_75t_L g7699 ( 
.A(n_7073),
.B(n_5932),
.Y(n_7699)
);

INVx3_ASAP7_75t_L g7700 ( 
.A(n_7458),
.Y(n_7700)
);

INVx2_ASAP7_75t_L g7701 ( 
.A(n_7034),
.Y(n_7701)
);

AND2x4_ASAP7_75t_L g7702 ( 
.A(n_7460),
.B(n_5541),
.Y(n_7702)
);

INVx2_ASAP7_75t_L g7703 ( 
.A(n_7036),
.Y(n_7703)
);

INVx1_ASAP7_75t_L g7704 ( 
.A(n_7178),
.Y(n_7704)
);

INVx2_ASAP7_75t_L g7705 ( 
.A(n_7038),
.Y(n_7705)
);

AND2x2_ASAP7_75t_L g7706 ( 
.A(n_7186),
.B(n_5627),
.Y(n_7706)
);

BUFx6f_ASAP7_75t_L g7707 ( 
.A(n_7459),
.Y(n_7707)
);

INVx1_ASAP7_75t_L g7708 ( 
.A(n_7181),
.Y(n_7708)
);

AND2x6_ASAP7_75t_L g7709 ( 
.A(n_7348),
.B(n_5649),
.Y(n_7709)
);

AND2x4_ASAP7_75t_L g7710 ( 
.A(n_7017),
.B(n_5552),
.Y(n_7710)
);

AND2x4_ASAP7_75t_L g7711 ( 
.A(n_7031),
.B(n_7088),
.Y(n_7711)
);

HB1xp67_ASAP7_75t_L g7712 ( 
.A(n_7344),
.Y(n_7712)
);

INVx1_ASAP7_75t_L g7713 ( 
.A(n_7183),
.Y(n_7713)
);

BUFx2_ASAP7_75t_L g7714 ( 
.A(n_7385),
.Y(n_7714)
);

BUFx8_ASAP7_75t_SL g7715 ( 
.A(n_7110),
.Y(n_7715)
);

HB1xp67_ASAP7_75t_L g7716 ( 
.A(n_7377),
.Y(n_7716)
);

INVx2_ASAP7_75t_L g7717 ( 
.A(n_7042),
.Y(n_7717)
);

BUFx2_ASAP7_75t_L g7718 ( 
.A(n_7386),
.Y(n_7718)
);

INVx2_ASAP7_75t_L g7719 ( 
.A(n_7043),
.Y(n_7719)
);

BUFx6f_ASAP7_75t_L g7720 ( 
.A(n_7461),
.Y(n_7720)
);

AND2x2_ASAP7_75t_L g7721 ( 
.A(n_6980),
.B(n_5686),
.Y(n_7721)
);

NAND2xp5_ASAP7_75t_L g7722 ( 
.A(n_7074),
.B(n_5982),
.Y(n_7722)
);

AND2x4_ASAP7_75t_L g7723 ( 
.A(n_7099),
.B(n_7102),
.Y(n_7723)
);

INVx2_ASAP7_75t_L g7724 ( 
.A(n_7046),
.Y(n_7724)
);

INVx2_ASAP7_75t_L g7725 ( 
.A(n_7048),
.Y(n_7725)
);

OAI22xp5_ASAP7_75t_SL g7726 ( 
.A1(n_7402),
.A2(n_5519),
.B1(n_5533),
.B2(n_5517),
.Y(n_7726)
);

BUFx3_ASAP7_75t_L g7727 ( 
.A(n_7213),
.Y(n_7727)
);

BUFx8_ASAP7_75t_L g7728 ( 
.A(n_7279),
.Y(n_7728)
);

BUFx6f_ASAP7_75t_L g7729 ( 
.A(n_7463),
.Y(n_7729)
);

NAND2xp5_ASAP7_75t_L g7730 ( 
.A(n_7075),
.B(n_7076),
.Y(n_7730)
);

CKINVDCx6p67_ASAP7_75t_R g7731 ( 
.A(n_6986),
.Y(n_7731)
);

INVx3_ASAP7_75t_L g7732 ( 
.A(n_7078),
.Y(n_7732)
);

BUFx6f_ASAP7_75t_L g7733 ( 
.A(n_6981),
.Y(n_7733)
);

AOI22xp5_ASAP7_75t_L g7734 ( 
.A1(n_7349),
.A2(n_5788),
.B1(n_5792),
.B2(n_5754),
.Y(n_7734)
);

NOR2xp33_ASAP7_75t_L g7735 ( 
.A(n_7352),
.B(n_5588),
.Y(n_7735)
);

INVx3_ASAP7_75t_L g7736 ( 
.A(n_7078),
.Y(n_7736)
);

INVx1_ASAP7_75t_L g7737 ( 
.A(n_7185),
.Y(n_7737)
);

INVx3_ASAP7_75t_L g7738 ( 
.A(n_6982),
.Y(n_7738)
);

BUFx2_ASAP7_75t_L g7739 ( 
.A(n_7408),
.Y(n_7739)
);

BUFx3_ASAP7_75t_L g7740 ( 
.A(n_7216),
.Y(n_7740)
);

BUFx6f_ASAP7_75t_L g7741 ( 
.A(n_6983),
.Y(n_7741)
);

INVx1_ASAP7_75t_L g7742 ( 
.A(n_7190),
.Y(n_7742)
);

BUFx6f_ASAP7_75t_L g7743 ( 
.A(n_6984),
.Y(n_7743)
);

INVx2_ASAP7_75t_L g7744 ( 
.A(n_7050),
.Y(n_7744)
);

NAND2xp5_ASAP7_75t_SL g7745 ( 
.A(n_7374),
.B(n_5152),
.Y(n_7745)
);

INVx2_ASAP7_75t_L g7746 ( 
.A(n_7057),
.Y(n_7746)
);

INVx2_ASAP7_75t_SL g7747 ( 
.A(n_7423),
.Y(n_7747)
);

HB1xp67_ASAP7_75t_L g7748 ( 
.A(n_7395),
.Y(n_7748)
);

INVx1_ASAP7_75t_L g7749 ( 
.A(n_7192),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7196),
.Y(n_7750)
);

AOI22xp5_ASAP7_75t_SL g7751 ( 
.A1(n_7232),
.A2(n_5617),
.B1(n_5620),
.B2(n_5574),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_7198),
.Y(n_7752)
);

AND2x4_ASAP7_75t_L g7753 ( 
.A(n_7104),
.B(n_7113),
.Y(n_7753)
);

INVx6_ASAP7_75t_L g7754 ( 
.A(n_7016),
.Y(n_7754)
);

AND2x4_ASAP7_75t_L g7755 ( 
.A(n_7357),
.B(n_7397),
.Y(n_7755)
);

OA21x2_ASAP7_75t_L g7756 ( 
.A1(n_7302),
.A2(n_6117),
.B(n_6069),
.Y(n_7756)
);

AOI22xp5_ASAP7_75t_L g7757 ( 
.A1(n_7355),
.A2(n_5855),
.B1(n_5890),
.B2(n_5812),
.Y(n_7757)
);

INVx2_ASAP7_75t_L g7758 ( 
.A(n_7059),
.Y(n_7758)
);

INVx2_ASAP7_75t_L g7759 ( 
.A(n_6990),
.Y(n_7759)
);

CKINVDCx5p33_ASAP7_75t_R g7760 ( 
.A(n_6972),
.Y(n_7760)
);

OA21x2_ASAP7_75t_L g7761 ( 
.A1(n_7304),
.A2(n_6260),
.B(n_6135),
.Y(n_7761)
);

NAND2x1p5_ASAP7_75t_L g7762 ( 
.A(n_7366),
.B(n_7372),
.Y(n_7762)
);

INVx1_ASAP7_75t_L g7763 ( 
.A(n_7199),
.Y(n_7763)
);

INVx5_ASAP7_75t_L g7764 ( 
.A(n_7288),
.Y(n_7764)
);

INVx5_ASAP7_75t_L g7765 ( 
.A(n_7323),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_7200),
.Y(n_7766)
);

AOI22xp5_ASAP7_75t_L g7767 ( 
.A1(n_7356),
.A2(n_5901),
.B1(n_5957),
.B2(n_5893),
.Y(n_7767)
);

CKINVDCx6p67_ASAP7_75t_R g7768 ( 
.A(n_7040),
.Y(n_7768)
);

BUFx6f_ASAP7_75t_L g7769 ( 
.A(n_6985),
.Y(n_7769)
);

NAND2xp5_ASAP7_75t_L g7770 ( 
.A(n_7077),
.B(n_7080),
.Y(n_7770)
);

AND2x2_ASAP7_75t_L g7771 ( 
.A(n_7136),
.B(n_5686),
.Y(n_7771)
);

INVx1_ASAP7_75t_L g7772 ( 
.A(n_7201),
.Y(n_7772)
);

OAI21x1_ASAP7_75t_L g7773 ( 
.A1(n_7307),
.A2(n_6291),
.B(n_6270),
.Y(n_7773)
);

INVx2_ASAP7_75t_L g7774 ( 
.A(n_6992),
.Y(n_7774)
);

INVx2_ASAP7_75t_SL g7775 ( 
.A(n_6979),
.Y(n_7775)
);

INVx2_ASAP7_75t_L g7776 ( 
.A(n_6993),
.Y(n_7776)
);

INVx3_ASAP7_75t_L g7777 ( 
.A(n_6987),
.Y(n_7777)
);

OA21x2_ASAP7_75t_L g7778 ( 
.A1(n_7310),
.A2(n_6319),
.B(n_6299),
.Y(n_7778)
);

AND2x4_ASAP7_75t_L g7779 ( 
.A(n_7361),
.B(n_5745),
.Y(n_7779)
);

BUFx2_ASAP7_75t_L g7780 ( 
.A(n_7187),
.Y(n_7780)
);

BUFx6f_ASAP7_75t_L g7781 ( 
.A(n_6988),
.Y(n_7781)
);

BUFx6f_ASAP7_75t_L g7782 ( 
.A(n_6989),
.Y(n_7782)
);

INVx1_ASAP7_75t_L g7783 ( 
.A(n_7202),
.Y(n_7783)
);

INVx2_ASAP7_75t_L g7784 ( 
.A(n_6996),
.Y(n_7784)
);

INVx1_ASAP7_75t_L g7785 ( 
.A(n_7206),
.Y(n_7785)
);

INVx2_ASAP7_75t_L g7786 ( 
.A(n_6997),
.Y(n_7786)
);

AND2x4_ASAP7_75t_L g7787 ( 
.A(n_7362),
.B(n_7363),
.Y(n_7787)
);

INVx3_ASAP7_75t_L g7788 ( 
.A(n_7214),
.Y(n_7788)
);

AND2x2_ASAP7_75t_L g7789 ( 
.A(n_7143),
.B(n_5886),
.Y(n_7789)
);

BUFx12f_ASAP7_75t_L g7790 ( 
.A(n_7391),
.Y(n_7790)
);

OAI22xp5_ASAP7_75t_L g7791 ( 
.A1(n_7365),
.A2(n_5154),
.B1(n_5158),
.B2(n_5157),
.Y(n_7791)
);

BUFx6f_ASAP7_75t_L g7792 ( 
.A(n_7215),
.Y(n_7792)
);

BUFx6f_ASAP7_75t_L g7793 ( 
.A(n_7217),
.Y(n_7793)
);

NAND2xp5_ASAP7_75t_L g7794 ( 
.A(n_7082),
.B(n_6336),
.Y(n_7794)
);

INVx2_ASAP7_75t_L g7795 ( 
.A(n_6999),
.Y(n_7795)
);

INVx2_ASAP7_75t_L g7796 ( 
.A(n_7000),
.Y(n_7796)
);

BUFx6f_ASAP7_75t_L g7797 ( 
.A(n_7219),
.Y(n_7797)
);

HB1xp67_ASAP7_75t_L g7798 ( 
.A(n_6950),
.Y(n_7798)
);

HB1xp67_ASAP7_75t_L g7799 ( 
.A(n_6969),
.Y(n_7799)
);

AND2x4_ASAP7_75t_L g7800 ( 
.A(n_7369),
.B(n_5826),
.Y(n_7800)
);

AOI22xp5_ASAP7_75t_L g7801 ( 
.A1(n_7370),
.A2(n_6007),
.B1(n_6029),
.B2(n_5988),
.Y(n_7801)
);

BUFx6f_ASAP7_75t_L g7802 ( 
.A(n_7221),
.Y(n_7802)
);

BUFx6f_ASAP7_75t_L g7803 ( 
.A(n_7222),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_7223),
.Y(n_7804)
);

AOI22xp5_ASAP7_75t_L g7805 ( 
.A1(n_7371),
.A2(n_6081),
.B1(n_6102),
.B2(n_6056),
.Y(n_7805)
);

AND2x2_ASAP7_75t_SL g7806 ( 
.A(n_7452),
.B(n_5120),
.Y(n_7806)
);

BUFx2_ASAP7_75t_L g7807 ( 
.A(n_7114),
.Y(n_7807)
);

INVx1_ASAP7_75t_L g7808 ( 
.A(n_7225),
.Y(n_7808)
);

BUFx6f_ASAP7_75t_L g7809 ( 
.A(n_7227),
.Y(n_7809)
);

INVx2_ASAP7_75t_L g7810 ( 
.A(n_7271),
.Y(n_7810)
);

NAND2xp5_ASAP7_75t_L g7811 ( 
.A(n_7083),
.B(n_7084),
.Y(n_7811)
);

AND2x4_ASAP7_75t_L g7812 ( 
.A(n_7375),
.B(n_5926),
.Y(n_7812)
);

OA21x2_ASAP7_75t_L g7813 ( 
.A1(n_7312),
.A2(n_5215),
.B(n_5207),
.Y(n_7813)
);

AND2x4_ASAP7_75t_L g7814 ( 
.A(n_7376),
.B(n_6037),
.Y(n_7814)
);

INVx2_ASAP7_75t_L g7815 ( 
.A(n_7273),
.Y(n_7815)
);

INVx1_ASAP7_75t_L g7816 ( 
.A(n_7085),
.Y(n_7816)
);

BUFx3_ASAP7_75t_L g7817 ( 
.A(n_7234),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_7086),
.Y(n_7818)
);

CKINVDCx5p33_ASAP7_75t_R g7819 ( 
.A(n_6974),
.Y(n_7819)
);

INVx2_ASAP7_75t_L g7820 ( 
.A(n_7274),
.Y(n_7820)
);

INVx2_ASAP7_75t_L g7821 ( 
.A(n_7275),
.Y(n_7821)
);

OAI22xp5_ASAP7_75t_L g7822 ( 
.A1(n_7379),
.A2(n_5165),
.B1(n_5166),
.B2(n_5160),
.Y(n_7822)
);

INVx2_ASAP7_75t_L g7823 ( 
.A(n_7276),
.Y(n_7823)
);

BUFx3_ASAP7_75t_L g7824 ( 
.A(n_7238),
.Y(n_7824)
);

AND2x2_ASAP7_75t_SL g7825 ( 
.A(n_7029),
.B(n_5193),
.Y(n_7825)
);

BUFx6f_ASAP7_75t_L g7826 ( 
.A(n_7087),
.Y(n_7826)
);

HB1xp67_ASAP7_75t_L g7827 ( 
.A(n_6995),
.Y(n_7827)
);

INVx3_ASAP7_75t_L g7828 ( 
.A(n_7107),
.Y(n_7828)
);

INVx2_ASAP7_75t_L g7829 ( 
.A(n_7230),
.Y(n_7829)
);

BUFx8_ASAP7_75t_L g7830 ( 
.A(n_7374),
.Y(n_7830)
);

INVx2_ASAP7_75t_SL g7831 ( 
.A(n_7194),
.Y(n_7831)
);

CKINVDCx5p33_ASAP7_75t_R g7832 ( 
.A(n_6977),
.Y(n_7832)
);

NOR2xp33_ASAP7_75t_SL g7833 ( 
.A(n_7263),
.B(n_5639),
.Y(n_7833)
);

BUFx3_ASAP7_75t_L g7834 ( 
.A(n_7247),
.Y(n_7834)
);

NAND2xp5_ASAP7_75t_L g7835 ( 
.A(n_7089),
.B(n_6281),
.Y(n_7835)
);

BUFx6f_ASAP7_75t_L g7836 ( 
.A(n_7090),
.Y(n_7836)
);

INVx1_ASAP7_75t_L g7837 ( 
.A(n_7091),
.Y(n_7837)
);

OA21x2_ASAP7_75t_L g7838 ( 
.A1(n_7316),
.A2(n_5219),
.B(n_5218),
.Y(n_7838)
);

INVx1_ASAP7_75t_L g7839 ( 
.A(n_7092),
.Y(n_7839)
);

CKINVDCx5p33_ASAP7_75t_R g7840 ( 
.A(n_6994),
.Y(n_7840)
);

AND2x2_ASAP7_75t_L g7841 ( 
.A(n_7176),
.B(n_5886),
.Y(n_7841)
);

BUFx6f_ASAP7_75t_L g7842 ( 
.A(n_7093),
.Y(n_7842)
);

AND2x4_ASAP7_75t_L g7843 ( 
.A(n_7381),
.B(n_6071),
.Y(n_7843)
);

BUFx6f_ASAP7_75t_L g7844 ( 
.A(n_7094),
.Y(n_7844)
);

BUFx6f_ASAP7_75t_L g7845 ( 
.A(n_7095),
.Y(n_7845)
);

AND2x2_ASAP7_75t_L g7846 ( 
.A(n_7205),
.B(n_6047),
.Y(n_7846)
);

NAND2xp5_ASAP7_75t_L g7847 ( 
.A(n_7097),
.B(n_6238),
.Y(n_7847)
);

INVx1_ASAP7_75t_L g7848 ( 
.A(n_7098),
.Y(n_7848)
);

INVxp67_ASAP7_75t_L g7849 ( 
.A(n_7413),
.Y(n_7849)
);

BUFx8_ASAP7_75t_SL g7850 ( 
.A(n_7139),
.Y(n_7850)
);

OA21x2_ASAP7_75t_L g7851 ( 
.A1(n_7318),
.A2(n_5225),
.B(n_5220),
.Y(n_7851)
);

INVx1_ASAP7_75t_L g7852 ( 
.A(n_7105),
.Y(n_7852)
);

BUFx12f_ASAP7_75t_L g7853 ( 
.A(n_7399),
.Y(n_7853)
);

CKINVDCx5p33_ASAP7_75t_R g7854 ( 
.A(n_7005),
.Y(n_7854)
);

INVx3_ASAP7_75t_L g7855 ( 
.A(n_7108),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_7106),
.Y(n_7856)
);

AND2x2_ASAP7_75t_L g7857 ( 
.A(n_7209),
.B(n_6047),
.Y(n_7857)
);

INVx1_ASAP7_75t_L g7858 ( 
.A(n_7248),
.Y(n_7858)
);

NOR2xp33_ASAP7_75t_L g7859 ( 
.A(n_7383),
.B(n_7384),
.Y(n_7859)
);

INVx1_ASAP7_75t_L g7860 ( 
.A(n_7250),
.Y(n_7860)
);

BUFx6f_ASAP7_75t_L g7861 ( 
.A(n_7235),
.Y(n_7861)
);

BUFx6f_ASAP7_75t_L g7862 ( 
.A(n_7236),
.Y(n_7862)
);

INVx3_ASAP7_75t_L g7863 ( 
.A(n_7111),
.Y(n_7863)
);

BUFx6f_ASAP7_75t_L g7864 ( 
.A(n_7239),
.Y(n_7864)
);

INVx6_ASAP7_75t_L g7865 ( 
.A(n_7382),
.Y(n_7865)
);

INVx2_ASAP7_75t_L g7866 ( 
.A(n_7240),
.Y(n_7866)
);

NAND2xp5_ASAP7_75t_L g7867 ( 
.A(n_7121),
.B(n_6422),
.Y(n_7867)
);

NOR2x1_ASAP7_75t_L g7868 ( 
.A(n_7387),
.B(n_5178),
.Y(n_7868)
);

INVx2_ASAP7_75t_L g7869 ( 
.A(n_7241),
.Y(n_7869)
);

INVx5_ASAP7_75t_L g7870 ( 
.A(n_6953),
.Y(n_7870)
);

INVx1_ASAP7_75t_L g7871 ( 
.A(n_7252),
.Y(n_7871)
);

INVx2_ASAP7_75t_L g7872 ( 
.A(n_7242),
.Y(n_7872)
);

CKINVDCx5p33_ASAP7_75t_R g7873 ( 
.A(n_7007),
.Y(n_7873)
);

INVx1_ASAP7_75t_L g7874 ( 
.A(n_7253),
.Y(n_7874)
);

BUFx12f_ASAP7_75t_L g7875 ( 
.A(n_7405),
.Y(n_7875)
);

BUFx6f_ASAP7_75t_L g7876 ( 
.A(n_7244),
.Y(n_7876)
);

INVx1_ASAP7_75t_L g7877 ( 
.A(n_7254),
.Y(n_7877)
);

CKINVDCx16_ASAP7_75t_R g7878 ( 
.A(n_7145),
.Y(n_7878)
);

OAI22xp5_ASAP7_75t_SL g7879 ( 
.A1(n_7147),
.A2(n_5658),
.B1(n_5659),
.B2(n_5643),
.Y(n_7879)
);

HB1xp67_ASAP7_75t_L g7880 ( 
.A(n_7006),
.Y(n_7880)
);

AND2x4_ASAP7_75t_L g7881 ( 
.A(n_7389),
.B(n_6449),
.Y(n_7881)
);

INVx2_ASAP7_75t_L g7882 ( 
.A(n_7245),
.Y(n_7882)
);

AND2x2_ASAP7_75t_L g7883 ( 
.A(n_7251),
.B(n_7410),
.Y(n_7883)
);

INVx1_ASAP7_75t_L g7884 ( 
.A(n_7255),
.Y(n_7884)
);

BUFx2_ASAP7_75t_L g7885 ( 
.A(n_7150),
.Y(n_7885)
);

OAI22xp5_ASAP7_75t_L g7886 ( 
.A1(n_7390),
.A2(n_5173),
.B1(n_5179),
.B2(n_5169),
.Y(n_7886)
);

INVx3_ASAP7_75t_L g7887 ( 
.A(n_7256),
.Y(n_7887)
);

BUFx8_ASAP7_75t_SL g7888 ( 
.A(n_7170),
.Y(n_7888)
);

AND2x2_ASAP7_75t_L g7889 ( 
.A(n_7414),
.B(n_6087),
.Y(n_7889)
);

NAND2xp5_ASAP7_75t_L g7890 ( 
.A(n_7123),
.B(n_6460),
.Y(n_7890)
);

AND2x2_ASAP7_75t_L g7891 ( 
.A(n_7416),
.B(n_6087),
.Y(n_7891)
);

HB1xp67_ASAP7_75t_L g7892 ( 
.A(n_7438),
.Y(n_7892)
);

AND2x4_ASAP7_75t_L g7893 ( 
.A(n_7392),
.B(n_5227),
.Y(n_7893)
);

INVx2_ASAP7_75t_L g7894 ( 
.A(n_7259),
.Y(n_7894)
);

NOR2xp33_ASAP7_75t_L g7895 ( 
.A(n_7394),
.B(n_5181),
.Y(n_7895)
);

BUFx6f_ASAP7_75t_L g7896 ( 
.A(n_7261),
.Y(n_7896)
);

OAI22xp5_ASAP7_75t_L g7897 ( 
.A1(n_7396),
.A2(n_5187),
.B1(n_5188),
.B2(n_5182),
.Y(n_7897)
);

INVx3_ASAP7_75t_L g7898 ( 
.A(n_7266),
.Y(n_7898)
);

OAI21x1_ASAP7_75t_L g7899 ( 
.A1(n_7398),
.A2(n_7401),
.B(n_7400),
.Y(n_7899)
);

AND2x2_ASAP7_75t_L g7900 ( 
.A(n_7320),
.B(n_6106),
.Y(n_7900)
);

OAI21x1_ASAP7_75t_L g7901 ( 
.A1(n_7403),
.A2(n_5209),
.B(n_5208),
.Y(n_7901)
);

INVx1_ASAP7_75t_L g7902 ( 
.A(n_7268),
.Y(n_7902)
);

NAND2xp5_ASAP7_75t_SL g7903 ( 
.A(n_7374),
.B(n_5190),
.Y(n_7903)
);

INVx2_ASAP7_75t_L g7904 ( 
.A(n_7321),
.Y(n_7904)
);

NAND2x1p5_ASAP7_75t_L g7905 ( 
.A(n_7409),
.B(n_6105),
.Y(n_7905)
);

INVx2_ASAP7_75t_L g7906 ( 
.A(n_7128),
.Y(n_7906)
);

INVx2_ASAP7_75t_L g7907 ( 
.A(n_7131),
.Y(n_7907)
);

NOR2xp33_ASAP7_75t_L g7908 ( 
.A(n_7411),
.B(n_5191),
.Y(n_7908)
);

NAND2xp5_ASAP7_75t_L g7909 ( 
.A(n_7134),
.B(n_5313),
.Y(n_7909)
);

BUFx6f_ASAP7_75t_L g7910 ( 
.A(n_7418),
.Y(n_7910)
);

CKINVDCx14_ASAP7_75t_R g7911 ( 
.A(n_7173),
.Y(n_7911)
);

INVx4_ASAP7_75t_L g7912 ( 
.A(n_7013),
.Y(n_7912)
);

BUFx6f_ASAP7_75t_L g7913 ( 
.A(n_7412),
.Y(n_7913)
);

BUFx2_ASAP7_75t_L g7914 ( 
.A(n_7179),
.Y(n_7914)
);

AND2x6_ASAP7_75t_L g7915 ( 
.A(n_7311),
.B(n_6115),
.Y(n_7915)
);

HB1xp67_ASAP7_75t_L g7916 ( 
.A(n_7439),
.Y(n_7916)
);

CKINVDCx6p67_ASAP7_75t_R g7917 ( 
.A(n_7001),
.Y(n_7917)
);

INVx1_ASAP7_75t_L g7918 ( 
.A(n_7140),
.Y(n_7918)
);

AND2x4_ASAP7_75t_L g7919 ( 
.A(n_7177),
.B(n_5228),
.Y(n_7919)
);

INVx1_ASAP7_75t_L g7920 ( 
.A(n_7193),
.Y(n_7920)
);

AND2x4_ASAP7_75t_L g7921 ( 
.A(n_7207),
.B(n_5229),
.Y(n_7921)
);

INVx1_ASAP7_75t_L g7922 ( 
.A(n_7212),
.Y(n_7922)
);

INVx1_ASAP7_75t_L g7923 ( 
.A(n_7270),
.Y(n_7923)
);

AND2x4_ASAP7_75t_L g7924 ( 
.A(n_7308),
.B(n_5231),
.Y(n_7924)
);

BUFx12f_ASAP7_75t_L g7925 ( 
.A(n_7407),
.Y(n_7925)
);

NAND2xp5_ASAP7_75t_L g7926 ( 
.A(n_7313),
.B(n_5332),
.Y(n_7926)
);

AND2x2_ASAP7_75t_L g7927 ( 
.A(n_7322),
.B(n_6106),
.Y(n_7927)
);

NAND2xp5_ASAP7_75t_L g7928 ( 
.A(n_7337),
.B(n_5350),
.Y(n_7928)
);

INVx1_ASAP7_75t_L g7929 ( 
.A(n_7324),
.Y(n_7929)
);

INVx3_ASAP7_75t_L g7930 ( 
.A(n_7039),
.Y(n_7930)
);

OA21x2_ASAP7_75t_L g7931 ( 
.A1(n_7041),
.A2(n_5237),
.B(n_5236),
.Y(n_7931)
);

AND2x4_ASAP7_75t_L g7932 ( 
.A(n_7358),
.B(n_5242),
.Y(n_7932)
);

INVx2_ASAP7_75t_L g7933 ( 
.A(n_7404),
.Y(n_7933)
);

AOI22xp5_ASAP7_75t_L g7934 ( 
.A1(n_7052),
.A2(n_6142),
.B1(n_6171),
.B2(n_6120),
.Y(n_7934)
);

INVx6_ASAP7_75t_L g7935 ( 
.A(n_7374),
.Y(n_7935)
);

AND2x4_ASAP7_75t_L g7936 ( 
.A(n_7246),
.B(n_5244),
.Y(n_7936)
);

BUFx12f_ASAP7_75t_L g7937 ( 
.A(n_7053),
.Y(n_7937)
);

INVx1_ASAP7_75t_L g7938 ( 
.A(n_7257),
.Y(n_7938)
);

INVx2_ASAP7_75t_L g7939 ( 
.A(n_7070),
.Y(n_7939)
);

AND2x4_ASAP7_75t_L g7940 ( 
.A(n_7281),
.B(n_5259),
.Y(n_7940)
);

INVx3_ASAP7_75t_L g7941 ( 
.A(n_7112),
.Y(n_7941)
);

CKINVDCx6p67_ASAP7_75t_R g7942 ( 
.A(n_7278),
.Y(n_7942)
);

BUFx6f_ASAP7_75t_L g7943 ( 
.A(n_7148),
.Y(n_7943)
);

BUFx6f_ASAP7_75t_L g7944 ( 
.A(n_7149),
.Y(n_7944)
);

INVx5_ASAP7_75t_L g7945 ( 
.A(n_7045),
.Y(n_7945)
);

INVx1_ASAP7_75t_L g7946 ( 
.A(n_7154),
.Y(n_7946)
);

AND2x2_ASAP7_75t_L g7947 ( 
.A(n_7374),
.B(n_6172),
.Y(n_7947)
);

AND2x2_ASAP7_75t_L g7948 ( 
.A(n_7156),
.B(n_6172),
.Y(n_7948)
);

NAND2xp5_ASAP7_75t_L g7949 ( 
.A(n_7157),
.B(n_5362),
.Y(n_7949)
);

INVx2_ASAP7_75t_L g7950 ( 
.A(n_7158),
.Y(n_7950)
);

INVx1_ASAP7_75t_L g7951 ( 
.A(n_7159),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_7163),
.Y(n_7952)
);

INVx3_ASAP7_75t_L g7953 ( 
.A(n_7174),
.Y(n_7953)
);

AND2x4_ASAP7_75t_L g7954 ( 
.A(n_7182),
.B(n_5275),
.Y(n_7954)
);

INVx2_ASAP7_75t_L g7955 ( 
.A(n_7189),
.Y(n_7955)
);

BUFx6f_ASAP7_75t_L g7956 ( 
.A(n_7195),
.Y(n_7956)
);

AND2x2_ASAP7_75t_L g7957 ( 
.A(n_7197),
.B(n_6211),
.Y(n_7957)
);

INVx1_ASAP7_75t_L g7958 ( 
.A(n_7204),
.Y(n_7958)
);

HB1xp67_ASAP7_75t_L g7959 ( 
.A(n_7208),
.Y(n_7959)
);

BUFx12f_ASAP7_75t_L g7960 ( 
.A(n_7218),
.Y(n_7960)
);

AOI22xp5_ASAP7_75t_L g7961 ( 
.A1(n_7233),
.A2(n_6283),
.B1(n_6354),
.B2(n_6235),
.Y(n_7961)
);

BUFx8_ASAP7_75t_SL g7962 ( 
.A(n_7051),
.Y(n_7962)
);

INVx2_ASAP7_75t_L g7963 ( 
.A(n_7237),
.Y(n_7963)
);

INVx6_ASAP7_75t_L g7964 ( 
.A(n_7119),
.Y(n_7964)
);

INVx3_ASAP7_75t_L g7965 ( 
.A(n_7243),
.Y(n_7965)
);

BUFx2_ASAP7_75t_L g7966 ( 
.A(n_7317),
.Y(n_7966)
);

OAI21x1_ASAP7_75t_L g7967 ( 
.A1(n_7351),
.A2(n_5447),
.B(n_5367),
.Y(n_7967)
);

INVx3_ASAP7_75t_L g7968 ( 
.A(n_7258),
.Y(n_7968)
);

OAI22xp5_ASAP7_75t_L g7969 ( 
.A1(n_7267),
.A2(n_5197),
.B1(n_5199),
.B2(n_5196),
.Y(n_7969)
);

NOR2xp33_ASAP7_75t_L g7970 ( 
.A(n_7269),
.B(n_5200),
.Y(n_7970)
);

CKINVDCx5p33_ASAP7_75t_R g7971 ( 
.A(n_7272),
.Y(n_7971)
);

INVx3_ASAP7_75t_L g7972 ( 
.A(n_7280),
.Y(n_7972)
);

HB1xp67_ASAP7_75t_L g7973 ( 
.A(n_7282),
.Y(n_7973)
);

INVx2_ASAP7_75t_L g7974 ( 
.A(n_7286),
.Y(n_7974)
);

OA21x2_ASAP7_75t_L g7975 ( 
.A1(n_7291),
.A2(n_5281),
.B(n_5280),
.Y(n_7975)
);

NOR2xp33_ASAP7_75t_L g7976 ( 
.A(n_7297),
.B(n_5201),
.Y(n_7976)
);

AND2x6_ASAP7_75t_L g7977 ( 
.A(n_7203),
.B(n_6357),
.Y(n_7977)
);

INVx5_ASAP7_75t_L g7978 ( 
.A(n_7220),
.Y(n_7978)
);

INVx6_ASAP7_75t_L g7979 ( 
.A(n_7072),
.Y(n_7979)
);

INVx1_ASAP7_75t_L g7980 ( 
.A(n_7303),
.Y(n_7980)
);

OA21x2_ASAP7_75t_L g7981 ( 
.A1(n_7306),
.A2(n_5295),
.B(n_5292),
.Y(n_7981)
);

BUFx6f_ASAP7_75t_L g7982 ( 
.A(n_7309),
.Y(n_7982)
);

BUFx3_ASAP7_75t_L g7983 ( 
.A(n_7325),
.Y(n_7983)
);

NOR2xp33_ASAP7_75t_L g7984 ( 
.A(n_7327),
.B(n_5204),
.Y(n_7984)
);

INVx3_ASAP7_75t_L g7985 ( 
.A(n_7330),
.Y(n_7985)
);

NAND2xp5_ASAP7_75t_L g7986 ( 
.A(n_7338),
.B(n_5486),
.Y(n_7986)
);

CKINVDCx5p33_ASAP7_75t_R g7987 ( 
.A(n_7342),
.Y(n_7987)
);

INVx1_ASAP7_75t_L g7988 ( 
.A(n_7350),
.Y(n_7988)
);

AND2x6_ASAP7_75t_L g7989 ( 
.A(n_7435),
.B(n_6361),
.Y(n_7989)
);

INVx2_ASAP7_75t_L g7990 ( 
.A(n_7455),
.Y(n_7990)
);

BUFx6f_ASAP7_75t_L g7991 ( 
.A(n_7457),
.Y(n_7991)
);

BUFx6f_ASAP7_75t_L g7992 ( 
.A(n_7465),
.Y(n_7992)
);

NAND2xp5_ASAP7_75t_L g7993 ( 
.A(n_7335),
.B(n_5495),
.Y(n_7993)
);

INVx3_ASAP7_75t_L g7994 ( 
.A(n_7336),
.Y(n_7994)
);

OAI22xp5_ASAP7_75t_L g7995 ( 
.A1(n_7437),
.A2(n_5205),
.B1(n_5212),
.B2(n_5211),
.Y(n_7995)
);

AND2x4_ASAP7_75t_L g7996 ( 
.A(n_7445),
.B(n_5299),
.Y(n_7996)
);

INVx2_ASAP7_75t_L g7997 ( 
.A(n_7453),
.Y(n_7997)
);

AND2x2_ASAP7_75t_L g7998 ( 
.A(n_7427),
.B(n_6211),
.Y(n_7998)
);

AND2x2_ASAP7_75t_L g7999 ( 
.A(n_7427),
.B(n_6344),
.Y(n_7999)
);

INVx2_ASAP7_75t_L g8000 ( 
.A(n_7081),
.Y(n_8000)
);

AND2x2_ASAP7_75t_L g8001 ( 
.A(n_7427),
.B(n_6344),
.Y(n_8001)
);

BUFx12f_ASAP7_75t_L g8002 ( 
.A(n_7431),
.Y(n_8002)
);

BUFx6f_ASAP7_75t_L g8003 ( 
.A(n_7440),
.Y(n_8003)
);

INVx3_ASAP7_75t_L g8004 ( 
.A(n_7044),
.Y(n_8004)
);

BUFx2_ASAP7_75t_L g8005 ( 
.A(n_7432),
.Y(n_8005)
);

INVx1_ASAP7_75t_L g8006 ( 
.A(n_7117),
.Y(n_8006)
);

AND2x2_ASAP7_75t_L g8007 ( 
.A(n_7427),
.B(n_6456),
.Y(n_8007)
);

INVx1_ASAP7_75t_L g8008 ( 
.A(n_7117),
.Y(n_8008)
);

INVx2_ASAP7_75t_L g8009 ( 
.A(n_7081),
.Y(n_8009)
);

INVx5_ASAP7_75t_L g8010 ( 
.A(n_7422),
.Y(n_8010)
);

BUFx3_ASAP7_75t_L g8011 ( 
.A(n_7434),
.Y(n_8011)
);

BUFx2_ASAP7_75t_L g8012 ( 
.A(n_7432),
.Y(n_8012)
);

INVx1_ASAP7_75t_L g8013 ( 
.A(n_7117),
.Y(n_8013)
);

AOI22xp5_ASAP7_75t_L g8014 ( 
.A1(n_6957),
.A2(n_6413),
.B1(n_6485),
.B2(n_6396),
.Y(n_8014)
);

INVx1_ASAP7_75t_L g8015 ( 
.A(n_7117),
.Y(n_8015)
);

BUFx6f_ASAP7_75t_L g8016 ( 
.A(n_7440),
.Y(n_8016)
);

NAND2xp5_ASAP7_75t_L g8017 ( 
.A(n_7014),
.B(n_5504),
.Y(n_8017)
);

INVx1_ASAP7_75t_L g8018 ( 
.A(n_7117),
.Y(n_8018)
);

INVx2_ASAP7_75t_L g8019 ( 
.A(n_7081),
.Y(n_8019)
);

OA21x2_ASAP7_75t_L g8020 ( 
.A1(n_7277),
.A2(n_5307),
.B(n_5306),
.Y(n_8020)
);

CKINVDCx5p33_ASAP7_75t_R g8021 ( 
.A(n_6949),
.Y(n_8021)
);

INVx1_ASAP7_75t_L g8022 ( 
.A(n_7117),
.Y(n_8022)
);

NOR2xp33_ASAP7_75t_L g8023 ( 
.A(n_7449),
.B(n_5213),
.Y(n_8023)
);

CKINVDCx20_ASAP7_75t_R g8024 ( 
.A(n_6955),
.Y(n_8024)
);

INVx1_ASAP7_75t_L g8025 ( 
.A(n_7117),
.Y(n_8025)
);

INVx2_ASAP7_75t_L g8026 ( 
.A(n_7081),
.Y(n_8026)
);

OA21x2_ASAP7_75t_L g8027 ( 
.A1(n_7277),
.A2(n_5319),
.B(n_5310),
.Y(n_8027)
);

BUFx6f_ASAP7_75t_L g8028 ( 
.A(n_7440),
.Y(n_8028)
);

AOI22xp5_ASAP7_75t_L g8029 ( 
.A1(n_6957),
.A2(n_5217),
.B1(n_5223),
.B2(n_5222),
.Y(n_8029)
);

BUFx12f_ASAP7_75t_L g8030 ( 
.A(n_7431),
.Y(n_8030)
);

BUFx6f_ASAP7_75t_L g8031 ( 
.A(n_7440),
.Y(n_8031)
);

NAND2xp5_ASAP7_75t_L g8032 ( 
.A(n_7014),
.B(n_5507),
.Y(n_8032)
);

INVx1_ASAP7_75t_L g8033 ( 
.A(n_7117),
.Y(n_8033)
);

BUFx3_ASAP7_75t_L g8034 ( 
.A(n_7434),
.Y(n_8034)
);

OAI21x1_ASAP7_75t_L g8035 ( 
.A1(n_7277),
.A2(n_5526),
.B(n_5520),
.Y(n_8035)
);

INVx2_ASAP7_75t_L g8036 ( 
.A(n_7081),
.Y(n_8036)
);

CKINVDCx5p33_ASAP7_75t_R g8037 ( 
.A(n_6949),
.Y(n_8037)
);

BUFx6f_ASAP7_75t_L g8038 ( 
.A(n_7440),
.Y(n_8038)
);

BUFx6f_ASAP7_75t_L g8039 ( 
.A(n_7440),
.Y(n_8039)
);

AOI22xp5_ASAP7_75t_L g8040 ( 
.A1(n_6957),
.A2(n_5226),
.B1(n_5232),
.B2(n_5230),
.Y(n_8040)
);

NAND2xp5_ASAP7_75t_L g8041 ( 
.A(n_7014),
.B(n_5647),
.Y(n_8041)
);

INVx2_ASAP7_75t_L g8042 ( 
.A(n_7081),
.Y(n_8042)
);

INVx2_ASAP7_75t_L g8043 ( 
.A(n_7081),
.Y(n_8043)
);

INVx1_ASAP7_75t_L g8044 ( 
.A(n_7117),
.Y(n_8044)
);

OAI22xp5_ASAP7_75t_SL g8045 ( 
.A1(n_7432),
.A2(n_5692),
.B1(n_5694),
.B2(n_5661),
.Y(n_8045)
);

INVx2_ASAP7_75t_L g8046 ( 
.A(n_7081),
.Y(n_8046)
);

BUFx6f_ASAP7_75t_L g8047 ( 
.A(n_7440),
.Y(n_8047)
);

INVx1_ASAP7_75t_L g8048 ( 
.A(n_7117),
.Y(n_8048)
);

AND2x4_ASAP7_75t_L g8049 ( 
.A(n_7434),
.B(n_5320),
.Y(n_8049)
);

BUFx6f_ASAP7_75t_L g8050 ( 
.A(n_7440),
.Y(n_8050)
);

INVx1_ASAP7_75t_L g8051 ( 
.A(n_7117),
.Y(n_8051)
);

INVx3_ASAP7_75t_L g8052 ( 
.A(n_7044),
.Y(n_8052)
);

NAND2xp5_ASAP7_75t_L g8053 ( 
.A(n_7014),
.B(n_5654),
.Y(n_8053)
);

BUFx6f_ASAP7_75t_L g8054 ( 
.A(n_7440),
.Y(n_8054)
);

NAND2xp5_ASAP7_75t_L g8055 ( 
.A(n_7014),
.B(n_5672),
.Y(n_8055)
);

INVx2_ASAP7_75t_SL g8056 ( 
.A(n_7428),
.Y(n_8056)
);

CKINVDCx5p33_ASAP7_75t_R g8057 ( 
.A(n_7672),
.Y(n_8057)
);

HB1xp67_ASAP7_75t_L g8058 ( 
.A(n_7486),
.Y(n_8058)
);

INVx2_ASAP7_75t_L g8059 ( 
.A(n_7548),
.Y(n_8059)
);

INVx3_ASAP7_75t_L g8060 ( 
.A(n_7534),
.Y(n_8060)
);

INVx1_ASAP7_75t_L g8061 ( 
.A(n_7478),
.Y(n_8061)
);

CKINVDCx5p33_ASAP7_75t_R g8062 ( 
.A(n_7715),
.Y(n_8062)
);

BUFx6f_ASAP7_75t_L g8063 ( 
.A(n_7488),
.Y(n_8063)
);

INVx1_ASAP7_75t_L g8064 ( 
.A(n_7492),
.Y(n_8064)
);

INVx1_ASAP7_75t_L g8065 ( 
.A(n_7500),
.Y(n_8065)
);

CKINVDCx5p33_ASAP7_75t_R g8066 ( 
.A(n_7850),
.Y(n_8066)
);

CKINVDCx5p33_ASAP7_75t_R g8067 ( 
.A(n_7888),
.Y(n_8067)
);

INVx2_ASAP7_75t_L g8068 ( 
.A(n_7519),
.Y(n_8068)
);

INVx1_ASAP7_75t_L g8069 ( 
.A(n_8048),
.Y(n_8069)
);

NAND2xp5_ASAP7_75t_L g8070 ( 
.A(n_8023),
.B(n_7477),
.Y(n_8070)
);

INVx1_ASAP7_75t_L g8071 ( 
.A(n_8051),
.Y(n_8071)
);

INVx2_ASAP7_75t_L g8072 ( 
.A(n_7524),
.Y(n_8072)
);

NOR2xp33_ASAP7_75t_L g8073 ( 
.A(n_7629),
.B(n_5234),
.Y(n_8073)
);

OAI21x1_ASAP7_75t_L g8074 ( 
.A1(n_7563),
.A2(n_5695),
.B(n_5673),
.Y(n_8074)
);

NAND2xp5_ASAP7_75t_SL g8075 ( 
.A(n_7601),
.B(n_5238),
.Y(n_8075)
);

INVx1_ASAP7_75t_L g8076 ( 
.A(n_7509),
.Y(n_8076)
);

INVx1_ASAP7_75t_L g8077 ( 
.A(n_7539),
.Y(n_8077)
);

NAND2xp5_ASAP7_75t_L g8078 ( 
.A(n_7906),
.B(n_5239),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_7545),
.Y(n_8079)
);

INVx1_ASAP7_75t_L g8080 ( 
.A(n_7549),
.Y(n_8080)
);

INVx1_ASAP7_75t_L g8081 ( 
.A(n_8044),
.Y(n_8081)
);

CKINVDCx5p33_ASAP7_75t_R g8082 ( 
.A(n_7962),
.Y(n_8082)
);

CKINVDCx20_ASAP7_75t_R g8083 ( 
.A(n_7586),
.Y(n_8083)
);

INVx1_ASAP7_75t_L g8084 ( 
.A(n_7550),
.Y(n_8084)
);

NAND2xp5_ASAP7_75t_L g8085 ( 
.A(n_7907),
.B(n_5241),
.Y(n_8085)
);

CKINVDCx20_ASAP7_75t_R g8086 ( 
.A(n_8024),
.Y(n_8086)
);

INVx1_ASAP7_75t_L g8087 ( 
.A(n_7556),
.Y(n_8087)
);

NOR2xp33_ASAP7_75t_L g8088 ( 
.A(n_7476),
.B(n_7949),
.Y(n_8088)
);

CKINVDCx5p33_ASAP7_75t_R g8089 ( 
.A(n_7508),
.Y(n_8089)
);

INVx1_ASAP7_75t_L g8090 ( 
.A(n_7561),
.Y(n_8090)
);

INVxp67_ASAP7_75t_L g8091 ( 
.A(n_7536),
.Y(n_8091)
);

CKINVDCx5p33_ASAP7_75t_R g8092 ( 
.A(n_7547),
.Y(n_8092)
);

INVx2_ASAP7_75t_L g8093 ( 
.A(n_7527),
.Y(n_8093)
);

AND2x4_ASAP7_75t_L g8094 ( 
.A(n_7483),
.B(n_5325),
.Y(n_8094)
);

INVx1_ASAP7_75t_L g8095 ( 
.A(n_7562),
.Y(n_8095)
);

CKINVDCx5p33_ASAP7_75t_R g8096 ( 
.A(n_7569),
.Y(n_8096)
);

NAND2xp5_ASAP7_75t_L g8097 ( 
.A(n_7816),
.B(n_5245),
.Y(n_8097)
);

CKINVDCx5p33_ASAP7_75t_R g8098 ( 
.A(n_7693),
.Y(n_8098)
);

CKINVDCx5p33_ASAP7_75t_R g8099 ( 
.A(n_7760),
.Y(n_8099)
);

INVx1_ASAP7_75t_L g8100 ( 
.A(n_7578),
.Y(n_8100)
);

INVx1_ASAP7_75t_L g8101 ( 
.A(n_7583),
.Y(n_8101)
);

CKINVDCx5p33_ASAP7_75t_R g8102 ( 
.A(n_7819),
.Y(n_8102)
);

INVx1_ASAP7_75t_L g8103 ( 
.A(n_7593),
.Y(n_8103)
);

NAND2xp5_ASAP7_75t_SL g8104 ( 
.A(n_8056),
.B(n_5246),
.Y(n_8104)
);

NAND2xp5_ASAP7_75t_L g8105 ( 
.A(n_7818),
.B(n_5247),
.Y(n_8105)
);

NAND2xp33_ASAP7_75t_L g8106 ( 
.A(n_7507),
.B(n_5248),
.Y(n_8106)
);

CKINVDCx5p33_ASAP7_75t_R g8107 ( 
.A(n_7832),
.Y(n_8107)
);

AND2x4_ASAP7_75t_L g8108 ( 
.A(n_8011),
.B(n_5337),
.Y(n_8108)
);

INVx2_ASAP7_75t_L g8109 ( 
.A(n_7537),
.Y(n_8109)
);

NOR2xp33_ASAP7_75t_L g8110 ( 
.A(n_7986),
.B(n_5249),
.Y(n_8110)
);

INVx2_ASAP7_75t_L g8111 ( 
.A(n_7538),
.Y(n_8111)
);

INVx1_ASAP7_75t_L g8112 ( 
.A(n_7609),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_7614),
.Y(n_8113)
);

INVx2_ASAP7_75t_L g8114 ( 
.A(n_7576),
.Y(n_8114)
);

BUFx6f_ASAP7_75t_L g8115 ( 
.A(n_7490),
.Y(n_8115)
);

INVx2_ASAP7_75t_L g8116 ( 
.A(n_7577),
.Y(n_8116)
);

INVx1_ASAP7_75t_L g8117 ( 
.A(n_7616),
.Y(n_8117)
);

CKINVDCx5p33_ASAP7_75t_R g8118 ( 
.A(n_7840),
.Y(n_8118)
);

INVx2_ASAP7_75t_L g8119 ( 
.A(n_7810),
.Y(n_8119)
);

INVx1_ASAP7_75t_L g8120 ( 
.A(n_7617),
.Y(n_8120)
);

CKINVDCx5p33_ASAP7_75t_R g8121 ( 
.A(n_7854),
.Y(n_8121)
);

INVx1_ASAP7_75t_L g8122 ( 
.A(n_7632),
.Y(n_8122)
);

INVx1_ASAP7_75t_L g8123 ( 
.A(n_7638),
.Y(n_8123)
);

AND2x2_ASAP7_75t_L g8124 ( 
.A(n_7520),
.B(n_5731),
.Y(n_8124)
);

CKINVDCx5p33_ASAP7_75t_R g8125 ( 
.A(n_7873),
.Y(n_8125)
);

INVx2_ASAP7_75t_L g8126 ( 
.A(n_7815),
.Y(n_8126)
);

INVx2_ASAP7_75t_L g8127 ( 
.A(n_7820),
.Y(n_8127)
);

CKINVDCx20_ASAP7_75t_R g8128 ( 
.A(n_7648),
.Y(n_8128)
);

CKINVDCx5p33_ASAP7_75t_R g8129 ( 
.A(n_7971),
.Y(n_8129)
);

CKINVDCx20_ASAP7_75t_R g8130 ( 
.A(n_7878),
.Y(n_8130)
);

INVx1_ASAP7_75t_L g8131 ( 
.A(n_7651),
.Y(n_8131)
);

CKINVDCx5p33_ASAP7_75t_R g8132 ( 
.A(n_7987),
.Y(n_8132)
);

CKINVDCx5p33_ASAP7_75t_R g8133 ( 
.A(n_8021),
.Y(n_8133)
);

INVx2_ASAP7_75t_L g8134 ( 
.A(n_7821),
.Y(n_8134)
);

AND2x2_ASAP7_75t_L g8135 ( 
.A(n_7501),
.B(n_5732),
.Y(n_8135)
);

CKINVDCx5p33_ASAP7_75t_R g8136 ( 
.A(n_8037),
.Y(n_8136)
);

INVx2_ASAP7_75t_L g8137 ( 
.A(n_7823),
.Y(n_8137)
);

INVx1_ASAP7_75t_L g8138 ( 
.A(n_7654),
.Y(n_8138)
);

CKINVDCx5p33_ASAP7_75t_R g8139 ( 
.A(n_7691),
.Y(n_8139)
);

AND2x2_ASAP7_75t_L g8140 ( 
.A(n_7485),
.B(n_7541),
.Y(n_8140)
);

CKINVDCx5p33_ASAP7_75t_R g8141 ( 
.A(n_7685),
.Y(n_8141)
);

INVx1_ASAP7_75t_L g8142 ( 
.A(n_7655),
.Y(n_8142)
);

INVx1_ASAP7_75t_L g8143 ( 
.A(n_7658),
.Y(n_8143)
);

INVx1_ASAP7_75t_L g8144 ( 
.A(n_7670),
.Y(n_8144)
);

CKINVDCx5p33_ASAP7_75t_R g8145 ( 
.A(n_7790),
.Y(n_8145)
);

CKINVDCx5p33_ASAP7_75t_R g8146 ( 
.A(n_7853),
.Y(n_8146)
);

INVxp67_ASAP7_75t_L g8147 ( 
.A(n_7883),
.Y(n_8147)
);

INVx2_ASAP7_75t_L g8148 ( 
.A(n_7525),
.Y(n_8148)
);

INVx1_ASAP7_75t_L g8149 ( 
.A(n_7676),
.Y(n_8149)
);

INVx1_ASAP7_75t_L g8150 ( 
.A(n_7679),
.Y(n_8150)
);

AND2x2_ASAP7_75t_L g8151 ( 
.A(n_7479),
.B(n_5739),
.Y(n_8151)
);

CKINVDCx5p33_ASAP7_75t_R g8152 ( 
.A(n_7875),
.Y(n_8152)
);

INVx1_ASAP7_75t_L g8153 ( 
.A(n_7681),
.Y(n_8153)
);

NOR2xp33_ASAP7_75t_R g8154 ( 
.A(n_7911),
.B(n_5758),
.Y(n_8154)
);

NAND2xp33_ASAP7_75t_R g8155 ( 
.A(n_7473),
.B(n_5250),
.Y(n_8155)
);

INVx1_ASAP7_75t_L g8156 ( 
.A(n_7684),
.Y(n_8156)
);

INVx6_ASAP7_75t_L g8157 ( 
.A(n_7600),
.Y(n_8157)
);

NAND2xp5_ASAP7_75t_L g8158 ( 
.A(n_7837),
.B(n_5253),
.Y(n_8158)
);

CKINVDCx20_ASAP7_75t_R g8159 ( 
.A(n_7942),
.Y(n_8159)
);

OA21x2_ASAP7_75t_L g8160 ( 
.A1(n_7899),
.A2(n_5341),
.B(n_5340),
.Y(n_8160)
);

NAND2xp5_ASAP7_75t_L g8161 ( 
.A(n_7839),
.B(n_5254),
.Y(n_8161)
);

CKINVDCx5p33_ASAP7_75t_R g8162 ( 
.A(n_7925),
.Y(n_8162)
);

INVx2_ASAP7_75t_L g8163 ( 
.A(n_7526),
.Y(n_8163)
);

CKINVDCx5p33_ASAP7_75t_R g8164 ( 
.A(n_7937),
.Y(n_8164)
);

INVx2_ASAP7_75t_L g8165 ( 
.A(n_7535),
.Y(n_8165)
);

INVx1_ASAP7_75t_L g8166 ( 
.A(n_7696),
.Y(n_8166)
);

HB1xp67_ASAP7_75t_L g8167 ( 
.A(n_7798),
.Y(n_8167)
);

NAND2xp5_ASAP7_75t_L g8168 ( 
.A(n_7848),
.B(n_5255),
.Y(n_8168)
);

BUFx2_ASAP7_75t_L g8169 ( 
.A(n_7799),
.Y(n_8169)
);

NOR2xp33_ASAP7_75t_R g8170 ( 
.A(n_8002),
.B(n_5834),
.Y(n_8170)
);

INVx1_ASAP7_75t_L g8171 ( 
.A(n_7704),
.Y(n_8171)
);

CKINVDCx5p33_ASAP7_75t_R g8172 ( 
.A(n_7960),
.Y(n_8172)
);

AND2x6_ASAP7_75t_L g8173 ( 
.A(n_7947),
.B(n_5343),
.Y(n_8173)
);

NOR2xp33_ASAP7_75t_L g8174 ( 
.A(n_7970),
.B(n_5257),
.Y(n_8174)
);

NAND2xp5_ASAP7_75t_L g8175 ( 
.A(n_7852),
.B(n_5261),
.Y(n_8175)
);

CKINVDCx20_ASAP7_75t_R g8176 ( 
.A(n_7917),
.Y(n_8176)
);

INVx3_ASAP7_75t_L g8177 ( 
.A(n_7499),
.Y(n_8177)
);

AND2x2_ASAP7_75t_L g8178 ( 
.A(n_7998),
.B(n_5838),
.Y(n_8178)
);

CKINVDCx5p33_ASAP7_75t_R g8179 ( 
.A(n_8030),
.Y(n_8179)
);

INVx1_ASAP7_75t_L g8180 ( 
.A(n_7708),
.Y(n_8180)
);

INVx1_ASAP7_75t_L g8181 ( 
.A(n_7713),
.Y(n_8181)
);

INVx1_ASAP7_75t_L g8182 ( 
.A(n_7737),
.Y(n_8182)
);

BUFx6f_ASAP7_75t_L g8183 ( 
.A(n_7502),
.Y(n_8183)
);

INVx2_ASAP7_75t_L g8184 ( 
.A(n_7540),
.Y(n_8184)
);

CKINVDCx20_ASAP7_75t_R g8185 ( 
.A(n_7731),
.Y(n_8185)
);

CKINVDCx5p33_ASAP7_75t_R g8186 ( 
.A(n_7564),
.Y(n_8186)
);

INVx1_ASAP7_75t_L g8187 ( 
.A(n_7742),
.Y(n_8187)
);

CKINVDCx20_ASAP7_75t_R g8188 ( 
.A(n_7768),
.Y(n_8188)
);

CKINVDCx20_ASAP7_75t_R g8189 ( 
.A(n_7641),
.Y(n_8189)
);

CKINVDCx20_ASAP7_75t_R g8190 ( 
.A(n_7807),
.Y(n_8190)
);

INVx3_ASAP7_75t_L g8191 ( 
.A(n_7503),
.Y(n_8191)
);

OA21x2_ASAP7_75t_L g8192 ( 
.A1(n_7574),
.A2(n_5357),
.B(n_5348),
.Y(n_8192)
);

CKINVDCx20_ASAP7_75t_R g8193 ( 
.A(n_7885),
.Y(n_8193)
);

AND2x2_ASAP7_75t_L g8194 ( 
.A(n_7999),
.B(n_5839),
.Y(n_8194)
);

INVx1_ASAP7_75t_L g8195 ( 
.A(n_7749),
.Y(n_8195)
);

INVx1_ASAP7_75t_L g8196 ( 
.A(n_7750),
.Y(n_8196)
);

AND2x2_ASAP7_75t_L g8197 ( 
.A(n_8001),
.B(n_5847),
.Y(n_8197)
);

CKINVDCx5p33_ASAP7_75t_R g8198 ( 
.A(n_7943),
.Y(n_8198)
);

INVx1_ASAP7_75t_L g8199 ( 
.A(n_7752),
.Y(n_8199)
);

AND2x4_ASAP7_75t_L g8200 ( 
.A(n_8034),
.B(n_5369),
.Y(n_8200)
);

INVx1_ASAP7_75t_L g8201 ( 
.A(n_7763),
.Y(n_8201)
);

NAND2xp5_ASAP7_75t_L g8202 ( 
.A(n_7856),
.B(n_5263),
.Y(n_8202)
);

CKINVDCx5p33_ASAP7_75t_R g8203 ( 
.A(n_7944),
.Y(n_8203)
);

INVx1_ASAP7_75t_L g8204 ( 
.A(n_7766),
.Y(n_8204)
);

HB1xp67_ASAP7_75t_L g8205 ( 
.A(n_7827),
.Y(n_8205)
);

INVx1_ASAP7_75t_L g8206 ( 
.A(n_7772),
.Y(n_8206)
);

INVx3_ASAP7_75t_L g8207 ( 
.A(n_7506),
.Y(n_8207)
);

AND2x2_ASAP7_75t_L g8208 ( 
.A(n_8007),
.B(n_5852),
.Y(n_8208)
);

CKINVDCx5p33_ASAP7_75t_R g8209 ( 
.A(n_7956),
.Y(n_8209)
);

CKINVDCx5p33_ASAP7_75t_R g8210 ( 
.A(n_7982),
.Y(n_8210)
);

NOR2xp33_ASAP7_75t_L g8211 ( 
.A(n_7976),
.B(n_5265),
.Y(n_8211)
);

INVx1_ASAP7_75t_L g8212 ( 
.A(n_7783),
.Y(n_8212)
);

AND2x6_ASAP7_75t_L g8213 ( 
.A(n_7755),
.B(n_5370),
.Y(n_8213)
);

NOR2xp33_ASAP7_75t_R g8214 ( 
.A(n_7994),
.B(n_5870),
.Y(n_8214)
);

INVx1_ASAP7_75t_L g8215 ( 
.A(n_7785),
.Y(n_8215)
);

INVx3_ASAP7_75t_L g8216 ( 
.A(n_8003),
.Y(n_8216)
);

CKINVDCx5p33_ASAP7_75t_R g8217 ( 
.A(n_7991),
.Y(n_8217)
);

NAND2xp5_ASAP7_75t_L g8218 ( 
.A(n_7918),
.B(n_5266),
.Y(n_8218)
);

INVx1_ASAP7_75t_L g8219 ( 
.A(n_7804),
.Y(n_8219)
);

INVx1_ASAP7_75t_L g8220 ( 
.A(n_7808),
.Y(n_8220)
);

INVx2_ASAP7_75t_L g8221 ( 
.A(n_7829),
.Y(n_8221)
);

CKINVDCx5p33_ASAP7_75t_R g8222 ( 
.A(n_7992),
.Y(n_8222)
);

CKINVDCx20_ASAP7_75t_R g8223 ( 
.A(n_7914),
.Y(n_8223)
);

INVx1_ASAP7_75t_L g8224 ( 
.A(n_8006),
.Y(n_8224)
);

BUFx6f_ASAP7_75t_L g8225 ( 
.A(n_8016),
.Y(n_8225)
);

INVx1_ASAP7_75t_L g8226 ( 
.A(n_8008),
.Y(n_8226)
);

INVx2_ASAP7_75t_L g8227 ( 
.A(n_7866),
.Y(n_8227)
);

CKINVDCx20_ASAP7_75t_R g8228 ( 
.A(n_7650),
.Y(n_8228)
);

OR2x2_ASAP7_75t_L g8229 ( 
.A(n_7880),
.B(n_7892),
.Y(n_8229)
);

CKINVDCx5p33_ASAP7_75t_R g8230 ( 
.A(n_7665),
.Y(n_8230)
);

BUFx8_ASAP7_75t_L g8231 ( 
.A(n_8005),
.Y(n_8231)
);

BUFx2_ASAP7_75t_L g8232 ( 
.A(n_7916),
.Y(n_8232)
);

CKINVDCx5p33_ASAP7_75t_R g8233 ( 
.A(n_7979),
.Y(n_8233)
);

INVx2_ASAP7_75t_L g8234 ( 
.A(n_7869),
.Y(n_8234)
);

HB1xp67_ASAP7_75t_L g8235 ( 
.A(n_7528),
.Y(n_8235)
);

BUFx6f_ASAP7_75t_L g8236 ( 
.A(n_8028),
.Y(n_8236)
);

INVx2_ASAP7_75t_L g8237 ( 
.A(n_7872),
.Y(n_8237)
);

CKINVDCx5p33_ASAP7_75t_R g8238 ( 
.A(n_7673),
.Y(n_8238)
);

NAND2xp5_ASAP7_75t_SL g8239 ( 
.A(n_7825),
.B(n_5268),
.Y(n_8239)
);

BUFx6f_ASAP7_75t_L g8240 ( 
.A(n_8031),
.Y(n_8240)
);

AND2x2_ASAP7_75t_L g8241 ( 
.A(n_7546),
.B(n_7589),
.Y(n_8241)
);

HB1xp67_ASAP7_75t_L g8242 ( 
.A(n_8012),
.Y(n_8242)
);

INVx2_ASAP7_75t_L g8243 ( 
.A(n_7882),
.Y(n_8243)
);

AND2x4_ASAP7_75t_L g8244 ( 
.A(n_7513),
.B(n_5379),
.Y(n_8244)
);

INVx1_ASAP7_75t_L g8245 ( 
.A(n_8013),
.Y(n_8245)
);

NOR2xp33_ASAP7_75t_L g8246 ( 
.A(n_7984),
.B(n_5270),
.Y(n_8246)
);

CKINVDCx20_ASAP7_75t_R g8247 ( 
.A(n_7727),
.Y(n_8247)
);

INVx2_ASAP7_75t_L g8248 ( 
.A(n_7553),
.Y(n_8248)
);

NAND2xp5_ASAP7_75t_L g8249 ( 
.A(n_7920),
.B(n_5274),
.Y(n_8249)
);

CKINVDCx5p33_ASAP7_75t_R g8250 ( 
.A(n_7740),
.Y(n_8250)
);

CKINVDCx5p33_ASAP7_75t_R g8251 ( 
.A(n_7817),
.Y(n_8251)
);

CKINVDCx20_ASAP7_75t_R g8252 ( 
.A(n_7824),
.Y(n_8252)
);

AND2x2_ASAP7_75t_L g8253 ( 
.A(n_7592),
.B(n_5910),
.Y(n_8253)
);

CKINVDCx5p33_ASAP7_75t_R g8254 ( 
.A(n_7834),
.Y(n_8254)
);

INVx3_ASAP7_75t_L g8255 ( 
.A(n_8038),
.Y(n_8255)
);

INVx1_ASAP7_75t_L g8256 ( 
.A(n_8015),
.Y(n_8256)
);

CKINVDCx5p33_ASAP7_75t_R g8257 ( 
.A(n_7983),
.Y(n_8257)
);

AND2x4_ASAP7_75t_L g8258 ( 
.A(n_7495),
.B(n_5386),
.Y(n_8258)
);

INVx2_ASAP7_75t_L g8259 ( 
.A(n_7554),
.Y(n_8259)
);

CKINVDCx20_ASAP7_75t_R g8260 ( 
.A(n_7714),
.Y(n_8260)
);

CKINVDCx5p33_ASAP7_75t_R g8261 ( 
.A(n_7661),
.Y(n_8261)
);

INVx1_ASAP7_75t_L g8262 ( 
.A(n_8018),
.Y(n_8262)
);

INVx3_ASAP7_75t_L g8263 ( 
.A(n_8039),
.Y(n_8263)
);

INVx1_ASAP7_75t_L g8264 ( 
.A(n_8022),
.Y(n_8264)
);

HB1xp67_ASAP7_75t_L g8265 ( 
.A(n_7996),
.Y(n_8265)
);

INVx2_ASAP7_75t_L g8266 ( 
.A(n_7565),
.Y(n_8266)
);

CKINVDCx5p33_ASAP7_75t_R g8267 ( 
.A(n_7912),
.Y(n_8267)
);

CKINVDCx5p33_ASAP7_75t_R g8268 ( 
.A(n_7930),
.Y(n_8268)
);

NOR2xp33_ASAP7_75t_L g8269 ( 
.A(n_7579),
.B(n_5276),
.Y(n_8269)
);

INVx4_ASAP7_75t_L g8270 ( 
.A(n_7643),
.Y(n_8270)
);

INVx2_ASAP7_75t_L g8271 ( 
.A(n_7567),
.Y(n_8271)
);

CKINVDCx5p33_ASAP7_75t_R g8272 ( 
.A(n_7941),
.Y(n_8272)
);

INVx1_ASAP7_75t_L g8273 ( 
.A(n_8025),
.Y(n_8273)
);

INVxp67_ASAP7_75t_SL g8274 ( 
.A(n_7732),
.Y(n_8274)
);

CKINVDCx5p33_ASAP7_75t_R g8275 ( 
.A(n_7953),
.Y(n_8275)
);

XOR2xp5_ASAP7_75t_L g8276 ( 
.A(n_7718),
.B(n_5925),
.Y(n_8276)
);

AND2x2_ASAP7_75t_L g8277 ( 
.A(n_7596),
.B(n_7687),
.Y(n_8277)
);

INVx1_ASAP7_75t_L g8278 ( 
.A(n_8033),
.Y(n_8278)
);

INVx1_ASAP7_75t_L g8279 ( 
.A(n_7736),
.Y(n_8279)
);

AND2x2_ASAP7_75t_L g8280 ( 
.A(n_7900),
.B(n_5930),
.Y(n_8280)
);

NAND2xp5_ASAP7_75t_L g8281 ( 
.A(n_7922),
.B(n_5277),
.Y(n_8281)
);

INVxp67_ASAP7_75t_L g8282 ( 
.A(n_7789),
.Y(n_8282)
);

OAI22xp5_ASAP7_75t_L g8283 ( 
.A1(n_7859),
.A2(n_7923),
.B1(n_8032),
.B2(n_8017),
.Y(n_8283)
);

CKINVDCx5p33_ASAP7_75t_R g8284 ( 
.A(n_7965),
.Y(n_8284)
);

INVx1_ASAP7_75t_L g8285 ( 
.A(n_7858),
.Y(n_8285)
);

CKINVDCx5p33_ASAP7_75t_R g8286 ( 
.A(n_7968),
.Y(n_8286)
);

CKINVDCx5p33_ASAP7_75t_R g8287 ( 
.A(n_7972),
.Y(n_8287)
);

NAND2xp5_ASAP7_75t_L g8288 ( 
.A(n_8041),
.B(n_5278),
.Y(n_8288)
);

CKINVDCx20_ASAP7_75t_R g8289 ( 
.A(n_7739),
.Y(n_8289)
);

CKINVDCx5p33_ASAP7_75t_R g8290 ( 
.A(n_7985),
.Y(n_8290)
);

BUFx2_ASAP7_75t_L g8291 ( 
.A(n_7507),
.Y(n_8291)
);

NOR2xp67_ASAP7_75t_L g8292 ( 
.A(n_7870),
.B(n_4325),
.Y(n_8292)
);

NAND2xp5_ASAP7_75t_SL g8293 ( 
.A(n_7619),
.B(n_5282),
.Y(n_8293)
);

INVx1_ASAP7_75t_L g8294 ( 
.A(n_7860),
.Y(n_8294)
);

INVxp67_ASAP7_75t_L g8295 ( 
.A(n_7841),
.Y(n_8295)
);

BUFx10_ASAP7_75t_L g8296 ( 
.A(n_7964),
.Y(n_8296)
);

INVx3_ASAP7_75t_L g8297 ( 
.A(n_8047),
.Y(n_8297)
);

CKINVDCx5p33_ASAP7_75t_R g8298 ( 
.A(n_7830),
.Y(n_8298)
);

INVx1_ASAP7_75t_L g8299 ( 
.A(n_7871),
.Y(n_8299)
);

AND2x4_ASAP7_75t_L g8300 ( 
.A(n_7504),
.B(n_5396),
.Y(n_8300)
);

INVx1_ASAP7_75t_L g8301 ( 
.A(n_7874),
.Y(n_8301)
);

INVx1_ASAP7_75t_L g8302 ( 
.A(n_7877),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_7884),
.Y(n_8303)
);

INVx1_ASAP7_75t_L g8304 ( 
.A(n_7902),
.Y(n_8304)
);

CKINVDCx20_ASAP7_75t_R g8305 ( 
.A(n_7966),
.Y(n_8305)
);

NAND2xp5_ASAP7_75t_L g8306 ( 
.A(n_8053),
.B(n_8055),
.Y(n_8306)
);

CKINVDCx5p33_ASAP7_75t_R g8307 ( 
.A(n_7588),
.Y(n_8307)
);

INVx1_ASAP7_75t_L g8308 ( 
.A(n_8020),
.Y(n_8308)
);

INVx1_ASAP7_75t_L g8309 ( 
.A(n_8027),
.Y(n_8309)
);

INVx1_ASAP7_75t_L g8310 ( 
.A(n_7759),
.Y(n_8310)
);

AND2x4_ASAP7_75t_L g8311 ( 
.A(n_8004),
.B(n_5397),
.Y(n_8311)
);

BUFx6f_ASAP7_75t_L g8312 ( 
.A(n_8050),
.Y(n_8312)
);

INVx1_ASAP7_75t_L g8313 ( 
.A(n_7774),
.Y(n_8313)
);

CKINVDCx5p33_ASAP7_75t_R g8314 ( 
.A(n_7959),
.Y(n_8314)
);

CKINVDCx5p33_ASAP7_75t_R g8315 ( 
.A(n_7973),
.Y(n_8315)
);

NAND2xp5_ASAP7_75t_SL g8316 ( 
.A(n_7913),
.B(n_5283),
.Y(n_8316)
);

CKINVDCx5p33_ASAP7_75t_R g8317 ( 
.A(n_7754),
.Y(n_8317)
);

AND2x2_ASAP7_75t_L g8318 ( 
.A(n_7846),
.B(n_5934),
.Y(n_8318)
);

BUFx10_ASAP7_75t_L g8319 ( 
.A(n_7532),
.Y(n_8319)
);

BUFx2_ASAP7_75t_L g8320 ( 
.A(n_7610),
.Y(n_8320)
);

INVx1_ASAP7_75t_L g8321 ( 
.A(n_7776),
.Y(n_8321)
);

NOR2xp67_ASAP7_75t_L g8322 ( 
.A(n_7945),
.B(n_4326),
.Y(n_8322)
);

CKINVDCx5p33_ASAP7_75t_R g8323 ( 
.A(n_7978),
.Y(n_8323)
);

NOR2xp67_ASAP7_75t_L g8324 ( 
.A(n_7764),
.B(n_4328),
.Y(n_8324)
);

INVx1_ASAP7_75t_L g8325 ( 
.A(n_7784),
.Y(n_8325)
);

INVx2_ASAP7_75t_L g8326 ( 
.A(n_7571),
.Y(n_8326)
);

NAND2xp5_ASAP7_75t_L g8327 ( 
.A(n_7904),
.B(n_5284),
.Y(n_8327)
);

CKINVDCx5p33_ASAP7_75t_R g8328 ( 
.A(n_7865),
.Y(n_8328)
);

NAND2xp33_ASAP7_75t_SL g8329 ( 
.A(n_7948),
.B(n_7957),
.Y(n_8329)
);

CKINVDCx5p33_ASAP7_75t_R g8330 ( 
.A(n_7611),
.Y(n_8330)
);

CKINVDCx20_ASAP7_75t_R g8331 ( 
.A(n_7628),
.Y(n_8331)
);

AND2x4_ASAP7_75t_L g8332 ( 
.A(n_8052),
.B(n_7518),
.Y(n_8332)
);

INVx2_ASAP7_75t_L g8333 ( 
.A(n_7575),
.Y(n_8333)
);

NOR2xp67_ASAP7_75t_L g8334 ( 
.A(n_7765),
.B(n_4329),
.Y(n_8334)
);

INVxp33_ASAP7_75t_SL g8335 ( 
.A(n_7726),
.Y(n_8335)
);

NOR2xp33_ASAP7_75t_L g8336 ( 
.A(n_7926),
.B(n_5285),
.Y(n_8336)
);

INVx2_ASAP7_75t_L g8337 ( 
.A(n_7786),
.Y(n_8337)
);

INVx1_ASAP7_75t_L g8338 ( 
.A(n_7795),
.Y(n_8338)
);

INVx2_ASAP7_75t_L g8339 ( 
.A(n_7796),
.Y(n_8339)
);

NOR2xp33_ASAP7_75t_L g8340 ( 
.A(n_7928),
.B(n_5288),
.Y(n_8340)
);

CKINVDCx5p33_ASAP7_75t_R g8341 ( 
.A(n_7612),
.Y(n_8341)
);

INVx1_ASAP7_75t_L g8342 ( 
.A(n_7788),
.Y(n_8342)
);

AND2x2_ASAP7_75t_L g8343 ( 
.A(n_7857),
.B(n_5944),
.Y(n_8343)
);

BUFx6f_ASAP7_75t_L g8344 ( 
.A(n_8054),
.Y(n_8344)
);

BUFx6f_ASAP7_75t_L g8345 ( 
.A(n_7517),
.Y(n_8345)
);

AND2x6_ASAP7_75t_L g8346 ( 
.A(n_7787),
.B(n_5402),
.Y(n_8346)
);

BUFx3_ASAP7_75t_L g8347 ( 
.A(n_7522),
.Y(n_8347)
);

AND2x2_ASAP7_75t_L g8348 ( 
.A(n_7889),
.B(n_5972),
.Y(n_8348)
);

INVx2_ASAP7_75t_L g8349 ( 
.A(n_7581),
.Y(n_8349)
);

CKINVDCx5p33_ASAP7_75t_R g8350 ( 
.A(n_7555),
.Y(n_8350)
);

BUFx3_ASAP7_75t_L g8351 ( 
.A(n_7523),
.Y(n_8351)
);

CKINVDCx5p33_ASAP7_75t_R g8352 ( 
.A(n_7728),
.Y(n_8352)
);

INVx2_ASAP7_75t_L g8353 ( 
.A(n_7590),
.Y(n_8353)
);

INVx2_ASAP7_75t_L g8354 ( 
.A(n_7594),
.Y(n_8354)
);

INVx1_ASAP7_75t_L g8355 ( 
.A(n_7894),
.Y(n_8355)
);

INVx1_ASAP7_75t_L g8356 ( 
.A(n_7595),
.Y(n_8356)
);

NOR2x1_ASAP7_75t_L g8357 ( 
.A(n_7993),
.B(n_5202),
.Y(n_8357)
);

CKINVDCx5p33_ASAP7_75t_R g8358 ( 
.A(n_7680),
.Y(n_8358)
);

INVx1_ASAP7_75t_L g8359 ( 
.A(n_7598),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_7607),
.Y(n_8360)
);

INVx2_ASAP7_75t_L g8361 ( 
.A(n_7618),
.Y(n_8361)
);

INVx1_ASAP7_75t_L g8362 ( 
.A(n_7624),
.Y(n_8362)
);

NAND2xp5_ASAP7_75t_L g8363 ( 
.A(n_7698),
.B(n_5291),
.Y(n_8363)
);

INVx1_ASAP7_75t_L g8364 ( 
.A(n_7627),
.Y(n_8364)
);

CKINVDCx5p33_ASAP7_75t_R g8365 ( 
.A(n_7939),
.Y(n_8365)
);

AND2x2_ASAP7_75t_L g8366 ( 
.A(n_7891),
.B(n_6009),
.Y(n_8366)
);

INVx2_ASAP7_75t_L g8367 ( 
.A(n_7636),
.Y(n_8367)
);

CKINVDCx5p33_ASAP7_75t_R g8368 ( 
.A(n_7950),
.Y(n_8368)
);

NAND2xp5_ASAP7_75t_L g8369 ( 
.A(n_7730),
.B(n_5293),
.Y(n_8369)
);

INVx1_ASAP7_75t_L g8370 ( 
.A(n_7644),
.Y(n_8370)
);

CKINVDCx20_ASAP7_75t_R g8371 ( 
.A(n_7558),
.Y(n_8371)
);

CKINVDCx20_ASAP7_75t_R g8372 ( 
.A(n_7879),
.Y(n_8372)
);

INVx1_ASAP7_75t_L g8373 ( 
.A(n_7645),
.Y(n_8373)
);

INVx1_ASAP7_75t_L g8374 ( 
.A(n_7647),
.Y(n_8374)
);

NAND2xp5_ASAP7_75t_SL g8375 ( 
.A(n_7689),
.B(n_5294),
.Y(n_8375)
);

INVx1_ASAP7_75t_L g8376 ( 
.A(n_7653),
.Y(n_8376)
);

INVx2_ASAP7_75t_L g8377 ( 
.A(n_7657),
.Y(n_8377)
);

INVx1_ASAP7_75t_L g8378 ( 
.A(n_7695),
.Y(n_8378)
);

INVx1_ASAP7_75t_L g8379 ( 
.A(n_7701),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7703),
.Y(n_8380)
);

INVx2_ASAP7_75t_L g8381 ( 
.A(n_7705),
.Y(n_8381)
);

INVx3_ASAP7_75t_L g8382 ( 
.A(n_7861),
.Y(n_8382)
);

NOR2xp33_ASAP7_75t_L g8383 ( 
.A(n_7484),
.B(n_5296),
.Y(n_8383)
);

INVx2_ASAP7_75t_L g8384 ( 
.A(n_7717),
.Y(n_8384)
);

NAND2xp33_ASAP7_75t_R g8385 ( 
.A(n_7931),
.B(n_5298),
.Y(n_8385)
);

INVx1_ASAP7_75t_L g8386 ( 
.A(n_7719),
.Y(n_8386)
);

BUFx6f_ASAP7_75t_L g8387 ( 
.A(n_7552),
.Y(n_8387)
);

INVx1_ASAP7_75t_L g8388 ( 
.A(n_7724),
.Y(n_8388)
);

INVx2_ASAP7_75t_L g8389 ( 
.A(n_7725),
.Y(n_8389)
);

CKINVDCx5p33_ASAP7_75t_R g8390 ( 
.A(n_7955),
.Y(n_8390)
);

INVx2_ASAP7_75t_L g8391 ( 
.A(n_7744),
.Y(n_8391)
);

INVx1_ASAP7_75t_L g8392 ( 
.A(n_7746),
.Y(n_8392)
);

NOR2xp33_ASAP7_75t_L g8393 ( 
.A(n_7482),
.B(n_5300),
.Y(n_8393)
);

INVx1_ASAP7_75t_L g8394 ( 
.A(n_7758),
.Y(n_8394)
);

BUFx2_ASAP7_75t_L g8395 ( 
.A(n_7610),
.Y(n_8395)
);

INVx2_ASAP7_75t_L g8396 ( 
.A(n_8035),
.Y(n_8396)
);

CKINVDCx5p33_ASAP7_75t_R g8397 ( 
.A(n_7963),
.Y(n_8397)
);

CKINVDCx5p33_ASAP7_75t_R g8398 ( 
.A(n_7974),
.Y(n_8398)
);

CKINVDCx20_ASAP7_75t_R g8399 ( 
.A(n_7511),
.Y(n_8399)
);

INVx1_ASAP7_75t_L g8400 ( 
.A(n_7828),
.Y(n_8400)
);

CKINVDCx5p33_ASAP7_75t_R g8401 ( 
.A(n_7990),
.Y(n_8401)
);

CKINVDCx20_ASAP7_75t_R g8402 ( 
.A(n_7531),
.Y(n_8402)
);

INVx1_ASAP7_75t_L g8403 ( 
.A(n_7855),
.Y(n_8403)
);

NAND2xp33_ASAP7_75t_L g8404 ( 
.A(n_7626),
.B(n_5301),
.Y(n_8404)
);

NAND2xp5_ASAP7_75t_L g8405 ( 
.A(n_7770),
.B(n_5303),
.Y(n_8405)
);

OA21x2_ASAP7_75t_L g8406 ( 
.A1(n_7901),
.A2(n_7585),
.B(n_7572),
.Y(n_8406)
);

INVx1_ASAP7_75t_L g8407 ( 
.A(n_7863),
.Y(n_8407)
);

INVx1_ASAP7_75t_L g8408 ( 
.A(n_7862),
.Y(n_8408)
);

INVx2_ASAP7_75t_L g8409 ( 
.A(n_7864),
.Y(n_8409)
);

CKINVDCx5p33_ASAP7_75t_R g8410 ( 
.A(n_7946),
.Y(n_8410)
);

CKINVDCx20_ASAP7_75t_R g8411 ( 
.A(n_7997),
.Y(n_8411)
);

INVx1_ASAP7_75t_L g8412 ( 
.A(n_7876),
.Y(n_8412)
);

AOI22xp5_ASAP7_75t_L g8413 ( 
.A1(n_7496),
.A2(n_6035),
.B1(n_6074),
.B2(n_6045),
.Y(n_8413)
);

INVx2_ASAP7_75t_L g8414 ( 
.A(n_7475),
.Y(n_8414)
);

INVx1_ASAP7_75t_L g8415 ( 
.A(n_7559),
.Y(n_8415)
);

CKINVDCx5p33_ASAP7_75t_R g8416 ( 
.A(n_7951),
.Y(n_8416)
);

CKINVDCx5p33_ASAP7_75t_R g8417 ( 
.A(n_7952),
.Y(n_8417)
);

NAND2xp5_ASAP7_75t_L g8418 ( 
.A(n_7811),
.B(n_5304),
.Y(n_8418)
);

CKINVDCx5p33_ASAP7_75t_R g8419 ( 
.A(n_7958),
.Y(n_8419)
);

BUFx6f_ASAP7_75t_L g8420 ( 
.A(n_7557),
.Y(n_8420)
);

CKINVDCx5p33_ASAP7_75t_R g8421 ( 
.A(n_7980),
.Y(n_8421)
);

INVx2_ASAP7_75t_L g8422 ( 
.A(n_7480),
.Y(n_8422)
);

CKINVDCx5p33_ASAP7_75t_R g8423 ( 
.A(n_7988),
.Y(n_8423)
);

OA21x2_ASAP7_75t_L g8424 ( 
.A1(n_7773),
.A2(n_5414),
.B(n_5411),
.Y(n_8424)
);

CKINVDCx5p33_ASAP7_75t_R g8425 ( 
.A(n_7780),
.Y(n_8425)
);

CKINVDCx5p33_ASAP7_75t_R g8426 ( 
.A(n_7626),
.Y(n_8426)
);

INVx1_ASAP7_75t_L g8427 ( 
.A(n_7560),
.Y(n_8427)
);

CKINVDCx5p33_ASAP7_75t_R g8428 ( 
.A(n_7989),
.Y(n_8428)
);

INVx1_ASAP7_75t_L g8429 ( 
.A(n_7620),
.Y(n_8429)
);

CKINVDCx5p33_ASAP7_75t_R g8430 ( 
.A(n_7989),
.Y(n_8430)
);

CKINVDCx5p33_ASAP7_75t_R g8431 ( 
.A(n_7977),
.Y(n_8431)
);

INVx1_ASAP7_75t_L g8432 ( 
.A(n_7623),
.Y(n_8432)
);

NOR2xp33_ASAP7_75t_R g8433 ( 
.A(n_7604),
.B(n_6084),
.Y(n_8433)
);

INVx1_ASAP7_75t_L g8434 ( 
.A(n_7639),
.Y(n_8434)
);

NAND2xp5_ASAP7_75t_L g8435 ( 
.A(n_7543),
.B(n_5309),
.Y(n_8435)
);

INVx3_ASAP7_75t_L g8436 ( 
.A(n_7582),
.Y(n_8436)
);

INVx1_ASAP7_75t_L g8437 ( 
.A(n_7656),
.Y(n_8437)
);

INVx1_ASAP7_75t_L g8438 ( 
.A(n_7667),
.Y(n_8438)
);

INVx3_ASAP7_75t_L g8439 ( 
.A(n_7584),
.Y(n_8439)
);

CKINVDCx5p33_ASAP7_75t_R g8440 ( 
.A(n_7977),
.Y(n_8440)
);

INVx1_ASAP7_75t_L g8441 ( 
.A(n_7700),
.Y(n_8441)
);

CKINVDCx5p33_ASAP7_75t_R g8442 ( 
.A(n_7625),
.Y(n_8442)
);

NAND2xp5_ASAP7_75t_L g8443 ( 
.A(n_7692),
.B(n_5311),
.Y(n_8443)
);

CKINVDCx5p33_ASAP7_75t_R g8444 ( 
.A(n_7666),
.Y(n_8444)
);

OA21x2_ASAP7_75t_L g8445 ( 
.A1(n_7967),
.A2(n_5419),
.B(n_5418),
.Y(n_8445)
);

INVx1_ASAP7_75t_L g8446 ( 
.A(n_7738),
.Y(n_8446)
);

AND2x2_ASAP7_75t_L g8447 ( 
.A(n_7771),
.B(n_6104),
.Y(n_8447)
);

NOR2xp33_ASAP7_75t_L g8448 ( 
.A(n_7895),
.B(n_5316),
.Y(n_8448)
);

INVx2_ASAP7_75t_L g8449 ( 
.A(n_7481),
.Y(n_8449)
);

CKINVDCx5p33_ASAP7_75t_R g8450 ( 
.A(n_7683),
.Y(n_8450)
);

CKINVDCx5p33_ASAP7_75t_R g8451 ( 
.A(n_7712),
.Y(n_8451)
);

BUFx8_ASAP7_75t_L g8452 ( 
.A(n_7915),
.Y(n_8452)
);

CKINVDCx5p33_ASAP7_75t_R g8453 ( 
.A(n_7716),
.Y(n_8453)
);

INVx3_ASAP7_75t_L g8454 ( 
.A(n_7606),
.Y(n_8454)
);

NAND2xp5_ASAP7_75t_L g8455 ( 
.A(n_7634),
.B(n_5321),
.Y(n_8455)
);

AND2x2_ASAP7_75t_L g8456 ( 
.A(n_7927),
.B(n_6110),
.Y(n_8456)
);

BUFx3_ASAP7_75t_L g8457 ( 
.A(n_7910),
.Y(n_8457)
);

CKINVDCx5p33_ASAP7_75t_R g8458 ( 
.A(n_7748),
.Y(n_8458)
);

INVx1_ASAP7_75t_L g8459 ( 
.A(n_7777),
.Y(n_8459)
);

NAND2xp5_ASAP7_75t_L g8460 ( 
.A(n_7677),
.B(n_5322),
.Y(n_8460)
);

AND2x2_ASAP7_75t_L g8461 ( 
.A(n_7775),
.B(n_6119),
.Y(n_8461)
);

AND2x2_ASAP7_75t_L g8462 ( 
.A(n_7831),
.B(n_6133),
.Y(n_8462)
);

INVx1_ASAP7_75t_L g8463 ( 
.A(n_7792),
.Y(n_8463)
);

HB1xp67_ASAP7_75t_L g8464 ( 
.A(n_7568),
.Y(n_8464)
);

OR2x2_ASAP7_75t_L g8465 ( 
.A(n_7995),
.B(n_5395),
.Y(n_8465)
);

INVx3_ASAP7_75t_L g8466 ( 
.A(n_7613),
.Y(n_8466)
);

CKINVDCx5p33_ASAP7_75t_R g8467 ( 
.A(n_7806),
.Y(n_8467)
);

INVx1_ASAP7_75t_L g8468 ( 
.A(n_7793),
.Y(n_8468)
);

CKINVDCx20_ASAP7_75t_R g8469 ( 
.A(n_7497),
.Y(n_8469)
);

CKINVDCx5p33_ASAP7_75t_R g8470 ( 
.A(n_7915),
.Y(n_8470)
);

CKINVDCx5p33_ASAP7_75t_R g8471 ( 
.A(n_7487),
.Y(n_8471)
);

NAND2xp5_ASAP7_75t_SL g8472 ( 
.A(n_7723),
.B(n_5324),
.Y(n_8472)
);

NOR2xp67_ASAP7_75t_L g8473 ( 
.A(n_7542),
.B(n_4330),
.Y(n_8473)
);

INVx1_ASAP7_75t_L g8474 ( 
.A(n_7797),
.Y(n_8474)
);

CKINVDCx20_ASAP7_75t_R g8475 ( 
.A(n_8045),
.Y(n_8475)
);

AND2x2_ASAP7_75t_L g8476 ( 
.A(n_8010),
.B(n_6160),
.Y(n_8476)
);

INVx1_ASAP7_75t_L g8477 ( 
.A(n_7802),
.Y(n_8477)
);

BUFx10_ASAP7_75t_L g8478 ( 
.A(n_7954),
.Y(n_8478)
);

INVx1_ASAP7_75t_L g8479 ( 
.A(n_7803),
.Y(n_8479)
);

AND2x4_ASAP7_75t_L g8480 ( 
.A(n_8049),
.B(n_5421),
.Y(n_8480)
);

INVx3_ASAP7_75t_L g8481 ( 
.A(n_7621),
.Y(n_8481)
);

HB1xp67_ASAP7_75t_L g8482 ( 
.A(n_7570),
.Y(n_8482)
);

CKINVDCx5p33_ASAP7_75t_R g8483 ( 
.A(n_7587),
.Y(n_8483)
);

INVx2_ASAP7_75t_L g8484 ( 
.A(n_7498),
.Y(n_8484)
);

INVx1_ASAP7_75t_L g8485 ( 
.A(n_7809),
.Y(n_8485)
);

INVx2_ASAP7_75t_L g8486 ( 
.A(n_7512),
.Y(n_8486)
);

CKINVDCx20_ASAP7_75t_R g8487 ( 
.A(n_7599),
.Y(n_8487)
);

INVx1_ASAP7_75t_L g8488 ( 
.A(n_7887),
.Y(n_8488)
);

INVxp67_ASAP7_75t_L g8489 ( 
.A(n_7615),
.Y(n_8489)
);

INVx1_ASAP7_75t_L g8490 ( 
.A(n_7898),
.Y(n_8490)
);

CKINVDCx5p33_ASAP7_75t_R g8491 ( 
.A(n_7969),
.Y(n_8491)
);

INVx1_ASAP7_75t_L g8492 ( 
.A(n_7813),
.Y(n_8492)
);

BUFx6f_ASAP7_75t_L g8493 ( 
.A(n_7630),
.Y(n_8493)
);

CKINVDCx8_ASAP7_75t_R g8494 ( 
.A(n_7675),
.Y(n_8494)
);

NAND2xp5_ASAP7_75t_L g8495 ( 
.A(n_7735),
.B(n_5326),
.Y(n_8495)
);

HB1xp67_ASAP7_75t_L g8496 ( 
.A(n_7975),
.Y(n_8496)
);

AND2x2_ASAP7_75t_L g8497 ( 
.A(n_7603),
.B(n_6181),
.Y(n_8497)
);

INVx2_ASAP7_75t_L g8498 ( 
.A(n_7515),
.Y(n_8498)
);

HB1xp67_ASAP7_75t_L g8499 ( 
.A(n_7981),
.Y(n_8499)
);

INVx1_ASAP7_75t_L g8500 ( 
.A(n_7838),
.Y(n_8500)
);

CKINVDCx5p33_ASAP7_75t_R g8501 ( 
.A(n_7933),
.Y(n_8501)
);

CKINVDCx16_ASAP7_75t_R g8502 ( 
.A(n_7833),
.Y(n_8502)
);

INVx1_ASAP7_75t_L g8503 ( 
.A(n_7851),
.Y(n_8503)
);

CKINVDCx5p33_ASAP7_75t_R g8504 ( 
.A(n_7929),
.Y(n_8504)
);

INVx1_ASAP7_75t_L g8505 ( 
.A(n_7847),
.Y(n_8505)
);

INVx2_ASAP7_75t_L g8506 ( 
.A(n_8000),
.Y(n_8506)
);

INVx2_ASAP7_75t_L g8507 ( 
.A(n_8009),
.Y(n_8507)
);

INVx2_ASAP7_75t_L g8508 ( 
.A(n_8019),
.Y(n_8508)
);

NAND2xp5_ASAP7_75t_SL g8509 ( 
.A(n_7753),
.B(n_5331),
.Y(n_8509)
);

NOR2xp33_ASAP7_75t_L g8510 ( 
.A(n_7908),
.B(n_5335),
.Y(n_8510)
);

CKINVDCx20_ASAP7_75t_R g8511 ( 
.A(n_7751),
.Y(n_8511)
);

BUFx6f_ASAP7_75t_L g8512 ( 
.A(n_7637),
.Y(n_8512)
);

INVx2_ASAP7_75t_L g8513 ( 
.A(n_8026),
.Y(n_8513)
);

INVx1_ASAP7_75t_L g8514 ( 
.A(n_7909),
.Y(n_8514)
);

CKINVDCx5p33_ASAP7_75t_R g8515 ( 
.A(n_7675),
.Y(n_8515)
);

NOR2xp67_ASAP7_75t_L g8516 ( 
.A(n_7747),
.B(n_4331),
.Y(n_8516)
);

NAND2xp5_ASAP7_75t_L g8517 ( 
.A(n_7711),
.B(n_5336),
.Y(n_8517)
);

INVx1_ASAP7_75t_L g8518 ( 
.A(n_7893),
.Y(n_8518)
);

INVx2_ASAP7_75t_L g8519 ( 
.A(n_8036),
.Y(n_8519)
);

INVx2_ASAP7_75t_L g8520 ( 
.A(n_8042),
.Y(n_8520)
);

INVx1_ASAP7_75t_L g8521 ( 
.A(n_8043),
.Y(n_8521)
);

NAND2xp5_ASAP7_75t_SL g8522 ( 
.A(n_7826),
.B(n_5344),
.Y(n_8522)
);

INVx1_ASAP7_75t_L g8523 ( 
.A(n_8046),
.Y(n_8523)
);

AND2x4_ASAP7_75t_L g8524 ( 
.A(n_7640),
.B(n_5425),
.Y(n_8524)
);

CKINVDCx5p33_ASAP7_75t_R g8525 ( 
.A(n_7709),
.Y(n_8525)
);

INVx1_ASAP7_75t_L g8526 ( 
.A(n_7849),
.Y(n_8526)
);

HB1xp67_ASAP7_75t_L g8527 ( 
.A(n_7936),
.Y(n_8527)
);

CKINVDCx5p33_ASAP7_75t_R g8528 ( 
.A(n_7709),
.Y(n_8528)
);

INVx2_ASAP7_75t_L g8529 ( 
.A(n_7669),
.Y(n_8529)
);

NOR2xp33_ASAP7_75t_R g8530 ( 
.A(n_7938),
.B(n_6205),
.Y(n_8530)
);

CKINVDCx5p33_ASAP7_75t_R g8531 ( 
.A(n_7631),
.Y(n_8531)
);

NOR2xp33_ASAP7_75t_L g8532 ( 
.A(n_8029),
.B(n_5345),
.Y(n_8532)
);

CKINVDCx5p33_ASAP7_75t_R g8533 ( 
.A(n_7608),
.Y(n_8533)
);

CKINVDCx5p33_ASAP7_75t_R g8534 ( 
.A(n_7935),
.Y(n_8534)
);

INVx2_ASAP7_75t_L g8535 ( 
.A(n_7836),
.Y(n_8535)
);

BUFx6f_ASAP7_75t_L g8536 ( 
.A(n_7649),
.Y(n_8536)
);

INVx1_ASAP7_75t_L g8537 ( 
.A(n_7493),
.Y(n_8537)
);

BUFx2_ASAP7_75t_L g8538 ( 
.A(n_7905),
.Y(n_8538)
);

CKINVDCx5p33_ASAP7_75t_R g8539 ( 
.A(n_7934),
.Y(n_8539)
);

HB1xp67_ASAP7_75t_L g8540 ( 
.A(n_7940),
.Y(n_8540)
);

INVxp67_ASAP7_75t_L g8541 ( 
.A(n_7529),
.Y(n_8541)
);

CKINVDCx20_ASAP7_75t_R g8542 ( 
.A(n_7745),
.Y(n_8542)
);

CKINVDCx5p33_ASAP7_75t_R g8543 ( 
.A(n_7961),
.Y(n_8543)
);

INVx2_ASAP7_75t_L g8544 ( 
.A(n_7842),
.Y(n_8544)
);

INVx1_ASAP7_75t_L g8545 ( 
.A(n_7505),
.Y(n_8545)
);

OR2x6_ASAP7_75t_L g8546 ( 
.A(n_7762),
.B(n_5427),
.Y(n_8546)
);

AND2x2_ASAP7_75t_L g8547 ( 
.A(n_8040),
.B(n_6239),
.Y(n_8547)
);

INVxp67_ASAP7_75t_L g8548 ( 
.A(n_7533),
.Y(n_8548)
);

NOR2xp33_ASAP7_75t_L g8549 ( 
.A(n_7903),
.B(n_5346),
.Y(n_8549)
);

NOR2xp33_ASAP7_75t_R g8550 ( 
.A(n_7721),
.B(n_6275),
.Y(n_8550)
);

INVx1_ASAP7_75t_L g8551 ( 
.A(n_7896),
.Y(n_8551)
);

CKINVDCx20_ASAP7_75t_R g8552 ( 
.A(n_7706),
.Y(n_8552)
);

INVx1_ASAP7_75t_L g8553 ( 
.A(n_7919),
.Y(n_8553)
);

INVx1_ASAP7_75t_L g8554 ( 
.A(n_7921),
.Y(n_8554)
);

AND2x2_ASAP7_75t_L g8555 ( 
.A(n_7494),
.B(n_6298),
.Y(n_8555)
);

CKINVDCx20_ASAP7_75t_R g8556 ( 
.A(n_7489),
.Y(n_8556)
);

CKINVDCx5p33_ASAP7_75t_R g8557 ( 
.A(n_7591),
.Y(n_8557)
);

INVx1_ASAP7_75t_L g8558 ( 
.A(n_7844),
.Y(n_8558)
);

AND2x2_ASAP7_75t_SL g8559 ( 
.A(n_8014),
.B(n_5728),
.Y(n_8559)
);

HB1xp67_ASAP7_75t_L g8560 ( 
.A(n_7924),
.Y(n_8560)
);

INVx1_ASAP7_75t_L g8561 ( 
.A(n_7845),
.Y(n_8561)
);

INVx1_ASAP7_75t_L g8562 ( 
.A(n_7867),
.Y(n_8562)
);

BUFx6f_ASAP7_75t_L g8563 ( 
.A(n_7659),
.Y(n_8563)
);

HB1xp67_ASAP7_75t_L g8564 ( 
.A(n_7932),
.Y(n_8564)
);

INVx2_ASAP7_75t_L g8565 ( 
.A(n_7544),
.Y(n_8565)
);

BUFx2_ASAP7_75t_L g8566 ( 
.A(n_7474),
.Y(n_8566)
);

INVx2_ASAP7_75t_L g8567 ( 
.A(n_7662),
.Y(n_8567)
);

NAND2xp5_ASAP7_75t_L g8568 ( 
.A(n_7521),
.B(n_5347),
.Y(n_8568)
);

CKINVDCx5p33_ASAP7_75t_R g8569 ( 
.A(n_7633),
.Y(n_8569)
);

CKINVDCx20_ASAP7_75t_R g8570 ( 
.A(n_7573),
.Y(n_8570)
);

AND2x6_ASAP7_75t_L g8571 ( 
.A(n_7868),
.B(n_5428),
.Y(n_8571)
);

NOR2xp67_ASAP7_75t_L g8572 ( 
.A(n_7791),
.B(n_4332),
.Y(n_8572)
);

INVx1_ASAP7_75t_L g8573 ( 
.A(n_7890),
.Y(n_8573)
);

AND2x4_ASAP7_75t_L g8574 ( 
.A(n_7663),
.B(n_5429),
.Y(n_8574)
);

INVx3_ASAP7_75t_L g8575 ( 
.A(n_7668),
.Y(n_8575)
);

HB1xp67_ASAP7_75t_L g8576 ( 
.A(n_7779),
.Y(n_8576)
);

INVx1_ASAP7_75t_L g8577 ( 
.A(n_7678),
.Y(n_8577)
);

CKINVDCx5p33_ASAP7_75t_R g8578 ( 
.A(n_7822),
.Y(n_8578)
);

AND2x4_ASAP7_75t_L g8579 ( 
.A(n_7682),
.B(n_5431),
.Y(n_8579)
);

CKINVDCx20_ASAP7_75t_R g8580 ( 
.A(n_7734),
.Y(n_8580)
);

AND2x2_ASAP7_75t_L g8581 ( 
.A(n_7491),
.B(n_6301),
.Y(n_8581)
);

INVx1_ASAP7_75t_L g8582 ( 
.A(n_7686),
.Y(n_8582)
);

CKINVDCx5p33_ASAP7_75t_R g8583 ( 
.A(n_7886),
.Y(n_8583)
);

BUFx6f_ASAP7_75t_L g8584 ( 
.A(n_7688),
.Y(n_8584)
);

INVx3_ASAP7_75t_L g8585 ( 
.A(n_7690),
.Y(n_8585)
);

INVx1_ASAP7_75t_L g8586 ( 
.A(n_7694),
.Y(n_8586)
);

NAND2xp33_ASAP7_75t_R g8587 ( 
.A(n_7800),
.B(n_5349),
.Y(n_8587)
);

NAND2xp5_ASAP7_75t_L g8588 ( 
.A(n_7510),
.B(n_5351),
.Y(n_8588)
);

INVx1_ASAP7_75t_L g8589 ( 
.A(n_7707),
.Y(n_8589)
);

INVx1_ASAP7_75t_L g8590 ( 
.A(n_7720),
.Y(n_8590)
);

INVx1_ASAP7_75t_L g8591 ( 
.A(n_7729),
.Y(n_8591)
);

BUFx6f_ASAP7_75t_L g8592 ( 
.A(n_7733),
.Y(n_8592)
);

CKINVDCx8_ASAP7_75t_R g8593 ( 
.A(n_7812),
.Y(n_8593)
);

BUFx2_ASAP7_75t_L g8594 ( 
.A(n_7642),
.Y(n_8594)
);

INVx2_ASAP7_75t_L g8595 ( 
.A(n_7741),
.Y(n_8595)
);

CKINVDCx20_ASAP7_75t_R g8596 ( 
.A(n_7757),
.Y(n_8596)
);

INVx1_ASAP7_75t_L g8597 ( 
.A(n_7743),
.Y(n_8597)
);

INVx1_ASAP7_75t_L g8598 ( 
.A(n_7769),
.Y(n_8598)
);

BUFx6f_ASAP7_75t_L g8599 ( 
.A(n_7781),
.Y(n_8599)
);

HB1xp67_ASAP7_75t_L g8600 ( 
.A(n_7814),
.Y(n_8600)
);

AND2x4_ASAP7_75t_L g8601 ( 
.A(n_7782),
.B(n_5435),
.Y(n_8601)
);

CKINVDCx20_ASAP7_75t_R g8602 ( 
.A(n_7767),
.Y(n_8602)
);

CKINVDCx5p33_ASAP7_75t_R g8603 ( 
.A(n_7897),
.Y(n_8603)
);

BUFx6f_ASAP7_75t_SL g8604 ( 
.A(n_7843),
.Y(n_8604)
);

NOR2xp33_ASAP7_75t_R g8605 ( 
.A(n_7530),
.B(n_6307),
.Y(n_8605)
);

CKINVDCx20_ASAP7_75t_R g8606 ( 
.A(n_7801),
.Y(n_8606)
);

NOR2xp33_ASAP7_75t_R g8607 ( 
.A(n_7635),
.B(n_6341),
.Y(n_8607)
);

CKINVDCx5p33_ASAP7_75t_R g8608 ( 
.A(n_7514),
.Y(n_8608)
);

CKINVDCx20_ASAP7_75t_R g8609 ( 
.A(n_7805),
.Y(n_8609)
);

INVx2_ASAP7_75t_L g8610 ( 
.A(n_7551),
.Y(n_8610)
);

INVx1_ASAP7_75t_L g8611 ( 
.A(n_7664),
.Y(n_8611)
);

INVx3_ASAP7_75t_L g8612 ( 
.A(n_7702),
.Y(n_8612)
);

CKINVDCx5p33_ASAP7_75t_R g8613 ( 
.A(n_7597),
.Y(n_8613)
);

INVx1_ASAP7_75t_L g8614 ( 
.A(n_7710),
.Y(n_8614)
);

INVx1_ASAP7_75t_L g8615 ( 
.A(n_7881),
.Y(n_8615)
);

INVx1_ASAP7_75t_L g8616 ( 
.A(n_7646),
.Y(n_8616)
);

INVx1_ASAP7_75t_L g8617 ( 
.A(n_7660),
.Y(n_8617)
);

CKINVDCx5p33_ASAP7_75t_R g8618 ( 
.A(n_7697),
.Y(n_8618)
);

BUFx6f_ASAP7_75t_L g8619 ( 
.A(n_7516),
.Y(n_8619)
);

INVx2_ASAP7_75t_L g8620 ( 
.A(n_7602),
.Y(n_8620)
);

INVx1_ASAP7_75t_L g8621 ( 
.A(n_8061),
.Y(n_8621)
);

AND2x2_ASAP7_75t_L g8622 ( 
.A(n_8140),
.B(n_7671),
.Y(n_8622)
);

INVx2_ASAP7_75t_L g8623 ( 
.A(n_8059),
.Y(n_8623)
);

INVx2_ASAP7_75t_L g8624 ( 
.A(n_8068),
.Y(n_8624)
);

INVx1_ASAP7_75t_L g8625 ( 
.A(n_8064),
.Y(n_8625)
);

INVx2_ASAP7_75t_L g8626 ( 
.A(n_8072),
.Y(n_8626)
);

NAND2xp5_ASAP7_75t_L g8627 ( 
.A(n_8070),
.B(n_7674),
.Y(n_8627)
);

INVx1_ASAP7_75t_L g8628 ( 
.A(n_8065),
.Y(n_8628)
);

BUFx6f_ASAP7_75t_L g8629 ( 
.A(n_8063),
.Y(n_8629)
);

INVx1_ASAP7_75t_L g8630 ( 
.A(n_8069),
.Y(n_8630)
);

INVx2_ASAP7_75t_L g8631 ( 
.A(n_8093),
.Y(n_8631)
);

NAND2x1_ASAP7_75t_L g8632 ( 
.A(n_8396),
.B(n_7652),
.Y(n_8632)
);

AOI22xp5_ASAP7_75t_L g8633 ( 
.A1(n_8241),
.A2(n_7722),
.B1(n_7794),
.B2(n_7699),
.Y(n_8633)
);

NAND2xp5_ASAP7_75t_SL g8634 ( 
.A(n_8277),
.B(n_7835),
.Y(n_8634)
);

HB1xp67_ASAP7_75t_L g8635 ( 
.A(n_8058),
.Y(n_8635)
);

OAI22xp5_ASAP7_75t_SL g8636 ( 
.A1(n_8469),
.A2(n_6384),
.B1(n_6400),
.B2(n_6365),
.Y(n_8636)
);

INVx3_ASAP7_75t_L g8637 ( 
.A(n_8387),
.Y(n_8637)
);

INVx3_ASAP7_75t_SL g8638 ( 
.A(n_8328),
.Y(n_8638)
);

INVxp67_ASAP7_75t_L g8639 ( 
.A(n_8060),
.Y(n_8639)
);

CKINVDCx8_ASAP7_75t_R g8640 ( 
.A(n_8186),
.Y(n_8640)
);

NAND2xp5_ASAP7_75t_L g8641 ( 
.A(n_8306),
.B(n_7566),
.Y(n_8641)
);

INVx1_ASAP7_75t_L g8642 ( 
.A(n_8071),
.Y(n_8642)
);

OR2x2_ASAP7_75t_L g8643 ( 
.A(n_8229),
.B(n_5353),
.Y(n_8643)
);

AND2x4_ASAP7_75t_L g8644 ( 
.A(n_8347),
.B(n_8351),
.Y(n_8644)
);

BUFx2_ASAP7_75t_L g8645 ( 
.A(n_8487),
.Y(n_8645)
);

INVx1_ASAP7_75t_L g8646 ( 
.A(n_8076),
.Y(n_8646)
);

OAI22xp5_ASAP7_75t_SL g8647 ( 
.A1(n_8475),
.A2(n_6408),
.B1(n_6417),
.B2(n_6403),
.Y(n_8647)
);

INVx1_ASAP7_75t_L g8648 ( 
.A(n_8077),
.Y(n_8648)
);

INVx1_ASAP7_75t_L g8649 ( 
.A(n_8079),
.Y(n_8649)
);

NOR2xp33_ASAP7_75t_SL g8650 ( 
.A(n_8089),
.B(n_6421),
.Y(n_8650)
);

BUFx6f_ASAP7_75t_L g8651 ( 
.A(n_8063),
.Y(n_8651)
);

AOI22xp5_ASAP7_75t_L g8652 ( 
.A1(n_8448),
.A2(n_7605),
.B1(n_7622),
.B2(n_7580),
.Y(n_8652)
);

AOI22xp5_ASAP7_75t_L g8653 ( 
.A1(n_8510),
.A2(n_7761),
.B1(n_7778),
.B2(n_7756),
.Y(n_8653)
);

INVx1_ASAP7_75t_L g8654 ( 
.A(n_8080),
.Y(n_8654)
);

NAND2xp5_ASAP7_75t_L g8655 ( 
.A(n_8514),
.B(n_5354),
.Y(n_8655)
);

INVx2_ASAP7_75t_L g8656 ( 
.A(n_8109),
.Y(n_8656)
);

INVx1_ASAP7_75t_L g8657 ( 
.A(n_8081),
.Y(n_8657)
);

INVx1_ASAP7_75t_L g8658 ( 
.A(n_8084),
.Y(n_8658)
);

NOR2xp33_ASAP7_75t_L g8659 ( 
.A(n_8088),
.B(n_6434),
.Y(n_8659)
);

BUFx8_ASAP7_75t_L g8660 ( 
.A(n_8604),
.Y(n_8660)
);

INVx1_ASAP7_75t_L g8661 ( 
.A(n_8087),
.Y(n_8661)
);

INVx2_ASAP7_75t_L g8662 ( 
.A(n_8111),
.Y(n_8662)
);

INVx1_ASAP7_75t_L g8663 ( 
.A(n_8090),
.Y(n_8663)
);

BUFx6f_ASAP7_75t_L g8664 ( 
.A(n_8115),
.Y(n_8664)
);

INVx1_ASAP7_75t_L g8665 ( 
.A(n_8095),
.Y(n_8665)
);

INVx1_ASAP7_75t_L g8666 ( 
.A(n_8100),
.Y(n_8666)
);

INVx1_ASAP7_75t_L g8667 ( 
.A(n_8101),
.Y(n_8667)
);

INVx2_ASAP7_75t_L g8668 ( 
.A(n_8248),
.Y(n_8668)
);

NAND2xp5_ASAP7_75t_L g8669 ( 
.A(n_8537),
.B(n_8545),
.Y(n_8669)
);

BUFx6f_ASAP7_75t_L g8670 ( 
.A(n_8115),
.Y(n_8670)
);

BUFx6f_ASAP7_75t_L g8671 ( 
.A(n_8183),
.Y(n_8671)
);

OAI22xp5_ASAP7_75t_SL g8672 ( 
.A1(n_8372),
.A2(n_6470),
.B1(n_6459),
.B2(n_5359),
.Y(n_8672)
);

INVx1_ASAP7_75t_L g8673 ( 
.A(n_8103),
.Y(n_8673)
);

AND2x6_ASAP7_75t_L g8674 ( 
.A(n_8562),
.B(n_5437),
.Y(n_8674)
);

AND2x2_ASAP7_75t_L g8675 ( 
.A(n_8235),
.B(n_5355),
.Y(n_8675)
);

INVx2_ASAP7_75t_L g8676 ( 
.A(n_8259),
.Y(n_8676)
);

INVx1_ASAP7_75t_L g8677 ( 
.A(n_8112),
.Y(n_8677)
);

NAND2xp5_ASAP7_75t_L g8678 ( 
.A(n_8616),
.B(n_5360),
.Y(n_8678)
);

NAND2xp5_ASAP7_75t_L g8679 ( 
.A(n_8617),
.B(n_5365),
.Y(n_8679)
);

AND2x2_ASAP7_75t_L g8680 ( 
.A(n_8280),
.B(n_5366),
.Y(n_8680)
);

HB1xp67_ASAP7_75t_L g8681 ( 
.A(n_8167),
.Y(n_8681)
);

INVx1_ASAP7_75t_L g8682 ( 
.A(n_8113),
.Y(n_8682)
);

INVx1_ASAP7_75t_L g8683 ( 
.A(n_8117),
.Y(n_8683)
);

INVx2_ASAP7_75t_L g8684 ( 
.A(n_8266),
.Y(n_8684)
);

NAND2xp5_ASAP7_75t_L g8685 ( 
.A(n_8573),
.B(n_5371),
.Y(n_8685)
);

NAND2xp33_ASAP7_75t_SL g8686 ( 
.A(n_8534),
.B(n_5372),
.Y(n_8686)
);

BUFx6f_ASAP7_75t_L g8687 ( 
.A(n_8183),
.Y(n_8687)
);

INVxp67_ASAP7_75t_L g8688 ( 
.A(n_8124),
.Y(n_8688)
);

BUFx2_ASAP7_75t_L g8689 ( 
.A(n_8169),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_8120),
.Y(n_8690)
);

INVx1_ASAP7_75t_SL g8691 ( 
.A(n_8232),
.Y(n_8691)
);

OAI22xp5_ASAP7_75t_SL g8692 ( 
.A1(n_8335),
.A2(n_5377),
.B1(n_5378),
.B2(n_5375),
.Y(n_8692)
);

INVx1_ASAP7_75t_L g8693 ( 
.A(n_8122),
.Y(n_8693)
);

NAND2xp5_ASAP7_75t_SL g8694 ( 
.A(n_8365),
.B(n_5380),
.Y(n_8694)
);

INVx1_ASAP7_75t_L g8695 ( 
.A(n_8123),
.Y(n_8695)
);

INVx1_ASAP7_75t_SL g8696 ( 
.A(n_8425),
.Y(n_8696)
);

BUFx6f_ASAP7_75t_L g8697 ( 
.A(n_8225),
.Y(n_8697)
);

INVx1_ASAP7_75t_L g8698 ( 
.A(n_8131),
.Y(n_8698)
);

NAND2xp5_ASAP7_75t_SL g8699 ( 
.A(n_8368),
.B(n_8390),
.Y(n_8699)
);

INVx1_ASAP7_75t_L g8700 ( 
.A(n_8138),
.Y(n_8700)
);

XNOR2xp5_ASAP7_75t_L g8701 ( 
.A(n_8083),
.B(n_4333),
.Y(n_8701)
);

HB1xp67_ASAP7_75t_L g8702 ( 
.A(n_8205),
.Y(n_8702)
);

INVx1_ASAP7_75t_L g8703 ( 
.A(n_8142),
.Y(n_8703)
);

NAND2xp5_ASAP7_75t_L g8704 ( 
.A(n_8283),
.B(n_5381),
.Y(n_8704)
);

INVx2_ASAP7_75t_L g8705 ( 
.A(n_8271),
.Y(n_8705)
);

HB1xp67_ASAP7_75t_L g8706 ( 
.A(n_8482),
.Y(n_8706)
);

NAND2xp5_ASAP7_75t_SL g8707 ( 
.A(n_8397),
.B(n_5383),
.Y(n_8707)
);

INVx2_ASAP7_75t_L g8708 ( 
.A(n_8326),
.Y(n_8708)
);

BUFx6f_ASAP7_75t_L g8709 ( 
.A(n_8225),
.Y(n_8709)
);

INVx1_ASAP7_75t_L g8710 ( 
.A(n_8143),
.Y(n_8710)
);

OAI22xp5_ASAP7_75t_L g8711 ( 
.A1(n_8548),
.A2(n_5389),
.B1(n_5390),
.B2(n_5385),
.Y(n_8711)
);

NOR2xp33_ASAP7_75t_L g8712 ( 
.A(n_8147),
.B(n_5391),
.Y(n_8712)
);

INVx2_ASAP7_75t_L g8713 ( 
.A(n_8333),
.Y(n_8713)
);

INVx1_ASAP7_75t_L g8714 ( 
.A(n_8144),
.Y(n_8714)
);

INVxp67_ASAP7_75t_L g8715 ( 
.A(n_8497),
.Y(n_8715)
);

AOI22xp5_ASAP7_75t_L g8716 ( 
.A1(n_8174),
.A2(n_5393),
.B1(n_5394),
.B2(n_5392),
.Y(n_8716)
);

AND2x2_ASAP7_75t_L g8717 ( 
.A(n_8151),
.B(n_5399),
.Y(n_8717)
);

NOR2xp33_ASAP7_75t_L g8718 ( 
.A(n_8091),
.B(n_5401),
.Y(n_8718)
);

AOI22xp5_ASAP7_75t_L g8719 ( 
.A1(n_8211),
.A2(n_5404),
.B1(n_5406),
.B2(n_5403),
.Y(n_8719)
);

INVx2_ASAP7_75t_L g8720 ( 
.A(n_8308),
.Y(n_8720)
);

BUFx6f_ASAP7_75t_SL g8721 ( 
.A(n_8319),
.Y(n_8721)
);

HB1xp67_ASAP7_75t_L g8722 ( 
.A(n_8464),
.Y(n_8722)
);

INVx1_ASAP7_75t_L g8723 ( 
.A(n_8149),
.Y(n_8723)
);

INVx1_ASAP7_75t_L g8724 ( 
.A(n_8150),
.Y(n_8724)
);

INVx1_ASAP7_75t_L g8725 ( 
.A(n_8153),
.Y(n_8725)
);

HB1xp67_ASAP7_75t_L g8726 ( 
.A(n_8265),
.Y(n_8726)
);

CKINVDCx20_ASAP7_75t_R g8727 ( 
.A(n_8086),
.Y(n_8727)
);

INVx3_ASAP7_75t_L g8728 ( 
.A(n_8387),
.Y(n_8728)
);

INVx1_ASAP7_75t_L g8729 ( 
.A(n_8156),
.Y(n_8729)
);

INVx1_ASAP7_75t_L g8730 ( 
.A(n_8166),
.Y(n_8730)
);

BUFx6f_ASAP7_75t_L g8731 ( 
.A(n_8236),
.Y(n_8731)
);

INVx2_ASAP7_75t_L g8732 ( 
.A(n_8309),
.Y(n_8732)
);

BUFx6f_ASAP7_75t_L g8733 ( 
.A(n_8236),
.Y(n_8733)
);

INVx1_ASAP7_75t_L g8734 ( 
.A(n_8171),
.Y(n_8734)
);

INVx1_ASAP7_75t_L g8735 ( 
.A(n_8180),
.Y(n_8735)
);

INVx1_ASAP7_75t_L g8736 ( 
.A(n_8181),
.Y(n_8736)
);

INVx1_ASAP7_75t_L g8737 ( 
.A(n_8182),
.Y(n_8737)
);

NAND2xp5_ASAP7_75t_L g8738 ( 
.A(n_8246),
.B(n_8383),
.Y(n_8738)
);

NAND2xp5_ASAP7_75t_SL g8739 ( 
.A(n_8398),
.B(n_5407),
.Y(n_8739)
);

OR2x2_ASAP7_75t_L g8740 ( 
.A(n_8253),
.B(n_5408),
.Y(n_8740)
);

INVx1_ASAP7_75t_L g8741 ( 
.A(n_8187),
.Y(n_8741)
);

INVx2_ASAP7_75t_L g8742 ( 
.A(n_8195),
.Y(n_8742)
);

INVx1_ASAP7_75t_L g8743 ( 
.A(n_8196),
.Y(n_8743)
);

INVx1_ASAP7_75t_L g8744 ( 
.A(n_8199),
.Y(n_8744)
);

NAND2xp5_ASAP7_75t_SL g8745 ( 
.A(n_8401),
.B(n_5410),
.Y(n_8745)
);

INVx1_ASAP7_75t_L g8746 ( 
.A(n_8201),
.Y(n_8746)
);

HB1xp67_ASAP7_75t_L g8747 ( 
.A(n_8242),
.Y(n_8747)
);

OAI22xp5_ASAP7_75t_SL g8748 ( 
.A1(n_8511),
.A2(n_8556),
.B1(n_8596),
.B2(n_8580),
.Y(n_8748)
);

HB1xp67_ASAP7_75t_L g8749 ( 
.A(n_8501),
.Y(n_8749)
);

NAND2xp5_ASAP7_75t_L g8750 ( 
.A(n_8393),
.B(n_5412),
.Y(n_8750)
);

NAND2xp5_ASAP7_75t_SL g8751 ( 
.A(n_8502),
.B(n_5415),
.Y(n_8751)
);

INVx1_ASAP7_75t_L g8752 ( 
.A(n_8204),
.Y(n_8752)
);

INVx1_ASAP7_75t_L g8753 ( 
.A(n_8206),
.Y(n_8753)
);

HB1xp67_ASAP7_75t_L g8754 ( 
.A(n_8483),
.Y(n_8754)
);

INVx1_ASAP7_75t_L g8755 ( 
.A(n_8212),
.Y(n_8755)
);

INVx2_ASAP7_75t_L g8756 ( 
.A(n_8215),
.Y(n_8756)
);

BUFx6f_ASAP7_75t_L g8757 ( 
.A(n_8240),
.Y(n_8757)
);

BUFx6f_ASAP7_75t_SL g8758 ( 
.A(n_8296),
.Y(n_8758)
);

INVx1_ASAP7_75t_L g8759 ( 
.A(n_8219),
.Y(n_8759)
);

INVx1_ASAP7_75t_L g8760 ( 
.A(n_8220),
.Y(n_8760)
);

NAND2xp5_ASAP7_75t_SL g8761 ( 
.A(n_8410),
.B(n_5417),
.Y(n_8761)
);

BUFx6f_ASAP7_75t_L g8762 ( 
.A(n_8240),
.Y(n_8762)
);

NAND2x1_ASAP7_75t_L g8763 ( 
.A(n_8565),
.B(n_6334),
.Y(n_8763)
);

INVx1_ASAP7_75t_L g8764 ( 
.A(n_8224),
.Y(n_8764)
);

INVx2_ASAP7_75t_L g8765 ( 
.A(n_8226),
.Y(n_8765)
);

NAND2xp33_ASAP7_75t_SL g8766 ( 
.A(n_8261),
.B(n_8267),
.Y(n_8766)
);

OAI22xp5_ASAP7_75t_SL g8767 ( 
.A1(n_8602),
.A2(n_5423),
.B1(n_5424),
.B2(n_5422),
.Y(n_8767)
);

BUFx2_ASAP7_75t_L g8768 ( 
.A(n_8190),
.Y(n_8768)
);

INVx2_ASAP7_75t_L g8769 ( 
.A(n_8245),
.Y(n_8769)
);

INVx1_ASAP7_75t_L g8770 ( 
.A(n_8256),
.Y(n_8770)
);

INVx1_ASAP7_75t_L g8771 ( 
.A(n_8262),
.Y(n_8771)
);

INVx1_ASAP7_75t_L g8772 ( 
.A(n_8264),
.Y(n_8772)
);

INVx1_ASAP7_75t_L g8773 ( 
.A(n_8273),
.Y(n_8773)
);

INVx2_ASAP7_75t_L g8774 ( 
.A(n_8278),
.Y(n_8774)
);

INVx1_ASAP7_75t_L g8775 ( 
.A(n_8285),
.Y(n_8775)
);

INVx2_ASAP7_75t_L g8776 ( 
.A(n_8294),
.Y(n_8776)
);

INVx1_ASAP7_75t_L g8777 ( 
.A(n_8299),
.Y(n_8777)
);

NAND2xp5_ASAP7_75t_SL g8778 ( 
.A(n_8416),
.B(n_5432),
.Y(n_8778)
);

INVx3_ASAP7_75t_L g8779 ( 
.A(n_8420),
.Y(n_8779)
);

INVx2_ASAP7_75t_L g8780 ( 
.A(n_8301),
.Y(n_8780)
);

HB1xp67_ASAP7_75t_L g8781 ( 
.A(n_8489),
.Y(n_8781)
);

INVx3_ASAP7_75t_L g8782 ( 
.A(n_8420),
.Y(n_8782)
);

INVx1_ASAP7_75t_L g8783 ( 
.A(n_8302),
.Y(n_8783)
);

INVx1_ASAP7_75t_L g8784 ( 
.A(n_8303),
.Y(n_8784)
);

HB1xp67_ASAP7_75t_L g8785 ( 
.A(n_8527),
.Y(n_8785)
);

HB1xp67_ASAP7_75t_L g8786 ( 
.A(n_8540),
.Y(n_8786)
);

INVx1_ASAP7_75t_L g8787 ( 
.A(n_8304),
.Y(n_8787)
);

NOR2xp33_ASAP7_75t_SL g8788 ( 
.A(n_8092),
.B(n_5433),
.Y(n_8788)
);

INVx1_ASAP7_75t_L g8789 ( 
.A(n_8355),
.Y(n_8789)
);

AOI22xp5_ASAP7_75t_L g8790 ( 
.A1(n_8173),
.A2(n_5441),
.B1(n_5442),
.B2(n_5436),
.Y(n_8790)
);

CKINVDCx16_ASAP7_75t_R g8791 ( 
.A(n_8154),
.Y(n_8791)
);

INVx1_ASAP7_75t_L g8792 ( 
.A(n_8356),
.Y(n_8792)
);

INVx1_ASAP7_75t_L g8793 ( 
.A(n_8359),
.Y(n_8793)
);

NAND2xp5_ASAP7_75t_SL g8794 ( 
.A(n_8417),
.B(n_5443),
.Y(n_8794)
);

BUFx3_ASAP7_75t_L g8795 ( 
.A(n_8345),
.Y(n_8795)
);

INVx1_ASAP7_75t_SL g8796 ( 
.A(n_8442),
.Y(n_8796)
);

BUFx6f_ASAP7_75t_L g8797 ( 
.A(n_8312),
.Y(n_8797)
);

AND2x2_ASAP7_75t_L g8798 ( 
.A(n_8178),
.B(n_5444),
.Y(n_8798)
);

INVx2_ASAP7_75t_L g8799 ( 
.A(n_8349),
.Y(n_8799)
);

INVx2_ASAP7_75t_L g8800 ( 
.A(n_8353),
.Y(n_8800)
);

INVx2_ASAP7_75t_L g8801 ( 
.A(n_8354),
.Y(n_8801)
);

INVx1_ASAP7_75t_L g8802 ( 
.A(n_8360),
.Y(n_8802)
);

AOI22xp5_ASAP7_75t_L g8803 ( 
.A1(n_8173),
.A2(n_5448),
.B1(n_5449),
.B2(n_5446),
.Y(n_8803)
);

INVx1_ASAP7_75t_L g8804 ( 
.A(n_8362),
.Y(n_8804)
);

BUFx3_ASAP7_75t_L g8805 ( 
.A(n_8345),
.Y(n_8805)
);

INVx3_ASAP7_75t_L g8806 ( 
.A(n_8493),
.Y(n_8806)
);

INVx1_ASAP7_75t_L g8807 ( 
.A(n_8364),
.Y(n_8807)
);

INVx2_ASAP7_75t_L g8808 ( 
.A(n_8361),
.Y(n_8808)
);

AOI22xp5_ASAP7_75t_L g8809 ( 
.A1(n_8173),
.A2(n_5452),
.B1(n_5459),
.B2(n_5451),
.Y(n_8809)
);

INVx1_ASAP7_75t_L g8810 ( 
.A(n_8370),
.Y(n_8810)
);

INVx2_ASAP7_75t_L g8811 ( 
.A(n_8367),
.Y(n_8811)
);

INVx1_ASAP7_75t_L g8812 ( 
.A(n_8373),
.Y(n_8812)
);

INVx3_ASAP7_75t_L g8813 ( 
.A(n_8493),
.Y(n_8813)
);

INVx2_ASAP7_75t_L g8814 ( 
.A(n_8377),
.Y(n_8814)
);

BUFx6f_ASAP7_75t_L g8815 ( 
.A(n_8312),
.Y(n_8815)
);

INVx1_ASAP7_75t_L g8816 ( 
.A(n_8374),
.Y(n_8816)
);

INVx1_ASAP7_75t_L g8817 ( 
.A(n_8376),
.Y(n_8817)
);

INVx1_ASAP7_75t_L g8818 ( 
.A(n_8378),
.Y(n_8818)
);

AND2x4_ASAP7_75t_L g8819 ( 
.A(n_8457),
.B(n_5438),
.Y(n_8819)
);

INVx2_ASAP7_75t_L g8820 ( 
.A(n_8381),
.Y(n_8820)
);

INVx2_ASAP7_75t_L g8821 ( 
.A(n_8384),
.Y(n_8821)
);

INVx1_ASAP7_75t_L g8822 ( 
.A(n_8379),
.Y(n_8822)
);

INVx1_ASAP7_75t_L g8823 ( 
.A(n_8380),
.Y(n_8823)
);

INVx1_ASAP7_75t_L g8824 ( 
.A(n_8386),
.Y(n_8824)
);

BUFx6f_ASAP7_75t_L g8825 ( 
.A(n_8344),
.Y(n_8825)
);

INVx2_ASAP7_75t_L g8826 ( 
.A(n_8389),
.Y(n_8826)
);

AND2x4_ASAP7_75t_L g8827 ( 
.A(n_8270),
.B(n_5445),
.Y(n_8827)
);

NAND2xp5_ASAP7_75t_L g8828 ( 
.A(n_8110),
.B(n_5464),
.Y(n_8828)
);

INVx1_ASAP7_75t_L g8829 ( 
.A(n_8388),
.Y(n_8829)
);

AOI22xp5_ASAP7_75t_L g8830 ( 
.A1(n_8505),
.A2(n_5472),
.B1(n_5475),
.B2(n_5466),
.Y(n_8830)
);

INVx1_ASAP7_75t_L g8831 ( 
.A(n_8392),
.Y(n_8831)
);

HB1xp67_ASAP7_75t_L g8832 ( 
.A(n_8560),
.Y(n_8832)
);

BUFx2_ASAP7_75t_L g8833 ( 
.A(n_8193),
.Y(n_8833)
);

INVx2_ASAP7_75t_L g8834 ( 
.A(n_8391),
.Y(n_8834)
);

HB1xp67_ASAP7_75t_L g8835 ( 
.A(n_8564),
.Y(n_8835)
);

INVx1_ASAP7_75t_L g8836 ( 
.A(n_8394),
.Y(n_8836)
);

NAND2xp33_ASAP7_75t_L g8837 ( 
.A(n_8268),
.B(n_8272),
.Y(n_8837)
);

OAI22xp5_ASAP7_75t_SL g8838 ( 
.A1(n_8606),
.A2(n_5480),
.B1(n_5481),
.B2(n_5478),
.Y(n_8838)
);

INVx1_ASAP7_75t_L g8839 ( 
.A(n_8310),
.Y(n_8839)
);

AOI22xp5_ASAP7_75t_L g8840 ( 
.A1(n_8532),
.A2(n_5484),
.B1(n_5485),
.B2(n_5482),
.Y(n_8840)
);

INVx1_ASAP7_75t_L g8841 ( 
.A(n_8313),
.Y(n_8841)
);

BUFx2_ASAP7_75t_L g8842 ( 
.A(n_8223),
.Y(n_8842)
);

INVx1_ASAP7_75t_L g8843 ( 
.A(n_8321),
.Y(n_8843)
);

INVx1_ASAP7_75t_L g8844 ( 
.A(n_8325),
.Y(n_8844)
);

NAND2xp5_ASAP7_75t_L g8845 ( 
.A(n_8336),
.B(n_5489),
.Y(n_8845)
);

INVx1_ASAP7_75t_L g8846 ( 
.A(n_8338),
.Y(n_8846)
);

INVx1_ASAP7_75t_L g8847 ( 
.A(n_8114),
.Y(n_8847)
);

INVx1_ASAP7_75t_L g8848 ( 
.A(n_8116),
.Y(n_8848)
);

INVxp67_ASAP7_75t_L g8849 ( 
.A(n_8194),
.Y(n_8849)
);

INVx1_ASAP7_75t_L g8850 ( 
.A(n_8119),
.Y(n_8850)
);

INVx3_ASAP7_75t_L g8851 ( 
.A(n_8512),
.Y(n_8851)
);

BUFx6f_ASAP7_75t_L g8852 ( 
.A(n_8344),
.Y(n_8852)
);

BUFx6f_ASAP7_75t_L g8853 ( 
.A(n_8512),
.Y(n_8853)
);

NAND2xp5_ASAP7_75t_L g8854 ( 
.A(n_8340),
.B(n_5490),
.Y(n_8854)
);

NAND2xp33_ASAP7_75t_SL g8855 ( 
.A(n_8557),
.B(n_5492),
.Y(n_8855)
);

AOI22xp5_ASAP7_75t_L g8856 ( 
.A1(n_8282),
.A2(n_5494),
.B1(n_5496),
.B2(n_5493),
.Y(n_8856)
);

INVx1_ASAP7_75t_L g8857 ( 
.A(n_8126),
.Y(n_8857)
);

NAND2xp5_ASAP7_75t_L g8858 ( 
.A(n_8288),
.B(n_5497),
.Y(n_8858)
);

NAND2xp5_ASAP7_75t_SL g8859 ( 
.A(n_8419),
.B(n_5498),
.Y(n_8859)
);

INVx1_ASAP7_75t_L g8860 ( 
.A(n_8127),
.Y(n_8860)
);

INVxp67_ASAP7_75t_L g8861 ( 
.A(n_8197),
.Y(n_8861)
);

INVx2_ASAP7_75t_L g8862 ( 
.A(n_8134),
.Y(n_8862)
);

INVx2_ASAP7_75t_L g8863 ( 
.A(n_8137),
.Y(n_8863)
);

INVx1_ASAP7_75t_L g8864 ( 
.A(n_8221),
.Y(n_8864)
);

INVx2_ASAP7_75t_L g8865 ( 
.A(n_8227),
.Y(n_8865)
);

NAND2xp5_ASAP7_75t_L g8866 ( 
.A(n_8435),
.B(n_5500),
.Y(n_8866)
);

BUFx3_ASAP7_75t_L g8867 ( 
.A(n_8317),
.Y(n_8867)
);

OAI22xp5_ASAP7_75t_SL g8868 ( 
.A1(n_8609),
.A2(n_5505),
.B1(n_5508),
.B2(n_5502),
.Y(n_8868)
);

INVx2_ASAP7_75t_L g8869 ( 
.A(n_8234),
.Y(n_8869)
);

INVx2_ASAP7_75t_L g8870 ( 
.A(n_8237),
.Y(n_8870)
);

INVx2_ASAP7_75t_L g8871 ( 
.A(n_8243),
.Y(n_8871)
);

NAND2xp5_ASAP7_75t_L g8872 ( 
.A(n_8073),
.B(n_5509),
.Y(n_8872)
);

OAI22xp5_ASAP7_75t_SL g8873 ( 
.A1(n_8570),
.A2(n_5513),
.B1(n_5514),
.B2(n_5512),
.Y(n_8873)
);

BUFx6f_ASAP7_75t_L g8874 ( 
.A(n_8536),
.Y(n_8874)
);

BUFx6f_ASAP7_75t_L g8875 ( 
.A(n_8536),
.Y(n_8875)
);

INVx1_ASAP7_75t_L g8876 ( 
.A(n_8337),
.Y(n_8876)
);

INVx2_ASAP7_75t_L g8877 ( 
.A(n_8339),
.Y(n_8877)
);

AND2x2_ASAP7_75t_L g8878 ( 
.A(n_8208),
.B(n_5518),
.Y(n_8878)
);

AND2x2_ASAP7_75t_L g8879 ( 
.A(n_8295),
.B(n_5522),
.Y(n_8879)
);

HB1xp67_ASAP7_75t_L g8880 ( 
.A(n_8444),
.Y(n_8880)
);

INVxp67_ASAP7_75t_L g8881 ( 
.A(n_8135),
.Y(n_8881)
);

INVx1_ASAP7_75t_L g8882 ( 
.A(n_8521),
.Y(n_8882)
);

INVx1_ASAP7_75t_SL g8883 ( 
.A(n_8450),
.Y(n_8883)
);

NAND2xp5_ASAP7_75t_L g8884 ( 
.A(n_8363),
.B(n_5528),
.Y(n_8884)
);

INVx3_ASAP7_75t_L g8885 ( 
.A(n_8563),
.Y(n_8885)
);

INVx1_ASAP7_75t_L g8886 ( 
.A(n_8523),
.Y(n_8886)
);

HB1xp67_ASAP7_75t_L g8887 ( 
.A(n_8451),
.Y(n_8887)
);

INVx2_ASAP7_75t_L g8888 ( 
.A(n_8529),
.Y(n_8888)
);

INVx1_ASAP7_75t_L g8889 ( 
.A(n_8414),
.Y(n_8889)
);

AOI22xp5_ASAP7_75t_L g8890 ( 
.A1(n_8496),
.A2(n_5532),
.B1(n_5534),
.B2(n_5531),
.Y(n_8890)
);

HB1xp67_ASAP7_75t_L g8891 ( 
.A(n_8453),
.Y(n_8891)
);

INVx1_ASAP7_75t_L g8892 ( 
.A(n_8422),
.Y(n_8892)
);

BUFx6f_ASAP7_75t_L g8893 ( 
.A(n_8563),
.Y(n_8893)
);

INVx3_ASAP7_75t_L g8894 ( 
.A(n_8584),
.Y(n_8894)
);

HB1xp67_ASAP7_75t_L g8895 ( 
.A(n_8458),
.Y(n_8895)
);

INVx1_ASAP7_75t_L g8896 ( 
.A(n_8449),
.Y(n_8896)
);

INVx1_ASAP7_75t_L g8897 ( 
.A(n_8484),
.Y(n_8897)
);

NOR2xp33_ASAP7_75t_L g8898 ( 
.A(n_8318),
.B(n_5535),
.Y(n_8898)
);

INVx8_ASAP7_75t_L g8899 ( 
.A(n_8213),
.Y(n_8899)
);

INVx1_ASAP7_75t_L g8900 ( 
.A(n_8486),
.Y(n_8900)
);

INVx2_ASAP7_75t_L g8901 ( 
.A(n_8148),
.Y(n_8901)
);

INVx3_ASAP7_75t_L g8902 ( 
.A(n_8584),
.Y(n_8902)
);

INVx1_ASAP7_75t_L g8903 ( 
.A(n_8498),
.Y(n_8903)
);

INVx1_ASAP7_75t_L g8904 ( 
.A(n_8506),
.Y(n_8904)
);

NAND2xp33_ASAP7_75t_SL g8905 ( 
.A(n_8569),
.B(n_5537),
.Y(n_8905)
);

INVx1_ASAP7_75t_SL g8906 ( 
.A(n_8461),
.Y(n_8906)
);

INVx2_ASAP7_75t_L g8907 ( 
.A(n_8163),
.Y(n_8907)
);

INVx2_ASAP7_75t_L g8908 ( 
.A(n_8165),
.Y(n_8908)
);

INVx1_ASAP7_75t_L g8909 ( 
.A(n_8507),
.Y(n_8909)
);

HB1xp67_ASAP7_75t_L g8910 ( 
.A(n_8094),
.Y(n_8910)
);

INVx1_ASAP7_75t_SL g8911 ( 
.A(n_8462),
.Y(n_8911)
);

NAND2xp5_ASAP7_75t_L g8912 ( 
.A(n_8369),
.B(n_5543),
.Y(n_8912)
);

OAI22xp5_ASAP7_75t_SL g8913 ( 
.A1(n_8539),
.A2(n_5545),
.B1(n_5550),
.B2(n_5544),
.Y(n_8913)
);

HB1xp67_ASAP7_75t_L g8914 ( 
.A(n_8108),
.Y(n_8914)
);

INVx1_ASAP7_75t_L g8915 ( 
.A(n_8508),
.Y(n_8915)
);

AND2x4_ASAP7_75t_L g8916 ( 
.A(n_8332),
.B(n_5453),
.Y(n_8916)
);

AND2x2_ASAP7_75t_L g8917 ( 
.A(n_8343),
.B(n_5553),
.Y(n_8917)
);

NOR2xp33_ASAP7_75t_SL g8918 ( 
.A(n_8096),
.B(n_5554),
.Y(n_8918)
);

INVx1_ASAP7_75t_L g8919 ( 
.A(n_8513),
.Y(n_8919)
);

INVx1_ASAP7_75t_L g8920 ( 
.A(n_8519),
.Y(n_8920)
);

INVx2_ASAP7_75t_L g8921 ( 
.A(n_8184),
.Y(n_8921)
);

INVx1_ASAP7_75t_L g8922 ( 
.A(n_8520),
.Y(n_8922)
);

CKINVDCx8_ASAP7_75t_R g8923 ( 
.A(n_8098),
.Y(n_8923)
);

INVx2_ASAP7_75t_L g8924 ( 
.A(n_8074),
.Y(n_8924)
);

HB1xp67_ASAP7_75t_L g8925 ( 
.A(n_8200),
.Y(n_8925)
);

INVx2_ASAP7_75t_L g8926 ( 
.A(n_8279),
.Y(n_8926)
);

INVx1_ASAP7_75t_L g8927 ( 
.A(n_8415),
.Y(n_8927)
);

INVx2_ASAP7_75t_L g8928 ( 
.A(n_8427),
.Y(n_8928)
);

INVx1_ASAP7_75t_L g8929 ( 
.A(n_8429),
.Y(n_8929)
);

INVx2_ASAP7_75t_L g8930 ( 
.A(n_8432),
.Y(n_8930)
);

INVx2_ASAP7_75t_L g8931 ( 
.A(n_8434),
.Y(n_8931)
);

INVx1_ASAP7_75t_L g8932 ( 
.A(n_8437),
.Y(n_8932)
);

INVx1_ASAP7_75t_L g8933 ( 
.A(n_8438),
.Y(n_8933)
);

NAND2xp5_ASAP7_75t_SL g8934 ( 
.A(n_8421),
.B(n_5557),
.Y(n_8934)
);

AND2x2_ASAP7_75t_L g8935 ( 
.A(n_8348),
.B(n_5558),
.Y(n_8935)
);

BUFx6f_ASAP7_75t_L g8936 ( 
.A(n_8592),
.Y(n_8936)
);

INVx1_ASAP7_75t_L g8937 ( 
.A(n_8441),
.Y(n_8937)
);

INVx1_ASAP7_75t_L g8938 ( 
.A(n_8446),
.Y(n_8938)
);

INVx1_ASAP7_75t_L g8939 ( 
.A(n_8459),
.Y(n_8939)
);

INVx2_ASAP7_75t_L g8940 ( 
.A(n_8492),
.Y(n_8940)
);

NAND2xp5_ASAP7_75t_L g8941 ( 
.A(n_8405),
.B(n_5559),
.Y(n_8941)
);

BUFx6f_ASAP7_75t_L g8942 ( 
.A(n_8592),
.Y(n_8942)
);

OAI22xp5_ASAP7_75t_SL g8943 ( 
.A1(n_8543),
.A2(n_8608),
.B1(n_8618),
.B2(n_8613),
.Y(n_8943)
);

AOI22xp5_ASAP7_75t_L g8944 ( 
.A1(n_8499),
.A2(n_5563),
.B1(n_5564),
.B2(n_5562),
.Y(n_8944)
);

NAND2xp5_ASAP7_75t_SL g8945 ( 
.A(n_8423),
.B(n_5565),
.Y(n_8945)
);

INVx1_ASAP7_75t_L g8946 ( 
.A(n_8342),
.Y(n_8946)
);

OAI22xp5_ASAP7_75t_SL g8947 ( 
.A1(n_8276),
.A2(n_5570),
.B1(n_5571),
.B2(n_5569),
.Y(n_8947)
);

CKINVDCx20_ASAP7_75t_R g8948 ( 
.A(n_8130),
.Y(n_8948)
);

HB1xp67_ASAP7_75t_L g8949 ( 
.A(n_8504),
.Y(n_8949)
);

INVx1_ASAP7_75t_L g8950 ( 
.A(n_8400),
.Y(n_8950)
);

NAND2xp5_ASAP7_75t_L g8951 ( 
.A(n_8418),
.B(n_5576),
.Y(n_8951)
);

OAI22xp5_ASAP7_75t_SL g8952 ( 
.A1(n_8491),
.A2(n_5579),
.B1(n_5582),
.B2(n_5578),
.Y(n_8952)
);

NOR2xp33_ASAP7_75t_L g8953 ( 
.A(n_8465),
.B(n_8447),
.Y(n_8953)
);

AOI22xp5_ASAP7_75t_L g8954 ( 
.A1(n_8329),
.A2(n_5585),
.B1(n_5586),
.B2(n_5584),
.Y(n_8954)
);

BUFx8_ASAP7_75t_L g8955 ( 
.A(n_8291),
.Y(n_8955)
);

BUFx6f_ASAP7_75t_L g8956 ( 
.A(n_8599),
.Y(n_8956)
);

OAI22xp5_ASAP7_75t_SL g8957 ( 
.A1(n_8531),
.A2(n_5591),
.B1(n_5593),
.B2(n_5589),
.Y(n_8957)
);

INVx1_ASAP7_75t_L g8958 ( 
.A(n_8403),
.Y(n_8958)
);

INVx2_ASAP7_75t_L g8959 ( 
.A(n_8500),
.Y(n_8959)
);

INVx1_ASAP7_75t_SL g8960 ( 
.A(n_8371),
.Y(n_8960)
);

BUFx2_ASAP7_75t_L g8961 ( 
.A(n_8411),
.Y(n_8961)
);

BUFx6f_ASAP7_75t_L g8962 ( 
.A(n_8599),
.Y(n_8962)
);

BUFx6f_ASAP7_75t_L g8963 ( 
.A(n_8478),
.Y(n_8963)
);

INVx2_ASAP7_75t_L g8964 ( 
.A(n_8503),
.Y(n_8964)
);

INVx1_ASAP7_75t_L g8965 ( 
.A(n_8407),
.Y(n_8965)
);

INVx3_ASAP7_75t_L g8966 ( 
.A(n_8382),
.Y(n_8966)
);

AOI22xp5_ASAP7_75t_L g8967 ( 
.A1(n_8549),
.A2(n_5600),
.B1(n_5601),
.B2(n_5599),
.Y(n_8967)
);

INVx1_ASAP7_75t_SL g8968 ( 
.A(n_8260),
.Y(n_8968)
);

INVx1_ASAP7_75t_L g8969 ( 
.A(n_8488),
.Y(n_8969)
);

BUFx6f_ASAP7_75t_L g8970 ( 
.A(n_8177),
.Y(n_8970)
);

OAI22xp5_ASAP7_75t_SL g8971 ( 
.A1(n_8578),
.A2(n_5603),
.B1(n_5606),
.B2(n_5602),
.Y(n_8971)
);

AND2x2_ASAP7_75t_L g8972 ( 
.A(n_8366),
.B(n_5608),
.Y(n_8972)
);

INVx1_ASAP7_75t_L g8973 ( 
.A(n_8490),
.Y(n_8973)
);

INVx8_ASAP7_75t_L g8974 ( 
.A(n_8213),
.Y(n_8974)
);

AND2x2_ASAP7_75t_L g8975 ( 
.A(n_8456),
.B(n_8269),
.Y(n_8975)
);

INVx3_ASAP7_75t_L g8976 ( 
.A(n_8436),
.Y(n_8976)
);

HB1xp67_ASAP7_75t_L g8977 ( 
.A(n_8576),
.Y(n_8977)
);

INVx1_ASAP7_75t_L g8978 ( 
.A(n_8553),
.Y(n_8978)
);

INVx1_ASAP7_75t_L g8979 ( 
.A(n_8554),
.Y(n_8979)
);

BUFx6f_ASAP7_75t_L g8980 ( 
.A(n_8191),
.Y(n_8980)
);

INVx8_ASAP7_75t_L g8981 ( 
.A(n_8213),
.Y(n_8981)
);

INVx3_ASAP7_75t_L g8982 ( 
.A(n_8439),
.Y(n_8982)
);

INVx6_ASAP7_75t_L g8983 ( 
.A(n_8231),
.Y(n_8983)
);

AND2x2_ASAP7_75t_L g8984 ( 
.A(n_8607),
.B(n_5611),
.Y(n_8984)
);

NAND2xp5_ASAP7_75t_L g8985 ( 
.A(n_8218),
.B(n_5614),
.Y(n_8985)
);

INVx1_ASAP7_75t_L g8986 ( 
.A(n_8274),
.Y(n_8986)
);

BUFx6f_ASAP7_75t_L g8987 ( 
.A(n_8207),
.Y(n_8987)
);

HB1xp67_ASAP7_75t_L g8988 ( 
.A(n_8600),
.Y(n_8988)
);

INVx3_ASAP7_75t_L g8989 ( 
.A(n_8454),
.Y(n_8989)
);

INVx1_ASAP7_75t_L g8990 ( 
.A(n_8258),
.Y(n_8990)
);

INVx1_ASAP7_75t_L g8991 ( 
.A(n_8300),
.Y(n_8991)
);

INVx1_ASAP7_75t_L g8992 ( 
.A(n_8311),
.Y(n_8992)
);

INVx2_ASAP7_75t_L g8993 ( 
.A(n_8192),
.Y(n_8993)
);

NOR2xp33_ASAP7_75t_L g8994 ( 
.A(n_8413),
.B(n_5615),
.Y(n_8994)
);

INVx1_ASAP7_75t_L g8995 ( 
.A(n_8526),
.Y(n_8995)
);

AOI22xp5_ASAP7_75t_L g8996 ( 
.A1(n_8542),
.A2(n_5619),
.B1(n_5624),
.B2(n_5618),
.Y(n_8996)
);

AND2x4_ASAP7_75t_L g8997 ( 
.A(n_8466),
.B(n_5454),
.Y(n_8997)
);

INVx1_ASAP7_75t_L g8998 ( 
.A(n_8518),
.Y(n_8998)
);

INVx1_ASAP7_75t_L g8999 ( 
.A(n_8244),
.Y(n_8999)
);

INVx8_ASAP7_75t_L g9000 ( 
.A(n_8198),
.Y(n_9000)
);

BUFx4f_ASAP7_75t_L g9001 ( 
.A(n_8157),
.Y(n_9001)
);

INVx1_ASAP7_75t_SL g9002 ( 
.A(n_8289),
.Y(n_9002)
);

INVxp67_ASAP7_75t_L g9003 ( 
.A(n_8581),
.Y(n_9003)
);

OA21x2_ASAP7_75t_L g9004 ( 
.A1(n_8620),
.A2(n_5460),
.B(n_5456),
.Y(n_9004)
);

HB1xp67_ASAP7_75t_L g9005 ( 
.A(n_8566),
.Y(n_9005)
);

INVx1_ASAP7_75t_L g9006 ( 
.A(n_8327),
.Y(n_9006)
);

AND2x2_ASAP7_75t_L g9007 ( 
.A(n_8275),
.B(n_5625),
.Y(n_9007)
);

INVx1_ASAP7_75t_L g9008 ( 
.A(n_8078),
.Y(n_9008)
);

NAND2xp5_ASAP7_75t_SL g9009 ( 
.A(n_8284),
.B(n_8286),
.Y(n_9009)
);

INVx1_ASAP7_75t_L g9010 ( 
.A(n_8085),
.Y(n_9010)
);

INVx2_ASAP7_75t_L g9011 ( 
.A(n_8610),
.Y(n_9011)
);

INVx1_ASAP7_75t_L g9012 ( 
.A(n_8249),
.Y(n_9012)
);

INVx1_ASAP7_75t_L g9013 ( 
.A(n_8281),
.Y(n_9013)
);

INVx1_ASAP7_75t_L g9014 ( 
.A(n_8097),
.Y(n_9014)
);

INVx2_ASAP7_75t_L g9015 ( 
.A(n_8619),
.Y(n_9015)
);

INVx1_ASAP7_75t_L g9016 ( 
.A(n_8105),
.Y(n_9016)
);

INVxp67_ASAP7_75t_L g9017 ( 
.A(n_8155),
.Y(n_9017)
);

INVx3_ASAP7_75t_L g9018 ( 
.A(n_8481),
.Y(n_9018)
);

INVx2_ASAP7_75t_L g9019 ( 
.A(n_8619),
.Y(n_9019)
);

OA22x2_ASAP7_75t_L g9020 ( 
.A1(n_8555),
.A2(n_5628),
.B1(n_5629),
.B2(n_5626),
.Y(n_9020)
);

INVx3_ASAP7_75t_SL g9021 ( 
.A(n_8203),
.Y(n_9021)
);

INVx3_ASAP7_75t_L g9022 ( 
.A(n_8575),
.Y(n_9022)
);

BUFx6f_ASAP7_75t_L g9023 ( 
.A(n_8216),
.Y(n_9023)
);

INVx1_ASAP7_75t_L g9024 ( 
.A(n_8158),
.Y(n_9024)
);

INVx3_ASAP7_75t_L g9025 ( 
.A(n_8585),
.Y(n_9025)
);

NAND2xp5_ASAP7_75t_L g9026 ( 
.A(n_8568),
.B(n_8455),
.Y(n_9026)
);

INVx1_ASAP7_75t_L g9027 ( 
.A(n_8161),
.Y(n_9027)
);

INVx1_ASAP7_75t_L g9028 ( 
.A(n_8168),
.Y(n_9028)
);

NAND2xp5_ASAP7_75t_SL g9029 ( 
.A(n_8287),
.B(n_8290),
.Y(n_9029)
);

AND2x6_ASAP7_75t_L g9030 ( 
.A(n_8357),
.B(n_5462),
.Y(n_9030)
);

NAND2xp5_ASAP7_75t_L g9031 ( 
.A(n_8460),
.B(n_5630),
.Y(n_9031)
);

INVx1_ASAP7_75t_L g9032 ( 
.A(n_8175),
.Y(n_9032)
);

INVx1_ASAP7_75t_L g9033 ( 
.A(n_8202),
.Y(n_9033)
);

INVx2_ASAP7_75t_L g9034 ( 
.A(n_8160),
.Y(n_9034)
);

NAND2xp5_ASAP7_75t_L g9035 ( 
.A(n_8495),
.B(n_5631),
.Y(n_9035)
);

INVx1_ASAP7_75t_L g9036 ( 
.A(n_8611),
.Y(n_9036)
);

INVx3_ASAP7_75t_L g9037 ( 
.A(n_8255),
.Y(n_9037)
);

BUFx2_ASAP7_75t_L g9038 ( 
.A(n_8305),
.Y(n_9038)
);

HB1xp67_ASAP7_75t_L g9039 ( 
.A(n_8524),
.Y(n_9039)
);

AOI22xp5_ASAP7_75t_L g9040 ( 
.A1(n_8583),
.A2(n_5635),
.B1(n_5637),
.B2(n_5633),
.Y(n_9040)
);

AOI22xp5_ASAP7_75t_L g9041 ( 
.A1(n_8603),
.A2(n_5642),
.B1(n_5644),
.B2(n_5638),
.Y(n_9041)
);

NAND2xp33_ASAP7_75t_SL g9042 ( 
.A(n_8426),
.B(n_5646),
.Y(n_9042)
);

INVx2_ASAP7_75t_L g9043 ( 
.A(n_8409),
.Y(n_9043)
);

INVx3_ASAP7_75t_L g9044 ( 
.A(n_8263),
.Y(n_9044)
);

INVx1_ASAP7_75t_L g9045 ( 
.A(n_8614),
.Y(n_9045)
);

HB1xp67_ASAP7_75t_L g9046 ( 
.A(n_8574),
.Y(n_9046)
);

INVx1_ASAP7_75t_L g9047 ( 
.A(n_8579),
.Y(n_9047)
);

INVx2_ASAP7_75t_L g9048 ( 
.A(n_8535),
.Y(n_9048)
);

INVx2_ASAP7_75t_L g9049 ( 
.A(n_8544),
.Y(n_9049)
);

INVx1_ASAP7_75t_L g9050 ( 
.A(n_8601),
.Y(n_9050)
);

AOI22xp5_ASAP7_75t_L g9051 ( 
.A1(n_8572),
.A2(n_5655),
.B1(n_5657),
.B2(n_5652),
.Y(n_9051)
);

BUFx6f_ASAP7_75t_L g9052 ( 
.A(n_8297),
.Y(n_9052)
);

INVx1_ASAP7_75t_L g9053 ( 
.A(n_8408),
.Y(n_9053)
);

INVx1_ASAP7_75t_SL g9054 ( 
.A(n_8350),
.Y(n_9054)
);

CKINVDCx5p33_ASAP7_75t_R g9055 ( 
.A(n_8099),
.Y(n_9055)
);

AND2x2_ASAP7_75t_L g9056 ( 
.A(n_8547),
.B(n_5660),
.Y(n_9056)
);

INVx2_ASAP7_75t_L g9057 ( 
.A(n_8412),
.Y(n_9057)
);

INVx1_ASAP7_75t_L g9058 ( 
.A(n_8463),
.Y(n_9058)
);

BUFx6f_ASAP7_75t_L g9059 ( 
.A(n_8233),
.Y(n_9059)
);

HB1xp67_ASAP7_75t_L g9060 ( 
.A(n_8209),
.Y(n_9060)
);

INVx2_ASAP7_75t_L g9061 ( 
.A(n_8445),
.Y(n_9061)
);

INVx2_ASAP7_75t_L g9062 ( 
.A(n_8468),
.Y(n_9062)
);

INVx2_ASAP7_75t_L g9063 ( 
.A(n_8474),
.Y(n_9063)
);

BUFx6f_ASAP7_75t_L g9064 ( 
.A(n_8593),
.Y(n_9064)
);

INVx1_ASAP7_75t_L g9065 ( 
.A(n_8477),
.Y(n_9065)
);

NAND2xp5_ASAP7_75t_SL g9066 ( 
.A(n_8443),
.B(n_5663),
.Y(n_9066)
);

INVx2_ASAP7_75t_L g9067 ( 
.A(n_8479),
.Y(n_9067)
);

OAI22xp5_ASAP7_75t_SL g9068 ( 
.A1(n_8533),
.A2(n_8467),
.B1(n_8525),
.B2(n_8515),
.Y(n_9068)
);

INVx2_ASAP7_75t_L g9069 ( 
.A(n_8485),
.Y(n_9069)
);

NAND2xp5_ASAP7_75t_L g9070 ( 
.A(n_8517),
.B(n_5666),
.Y(n_9070)
);

NAND2xp5_ASAP7_75t_L g9071 ( 
.A(n_8559),
.B(n_5669),
.Y(n_9071)
);

INVx3_ASAP7_75t_L g9072 ( 
.A(n_8567),
.Y(n_9072)
);

NAND2xp5_ASAP7_75t_SL g9073 ( 
.A(n_8433),
.B(n_8330),
.Y(n_9073)
);

INVx1_ASAP7_75t_L g9074 ( 
.A(n_8551),
.Y(n_9074)
);

OAI22xp5_ASAP7_75t_L g9075 ( 
.A1(n_8588),
.A2(n_5674),
.B1(n_5675),
.B2(n_5670),
.Y(n_9075)
);

INVx3_ASAP7_75t_L g9076 ( 
.A(n_8595),
.Y(n_9076)
);

INVx1_ASAP7_75t_L g9077 ( 
.A(n_8558),
.Y(n_9077)
);

INVx3_ASAP7_75t_L g9078 ( 
.A(n_8561),
.Y(n_9078)
);

INVx1_ASAP7_75t_L g9079 ( 
.A(n_8480),
.Y(n_9079)
);

INVx1_ASAP7_75t_L g9080 ( 
.A(n_8612),
.Y(n_9080)
);

INVx1_ASAP7_75t_L g9081 ( 
.A(n_8577),
.Y(n_9081)
);

INVx1_ASAP7_75t_L g9082 ( 
.A(n_8582),
.Y(n_9082)
);

AOI22xp5_ASAP7_75t_L g9083 ( 
.A1(n_8541),
.A2(n_5678),
.B1(n_5680),
.B2(n_5677),
.Y(n_9083)
);

INVx1_ASAP7_75t_L g9084 ( 
.A(n_8586),
.Y(n_9084)
);

INVx3_ASAP7_75t_L g9085 ( 
.A(n_8589),
.Y(n_9085)
);

INVx2_ASAP7_75t_L g9086 ( 
.A(n_8590),
.Y(n_9086)
);

INVxp67_ASAP7_75t_L g9087 ( 
.A(n_8476),
.Y(n_9087)
);

BUFx6f_ASAP7_75t_L g9088 ( 
.A(n_8157),
.Y(n_9088)
);

INVxp67_ASAP7_75t_L g9089 ( 
.A(n_8587),
.Y(n_9089)
);

INVx2_ASAP7_75t_L g9090 ( 
.A(n_8591),
.Y(n_9090)
);

INVx1_ASAP7_75t_L g9091 ( 
.A(n_8597),
.Y(n_9091)
);

INVx1_ASAP7_75t_L g9092 ( 
.A(n_8598),
.Y(n_9092)
);

INVx2_ASAP7_75t_L g9093 ( 
.A(n_8424),
.Y(n_9093)
);

INVx2_ASAP7_75t_L g9094 ( 
.A(n_8406),
.Y(n_9094)
);

INVx1_ASAP7_75t_L g9095 ( 
.A(n_8615),
.Y(n_9095)
);

BUFx2_ASAP7_75t_L g9096 ( 
.A(n_8214),
.Y(n_9096)
);

NAND2xp5_ASAP7_75t_SL g9097 ( 
.A(n_8341),
.B(n_5682),
.Y(n_9097)
);

HB1xp67_ASAP7_75t_L g9098 ( 
.A(n_8210),
.Y(n_9098)
);

INVx5_ASAP7_75t_L g9099 ( 
.A(n_8546),
.Y(n_9099)
);

INVx3_ASAP7_75t_L g9100 ( 
.A(n_8217),
.Y(n_9100)
);

AND2x4_ASAP7_75t_L g9101 ( 
.A(n_8594),
.B(n_5465),
.Y(n_9101)
);

BUFx6f_ASAP7_75t_L g9102 ( 
.A(n_8222),
.Y(n_9102)
);

AND2x2_ASAP7_75t_L g9103 ( 
.A(n_8538),
.B(n_5683),
.Y(n_9103)
);

AND2x4_ASAP7_75t_L g9104 ( 
.A(n_8228),
.B(n_5469),
.Y(n_9104)
);

NAND2xp5_ASAP7_75t_SL g9105 ( 
.A(n_8605),
.B(n_5684),
.Y(n_9105)
);

CKINVDCx20_ASAP7_75t_R g9106 ( 
.A(n_8128),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_8472),
.Y(n_9107)
);

INVx1_ASAP7_75t_L g9108 ( 
.A(n_8509),
.Y(n_9108)
);

BUFx3_ASAP7_75t_SL g9109 ( 
.A(n_8385),
.Y(n_9109)
);

BUFx6f_ASAP7_75t_L g9110 ( 
.A(n_8320),
.Y(n_9110)
);

INVx1_ASAP7_75t_L g9111 ( 
.A(n_8516),
.Y(n_9111)
);

INVx1_ASAP7_75t_L g9112 ( 
.A(n_8522),
.Y(n_9112)
);

BUFx6f_ASAP7_75t_L g9113 ( 
.A(n_8395),
.Y(n_9113)
);

INVx2_ASAP7_75t_L g9114 ( 
.A(n_8346),
.Y(n_9114)
);

INVx1_ASAP7_75t_L g9115 ( 
.A(n_8571),
.Y(n_9115)
);

INVx1_ASAP7_75t_L g9116 ( 
.A(n_8571),
.Y(n_9116)
);

INVx2_ASAP7_75t_L g9117 ( 
.A(n_8346),
.Y(n_9117)
);

INVx1_ASAP7_75t_L g9118 ( 
.A(n_8571),
.Y(n_9118)
);

INVx1_ASAP7_75t_L g9119 ( 
.A(n_8346),
.Y(n_9119)
);

OAI22xp5_ASAP7_75t_SL g9120 ( 
.A1(n_8528),
.A2(n_5689),
.B1(n_5696),
.B2(n_5687),
.Y(n_9120)
);

NAND2xp5_ASAP7_75t_L g9121 ( 
.A(n_8239),
.B(n_5699),
.Y(n_9121)
);

INVx2_ASAP7_75t_L g9122 ( 
.A(n_8316),
.Y(n_9122)
);

INVx2_ASAP7_75t_L g9123 ( 
.A(n_8104),
.Y(n_9123)
);

XOR2xp5_ASAP7_75t_L g9124 ( 
.A(n_8247),
.B(n_4334),
.Y(n_9124)
);

INVxp67_ASAP7_75t_L g9125 ( 
.A(n_8375),
.Y(n_9125)
);

INVx1_ASAP7_75t_L g9126 ( 
.A(n_8324),
.Y(n_9126)
);

BUFx6f_ASAP7_75t_L g9127 ( 
.A(n_8546),
.Y(n_9127)
);

INVx1_ASAP7_75t_L g9128 ( 
.A(n_8334),
.Y(n_9128)
);

NAND2xp5_ASAP7_75t_L g9129 ( 
.A(n_8293),
.B(n_5700),
.Y(n_9129)
);

INVx1_ASAP7_75t_L g9130 ( 
.A(n_8473),
.Y(n_9130)
);

INVx1_ASAP7_75t_L g9131 ( 
.A(n_8292),
.Y(n_9131)
);

INVx2_ASAP7_75t_L g9132 ( 
.A(n_8307),
.Y(n_9132)
);

NAND2xp5_ASAP7_75t_L g9133 ( 
.A(n_8322),
.B(n_5702),
.Y(n_9133)
);

INVx1_ASAP7_75t_L g9134 ( 
.A(n_8106),
.Y(n_9134)
);

INVx2_ASAP7_75t_L g9135 ( 
.A(n_8075),
.Y(n_9135)
);

INVx1_ASAP7_75t_L g9136 ( 
.A(n_8404),
.Y(n_9136)
);

BUFx2_ASAP7_75t_L g9137 ( 
.A(n_8252),
.Y(n_9137)
);

INVx1_ASAP7_75t_L g9138 ( 
.A(n_8314),
.Y(n_9138)
);

INVx1_ASAP7_75t_L g9139 ( 
.A(n_8315),
.Y(n_9139)
);

INVx2_ASAP7_75t_L g9140 ( 
.A(n_8238),
.Y(n_9140)
);

NAND2xp33_ASAP7_75t_SL g9141 ( 
.A(n_8428),
.B(n_5704),
.Y(n_9141)
);

INVx3_ASAP7_75t_SL g9142 ( 
.A(n_8102),
.Y(n_9142)
);

NAND2xp33_ASAP7_75t_SL g9143 ( 
.A(n_8430),
.B(n_8552),
.Y(n_9143)
);

NAND2xp5_ASAP7_75t_SL g9144 ( 
.A(n_8139),
.B(n_5705),
.Y(n_9144)
);

AND2x4_ASAP7_75t_L g9145 ( 
.A(n_8189),
.B(n_5470),
.Y(n_9145)
);

BUFx6f_ASAP7_75t_L g9146 ( 
.A(n_8107),
.Y(n_9146)
);

INVx3_ASAP7_75t_L g9147 ( 
.A(n_8250),
.Y(n_9147)
);

INVx3_ASAP7_75t_L g9148 ( 
.A(n_8251),
.Y(n_9148)
);

INVx2_ASAP7_75t_L g9149 ( 
.A(n_8254),
.Y(n_9149)
);

INVx1_ASAP7_75t_L g9150 ( 
.A(n_8471),
.Y(n_9150)
);

INVx1_ASAP7_75t_L g9151 ( 
.A(n_8257),
.Y(n_9151)
);

INVx1_ASAP7_75t_L g9152 ( 
.A(n_8494),
.Y(n_9152)
);

AND2x2_ASAP7_75t_L g9153 ( 
.A(n_8118),
.B(n_5706),
.Y(n_9153)
);

INVx1_ASAP7_75t_L g9154 ( 
.A(n_8121),
.Y(n_9154)
);

INVx1_ASAP7_75t_L g9155 ( 
.A(n_8125),
.Y(n_9155)
);

INVx1_ASAP7_75t_L g9156 ( 
.A(n_8129),
.Y(n_9156)
);

OR2x2_ASAP7_75t_L g9157 ( 
.A(n_8132),
.B(n_5708),
.Y(n_9157)
);

OAI22xp5_ASAP7_75t_SL g9158 ( 
.A1(n_8431),
.A2(n_5712),
.B1(n_5713),
.B2(n_5710),
.Y(n_9158)
);

NOR2xp33_ASAP7_75t_L g9159 ( 
.A(n_8133),
.B(n_5715),
.Y(n_9159)
);

INVx1_ASAP7_75t_L g9160 ( 
.A(n_8136),
.Y(n_9160)
);

XOR2xp5_ASAP7_75t_L g9161 ( 
.A(n_8057),
.B(n_4335),
.Y(n_9161)
);

INVx1_ASAP7_75t_L g9162 ( 
.A(n_8440),
.Y(n_9162)
);

NAND2xp5_ASAP7_75t_L g9163 ( 
.A(n_8550),
.B(n_5717),
.Y(n_9163)
);

INVx1_ASAP7_75t_L g9164 ( 
.A(n_8470),
.Y(n_9164)
);

HB1xp67_ASAP7_75t_L g9165 ( 
.A(n_8530),
.Y(n_9165)
);

INVx2_ASAP7_75t_L g9166 ( 
.A(n_8323),
.Y(n_9166)
);

INVx1_ASAP7_75t_L g9167 ( 
.A(n_8298),
.Y(n_9167)
);

BUFx6f_ASAP7_75t_L g9168 ( 
.A(n_8230),
.Y(n_9168)
);

NAND2xp5_ASAP7_75t_L g9169 ( 
.A(n_8170),
.B(n_5718),
.Y(n_9169)
);

INVx1_ASAP7_75t_L g9170 ( 
.A(n_8176),
.Y(n_9170)
);

BUFx6f_ASAP7_75t_SL g9171 ( 
.A(n_8331),
.Y(n_9171)
);

INVx1_ASAP7_75t_L g9172 ( 
.A(n_8179),
.Y(n_9172)
);

INVx1_ASAP7_75t_L g9173 ( 
.A(n_8141),
.Y(n_9173)
);

NAND2xp5_ASAP7_75t_L g9174 ( 
.A(n_8145),
.B(n_5719),
.Y(n_9174)
);

NAND2xp33_ASAP7_75t_SL g9175 ( 
.A(n_8185),
.B(n_8188),
.Y(n_9175)
);

BUFx4f_ASAP7_75t_L g9176 ( 
.A(n_9102),
.Y(n_9176)
);

NAND2xp33_ASAP7_75t_L g9177 ( 
.A(n_8738),
.B(n_8062),
.Y(n_9177)
);

BUFx6f_ASAP7_75t_L g9178 ( 
.A(n_8629),
.Y(n_9178)
);

INVx3_ASAP7_75t_L g9179 ( 
.A(n_9102),
.Y(n_9179)
);

BUFx3_ASAP7_75t_L g9180 ( 
.A(n_9000),
.Y(n_9180)
);

BUFx3_ASAP7_75t_L g9181 ( 
.A(n_9000),
.Y(n_9181)
);

NOR2xp33_ASAP7_75t_L g9182 ( 
.A(n_8659),
.B(n_8066),
.Y(n_9182)
);

INVx2_ASAP7_75t_L g9183 ( 
.A(n_8888),
.Y(n_9183)
);

OAI22xp33_ASAP7_75t_L g9184 ( 
.A1(n_8669),
.A2(n_8152),
.B1(n_8162),
.B2(n_8146),
.Y(n_9184)
);

INVx1_ASAP7_75t_L g9185 ( 
.A(n_8621),
.Y(n_9185)
);

INVx2_ASAP7_75t_SL g9186 ( 
.A(n_8689),
.Y(n_9186)
);

AND2x4_ASAP7_75t_L g9187 ( 
.A(n_8644),
.B(n_8159),
.Y(n_9187)
);

INVx1_ASAP7_75t_L g9188 ( 
.A(n_8625),
.Y(n_9188)
);

INVx5_ASAP7_75t_L g9189 ( 
.A(n_9146),
.Y(n_9189)
);

AND2x4_ASAP7_75t_L g9190 ( 
.A(n_8867),
.B(n_8067),
.Y(n_9190)
);

INVx1_ASAP7_75t_L g9191 ( 
.A(n_8628),
.Y(n_9191)
);

INVx1_ASAP7_75t_L g9192 ( 
.A(n_8630),
.Y(n_9192)
);

OR2x6_ASAP7_75t_L g9193 ( 
.A(n_9059),
.B(n_8164),
.Y(n_9193)
);

INVx2_ASAP7_75t_SL g9194 ( 
.A(n_8853),
.Y(n_9194)
);

BUFx6f_ASAP7_75t_L g9195 ( 
.A(n_8629),
.Y(n_9195)
);

NAND2xp5_ASAP7_75t_L g9196 ( 
.A(n_8627),
.B(n_5721),
.Y(n_9196)
);

INVx2_ASAP7_75t_L g9197 ( 
.A(n_8720),
.Y(n_9197)
);

BUFx2_ASAP7_75t_L g9198 ( 
.A(n_8961),
.Y(n_9198)
);

INVx1_ASAP7_75t_L g9199 ( 
.A(n_8642),
.Y(n_9199)
);

INVx2_ASAP7_75t_L g9200 ( 
.A(n_8732),
.Y(n_9200)
);

INVx1_ASAP7_75t_L g9201 ( 
.A(n_8646),
.Y(n_9201)
);

INVx1_ASAP7_75t_L g9202 ( 
.A(n_8648),
.Y(n_9202)
);

INVx2_ASAP7_75t_L g9203 ( 
.A(n_8742),
.Y(n_9203)
);

CKINVDCx5p33_ASAP7_75t_R g9204 ( 
.A(n_9055),
.Y(n_9204)
);

NAND3xp33_ASAP7_75t_L g9205 ( 
.A(n_8994),
.B(n_8452),
.C(n_8082),
.Y(n_9205)
);

INVx4_ASAP7_75t_L g9206 ( 
.A(n_9059),
.Y(n_9206)
);

INVx2_ASAP7_75t_L g9207 ( 
.A(n_8756),
.Y(n_9207)
);

INVx2_ASAP7_75t_L g9208 ( 
.A(n_8765),
.Y(n_9208)
);

AND2x2_ASAP7_75t_L g9209 ( 
.A(n_8622),
.B(n_8172),
.Y(n_9209)
);

NOR2xp33_ASAP7_75t_L g9210 ( 
.A(n_9012),
.B(n_8358),
.Y(n_9210)
);

CKINVDCx5p33_ASAP7_75t_R g9211 ( 
.A(n_8923),
.Y(n_9211)
);

NOR2xp33_ASAP7_75t_L g9212 ( 
.A(n_9013),
.B(n_8352),
.Y(n_9212)
);

INVx1_ASAP7_75t_L g9213 ( 
.A(n_8649),
.Y(n_9213)
);

INVxp67_ASAP7_75t_SL g9214 ( 
.A(n_8681),
.Y(n_9214)
);

INVx1_ASAP7_75t_L g9215 ( 
.A(n_8654),
.Y(n_9215)
);

INVx1_ASAP7_75t_L g9216 ( 
.A(n_8657),
.Y(n_9216)
);

INVx1_ASAP7_75t_L g9217 ( 
.A(n_8658),
.Y(n_9217)
);

NAND2xp5_ASAP7_75t_SL g9218 ( 
.A(n_8975),
.B(n_5723),
.Y(n_9218)
);

NOR2xp33_ASAP7_75t_L g9219 ( 
.A(n_8953),
.B(n_5724),
.Y(n_9219)
);

NAND2xp33_ASAP7_75t_SL g9220 ( 
.A(n_9142),
.B(n_8399),
.Y(n_9220)
);

AND2x4_ASAP7_75t_L g9221 ( 
.A(n_8795),
.B(n_8402),
.Y(n_9221)
);

INVx2_ASAP7_75t_L g9222 ( 
.A(n_8769),
.Y(n_9222)
);

NAND2xp5_ASAP7_75t_L g9223 ( 
.A(n_9014),
.B(n_5725),
.Y(n_9223)
);

BUFx3_ASAP7_75t_L g9224 ( 
.A(n_8805),
.Y(n_9224)
);

INVx1_ASAP7_75t_L g9225 ( 
.A(n_8661),
.Y(n_9225)
);

AND2x6_ASAP7_75t_L g9226 ( 
.A(n_9146),
.B(n_5471),
.Y(n_9226)
);

NAND2xp5_ASAP7_75t_SL g9227 ( 
.A(n_9016),
.B(n_5726),
.Y(n_9227)
);

INVx1_ASAP7_75t_SL g9228 ( 
.A(n_8691),
.Y(n_9228)
);

AND2x6_ASAP7_75t_L g9229 ( 
.A(n_9154),
.B(n_5473),
.Y(n_9229)
);

AND2x4_ASAP7_75t_L g9230 ( 
.A(n_9100),
.B(n_5487),
.Y(n_9230)
);

BUFx6f_ASAP7_75t_L g9231 ( 
.A(n_8651),
.Y(n_9231)
);

INVxp67_ASAP7_75t_SL g9232 ( 
.A(n_8702),
.Y(n_9232)
);

BUFx2_ASAP7_75t_L g9233 ( 
.A(n_8635),
.Y(n_9233)
);

INVx1_ASAP7_75t_L g9234 ( 
.A(n_8663),
.Y(n_9234)
);

NAND2xp5_ASAP7_75t_L g9235 ( 
.A(n_9024),
.B(n_5727),
.Y(n_9235)
);

NAND2xp5_ASAP7_75t_L g9236 ( 
.A(n_9027),
.B(n_5729),
.Y(n_9236)
);

AND2x2_ASAP7_75t_L g9237 ( 
.A(n_9056),
.B(n_5730),
.Y(n_9237)
);

AOI22xp33_ASAP7_75t_L g9238 ( 
.A1(n_8704),
.A2(n_5787),
.B1(n_5846),
.B2(n_5784),
.Y(n_9238)
);

INVx1_ASAP7_75t_L g9239 ( 
.A(n_8665),
.Y(n_9239)
);

AND2x4_ASAP7_75t_L g9240 ( 
.A(n_8963),
.B(n_5510),
.Y(n_9240)
);

AND2x2_ASAP7_75t_L g9241 ( 
.A(n_8984),
.B(n_5733),
.Y(n_9241)
);

OAI21xp33_ASAP7_75t_L g9242 ( 
.A1(n_8840),
.A2(n_5735),
.B(n_5734),
.Y(n_9242)
);

INVx1_ASAP7_75t_L g9243 ( 
.A(n_8666),
.Y(n_9243)
);

INVx1_ASAP7_75t_L g9244 ( 
.A(n_8667),
.Y(n_9244)
);

INVx2_ASAP7_75t_L g9245 ( 
.A(n_8774),
.Y(n_9245)
);

AND2x2_ASAP7_75t_L g9246 ( 
.A(n_8717),
.B(n_5736),
.Y(n_9246)
);

INVx3_ASAP7_75t_L g9247 ( 
.A(n_8853),
.Y(n_9247)
);

BUFx3_ASAP7_75t_L g9248 ( 
.A(n_8874),
.Y(n_9248)
);

CKINVDCx5p33_ASAP7_75t_R g9249 ( 
.A(n_8727),
.Y(n_9249)
);

NAND2xp5_ASAP7_75t_L g9250 ( 
.A(n_9028),
.B(n_5737),
.Y(n_9250)
);

AND2x6_ASAP7_75t_L g9251 ( 
.A(n_9155),
.B(n_5511),
.Y(n_9251)
);

INVx1_ASAP7_75t_L g9252 ( 
.A(n_8673),
.Y(n_9252)
);

INVx2_ASAP7_75t_L g9253 ( 
.A(n_8776),
.Y(n_9253)
);

NOR2x1p5_ASAP7_75t_L g9254 ( 
.A(n_9088),
.B(n_5740),
.Y(n_9254)
);

INVx3_ASAP7_75t_L g9255 ( 
.A(n_8874),
.Y(n_9255)
);

AND2x4_ASAP7_75t_L g9256 ( 
.A(n_8963),
.B(n_5524),
.Y(n_9256)
);

AND2x2_ASAP7_75t_L g9257 ( 
.A(n_8798),
.B(n_5746),
.Y(n_9257)
);

AOI21x1_ASAP7_75t_L g9258 ( 
.A1(n_8632),
.A2(n_5530),
.B(n_5525),
.Y(n_9258)
);

NAND2xp5_ASAP7_75t_L g9259 ( 
.A(n_9032),
.B(n_5747),
.Y(n_9259)
);

INVx2_ASAP7_75t_L g9260 ( 
.A(n_8780),
.Y(n_9260)
);

BUFx6f_ASAP7_75t_L g9261 ( 
.A(n_8651),
.Y(n_9261)
);

AND2x2_ASAP7_75t_L g9262 ( 
.A(n_8878),
.B(n_5752),
.Y(n_9262)
);

CKINVDCx5p33_ASAP7_75t_R g9263 ( 
.A(n_8638),
.Y(n_9263)
);

NOR2xp33_ASAP7_75t_L g9264 ( 
.A(n_9033),
.B(n_9017),
.Y(n_9264)
);

INVx2_ASAP7_75t_L g9265 ( 
.A(n_8940),
.Y(n_9265)
);

BUFx4f_ASAP7_75t_L g9266 ( 
.A(n_9021),
.Y(n_9266)
);

BUFx3_ASAP7_75t_L g9267 ( 
.A(n_8875),
.Y(n_9267)
);

BUFx6f_ASAP7_75t_L g9268 ( 
.A(n_8664),
.Y(n_9268)
);

OR2x6_ASAP7_75t_L g9269 ( 
.A(n_9088),
.B(n_8899),
.Y(n_9269)
);

INVx1_ASAP7_75t_L g9270 ( 
.A(n_8677),
.Y(n_9270)
);

INVx4_ASAP7_75t_SL g9271 ( 
.A(n_8983),
.Y(n_9271)
);

NAND2xp5_ASAP7_75t_L g9272 ( 
.A(n_9026),
.B(n_9008),
.Y(n_9272)
);

NAND3xp33_ASAP7_75t_SL g9273 ( 
.A(n_8716),
.B(n_5757),
.C(n_5753),
.Y(n_9273)
);

INVxp67_ASAP7_75t_SL g9274 ( 
.A(n_8706),
.Y(n_9274)
);

INVx1_ASAP7_75t_SL g9275 ( 
.A(n_8749),
.Y(n_9275)
);

NOR2xp33_ASAP7_75t_L g9276 ( 
.A(n_9010),
.B(n_5761),
.Y(n_9276)
);

NAND2xp5_ASAP7_75t_L g9277 ( 
.A(n_8641),
.B(n_5763),
.Y(n_9277)
);

INVx2_ASAP7_75t_L g9278 ( 
.A(n_8959),
.Y(n_9278)
);

INVx2_ASAP7_75t_L g9279 ( 
.A(n_8964),
.Y(n_9279)
);

NAND2xp5_ASAP7_75t_SL g9280 ( 
.A(n_9125),
.B(n_5766),
.Y(n_9280)
);

INVx2_ASAP7_75t_L g9281 ( 
.A(n_9011),
.Y(n_9281)
);

INVx1_ASAP7_75t_SL g9282 ( 
.A(n_8796),
.Y(n_9282)
);

INVx4_ASAP7_75t_L g9283 ( 
.A(n_8875),
.Y(n_9283)
);

BUFx6f_ASAP7_75t_L g9284 ( 
.A(n_8664),
.Y(n_9284)
);

INVx1_ASAP7_75t_L g9285 ( 
.A(n_8682),
.Y(n_9285)
);

INVx2_ASAP7_75t_L g9286 ( 
.A(n_8623),
.Y(n_9286)
);

AOI22xp33_ASAP7_75t_L g9287 ( 
.A1(n_9006),
.A2(n_5915),
.B1(n_5922),
.B2(n_5864),
.Y(n_9287)
);

AOI22x1_ASAP7_75t_L g9288 ( 
.A1(n_9134),
.A2(n_5546),
.B1(n_5548),
.B2(n_5540),
.Y(n_9288)
);

AND2x4_ASAP7_75t_L g9289 ( 
.A(n_9047),
.B(n_9050),
.Y(n_9289)
);

NAND2xp5_ASAP7_75t_L g9290 ( 
.A(n_8828),
.B(n_8750),
.Y(n_9290)
);

INVx4_ASAP7_75t_L g9291 ( 
.A(n_8893),
.Y(n_9291)
);

BUFx6f_ASAP7_75t_L g9292 ( 
.A(n_8670),
.Y(n_9292)
);

INVx1_ASAP7_75t_L g9293 ( 
.A(n_8683),
.Y(n_9293)
);

INVx2_ASAP7_75t_L g9294 ( 
.A(n_8624),
.Y(n_9294)
);

INVx2_ASAP7_75t_L g9295 ( 
.A(n_8626),
.Y(n_9295)
);

INVx2_ASAP7_75t_L g9296 ( 
.A(n_8631),
.Y(n_9296)
);

NAND2xp33_ASAP7_75t_L g9297 ( 
.A(n_9136),
.B(n_5767),
.Y(n_9297)
);

INVx1_ASAP7_75t_L g9298 ( 
.A(n_8690),
.Y(n_9298)
);

INVx2_ASAP7_75t_L g9299 ( 
.A(n_8656),
.Y(n_9299)
);

INVx1_ASAP7_75t_L g9300 ( 
.A(n_8693),
.Y(n_9300)
);

INVx5_ASAP7_75t_L g9301 ( 
.A(n_9168),
.Y(n_9301)
);

INVx2_ASAP7_75t_L g9302 ( 
.A(n_8662),
.Y(n_9302)
);

BUFx2_ASAP7_75t_L g9303 ( 
.A(n_8747),
.Y(n_9303)
);

NAND2xp5_ASAP7_75t_L g9304 ( 
.A(n_8845),
.B(n_5769),
.Y(n_9304)
);

AND2x2_ASAP7_75t_L g9305 ( 
.A(n_8917),
.B(n_5772),
.Y(n_9305)
);

BUFx10_ASAP7_75t_L g9306 ( 
.A(n_8758),
.Y(n_9306)
);

BUFx2_ASAP7_75t_L g9307 ( 
.A(n_8645),
.Y(n_9307)
);

NAND2xp5_ASAP7_75t_L g9308 ( 
.A(n_8854),
.B(n_5774),
.Y(n_9308)
);

NAND2xp5_ASAP7_75t_L g9309 ( 
.A(n_8872),
.B(n_8884),
.Y(n_9309)
);

INVx1_ASAP7_75t_SL g9310 ( 
.A(n_8883),
.Y(n_9310)
);

NOR2xp33_ASAP7_75t_SL g9311 ( 
.A(n_8640),
.B(n_5776),
.Y(n_9311)
);

NOR2xp33_ASAP7_75t_L g9312 ( 
.A(n_9089),
.B(n_5778),
.Y(n_9312)
);

BUFx3_ASAP7_75t_L g9313 ( 
.A(n_8893),
.Y(n_9313)
);

NAND2xp5_ASAP7_75t_L g9314 ( 
.A(n_8912),
.B(n_5782),
.Y(n_9314)
);

INVx2_ASAP7_75t_L g9315 ( 
.A(n_8668),
.Y(n_9315)
);

INVx1_ASAP7_75t_L g9316 ( 
.A(n_8695),
.Y(n_9316)
);

INVx2_ASAP7_75t_L g9317 ( 
.A(n_8676),
.Y(n_9317)
);

BUFx3_ASAP7_75t_L g9318 ( 
.A(n_8936),
.Y(n_9318)
);

INVx4_ASAP7_75t_L g9319 ( 
.A(n_8936),
.Y(n_9319)
);

NAND2xp5_ASAP7_75t_SL g9320 ( 
.A(n_8650),
.B(n_8906),
.Y(n_9320)
);

INVx1_ASAP7_75t_L g9321 ( 
.A(n_8698),
.Y(n_9321)
);

NAND2xp5_ASAP7_75t_L g9322 ( 
.A(n_8941),
.B(n_5785),
.Y(n_9322)
);

INVx1_ASAP7_75t_L g9323 ( 
.A(n_8700),
.Y(n_9323)
);

AND2x2_ASAP7_75t_L g9324 ( 
.A(n_8680),
.B(n_5790),
.Y(n_9324)
);

AND2x2_ASAP7_75t_L g9325 ( 
.A(n_8935),
.B(n_5794),
.Y(n_9325)
);

NAND2xp5_ASAP7_75t_L g9326 ( 
.A(n_8951),
.B(n_5795),
.Y(n_9326)
);

BUFx4f_ASAP7_75t_L g9327 ( 
.A(n_9168),
.Y(n_9327)
);

INVx2_ASAP7_75t_L g9328 ( 
.A(n_8684),
.Y(n_9328)
);

AND2x4_ASAP7_75t_SL g9329 ( 
.A(n_9060),
.B(n_5556),
.Y(n_9329)
);

INVx2_ASAP7_75t_L g9330 ( 
.A(n_8705),
.Y(n_9330)
);

INVx1_ASAP7_75t_L g9331 ( 
.A(n_8703),
.Y(n_9331)
);

INVx3_ASAP7_75t_L g9332 ( 
.A(n_8942),
.Y(n_9332)
);

NAND2xp5_ASAP7_75t_SL g9333 ( 
.A(n_8911),
.B(n_5796),
.Y(n_9333)
);

BUFx2_ASAP7_75t_L g9334 ( 
.A(n_8768),
.Y(n_9334)
);

BUFx10_ASAP7_75t_L g9335 ( 
.A(n_8721),
.Y(n_9335)
);

INVx2_ASAP7_75t_L g9336 ( 
.A(n_8708),
.Y(n_9336)
);

NAND2xp5_ASAP7_75t_L g9337 ( 
.A(n_8866),
.B(n_5798),
.Y(n_9337)
);

INVx1_ASAP7_75t_L g9338 ( 
.A(n_8710),
.Y(n_9338)
);

NAND2xp5_ASAP7_75t_SL g9339 ( 
.A(n_8995),
.B(n_8949),
.Y(n_9339)
);

NOR2xp33_ASAP7_75t_L g9340 ( 
.A(n_8699),
.B(n_5799),
.Y(n_9340)
);

BUFx6f_ASAP7_75t_L g9341 ( 
.A(n_8670),
.Y(n_9341)
);

BUFx6f_ASAP7_75t_L g9342 ( 
.A(n_8671),
.Y(n_9342)
);

INVx1_ASAP7_75t_L g9343 ( 
.A(n_8714),
.Y(n_9343)
);

INVx2_ASAP7_75t_L g9344 ( 
.A(n_8713),
.Y(n_9344)
);

NAND2xp5_ASAP7_75t_L g9345 ( 
.A(n_8858),
.B(n_5800),
.Y(n_9345)
);

INVx4_ASAP7_75t_L g9346 ( 
.A(n_8942),
.Y(n_9346)
);

NOR2xp33_ASAP7_75t_SL g9347 ( 
.A(n_9001),
.B(n_5801),
.Y(n_9347)
);

INVx1_ASAP7_75t_L g9348 ( 
.A(n_8723),
.Y(n_9348)
);

INVx3_ASAP7_75t_L g9349 ( 
.A(n_8956),
.Y(n_9349)
);

AO22x2_ASAP7_75t_L g9350 ( 
.A1(n_9109),
.A2(n_9116),
.B1(n_9118),
.B2(n_9115),
.Y(n_9350)
);

AND2x2_ASAP7_75t_L g9351 ( 
.A(n_8972),
.B(n_5803),
.Y(n_9351)
);

BUFx6f_ASAP7_75t_L g9352 ( 
.A(n_8671),
.Y(n_9352)
);

OR2x2_ASAP7_75t_L g9353 ( 
.A(n_8960),
.B(n_5804),
.Y(n_9353)
);

NAND2xp5_ASAP7_75t_SL g9354 ( 
.A(n_9147),
.B(n_5808),
.Y(n_9354)
);

INVx4_ASAP7_75t_L g9355 ( 
.A(n_8956),
.Y(n_9355)
);

INVx2_ASAP7_75t_L g9356 ( 
.A(n_8799),
.Y(n_9356)
);

AOI22xp33_ASAP7_75t_L g9357 ( 
.A1(n_8674),
.A2(n_5986),
.B1(n_5993),
.B2(n_5956),
.Y(n_9357)
);

INVx2_ASAP7_75t_L g9358 ( 
.A(n_8800),
.Y(n_9358)
);

INVx1_ASAP7_75t_L g9359 ( 
.A(n_8724),
.Y(n_9359)
);

INVx1_ASAP7_75t_L g9360 ( 
.A(n_8725),
.Y(n_9360)
);

NOR2xp33_ASAP7_75t_L g9361 ( 
.A(n_8943),
.B(n_5809),
.Y(n_9361)
);

INVx1_ASAP7_75t_L g9362 ( 
.A(n_8729),
.Y(n_9362)
);

INVx1_ASAP7_75t_L g9363 ( 
.A(n_8730),
.Y(n_9363)
);

NAND2xp33_ASAP7_75t_L g9364 ( 
.A(n_8674),
.B(n_5811),
.Y(n_9364)
);

BUFx6f_ASAP7_75t_L g9365 ( 
.A(n_8687),
.Y(n_9365)
);

INVx4_ASAP7_75t_L g9366 ( 
.A(n_8962),
.Y(n_9366)
);

NAND2xp5_ASAP7_75t_L g9367 ( 
.A(n_9031),
.B(n_9035),
.Y(n_9367)
);

BUFx3_ASAP7_75t_L g9368 ( 
.A(n_8962),
.Y(n_9368)
);

INVx4_ASAP7_75t_L g9369 ( 
.A(n_8687),
.Y(n_9369)
);

INVx2_ASAP7_75t_L g9370 ( 
.A(n_8801),
.Y(n_9370)
);

BUFx6f_ASAP7_75t_L g9371 ( 
.A(n_8697),
.Y(n_9371)
);

BUFx10_ASAP7_75t_L g9372 ( 
.A(n_9171),
.Y(n_9372)
);

OR2x2_ASAP7_75t_L g9373 ( 
.A(n_8968),
.B(n_5815),
.Y(n_9373)
);

NOR2xp33_ASAP7_75t_L g9374 ( 
.A(n_8849),
.B(n_8861),
.Y(n_9374)
);

INVx2_ASAP7_75t_L g9375 ( 
.A(n_8808),
.Y(n_9375)
);

INVx2_ASAP7_75t_L g9376 ( 
.A(n_8811),
.Y(n_9376)
);

INVx1_ASAP7_75t_L g9377 ( 
.A(n_8734),
.Y(n_9377)
);

INVx4_ASAP7_75t_L g9378 ( 
.A(n_8697),
.Y(n_9378)
);

INVx4_ASAP7_75t_L g9379 ( 
.A(n_8709),
.Y(n_9379)
);

INVx1_ASAP7_75t_L g9380 ( 
.A(n_8735),
.Y(n_9380)
);

NAND2xp5_ASAP7_75t_L g9381 ( 
.A(n_8736),
.B(n_5817),
.Y(n_9381)
);

INVx4_ASAP7_75t_L g9382 ( 
.A(n_8709),
.Y(n_9382)
);

NAND2xp5_ASAP7_75t_L g9383 ( 
.A(n_8737),
.B(n_5818),
.Y(n_9383)
);

NAND2xp5_ASAP7_75t_SL g9384 ( 
.A(n_9148),
.B(n_9132),
.Y(n_9384)
);

INVx2_ASAP7_75t_L g9385 ( 
.A(n_8814),
.Y(n_9385)
);

INVx2_ASAP7_75t_L g9386 ( 
.A(n_8820),
.Y(n_9386)
);

AND2x6_ASAP7_75t_L g9387 ( 
.A(n_9156),
.B(n_5560),
.Y(n_9387)
);

AND2x4_ASAP7_75t_L g9388 ( 
.A(n_9110),
.B(n_5561),
.Y(n_9388)
);

INVx4_ASAP7_75t_L g9389 ( 
.A(n_8731),
.Y(n_9389)
);

INVx2_ASAP7_75t_L g9390 ( 
.A(n_8821),
.Y(n_9390)
);

INVx2_ASAP7_75t_L g9391 ( 
.A(n_8826),
.Y(n_9391)
);

INVx4_ASAP7_75t_L g9392 ( 
.A(n_8731),
.Y(n_9392)
);

BUFx3_ASAP7_75t_L g9393 ( 
.A(n_8733),
.Y(n_9393)
);

INVx2_ASAP7_75t_L g9394 ( 
.A(n_8834),
.Y(n_9394)
);

INVx1_ASAP7_75t_L g9395 ( 
.A(n_8741),
.Y(n_9395)
);

BUFx3_ASAP7_75t_L g9396 ( 
.A(n_8733),
.Y(n_9396)
);

INVx1_ASAP7_75t_L g9397 ( 
.A(n_8743),
.Y(n_9397)
);

INVx2_ASAP7_75t_SL g9398 ( 
.A(n_8757),
.Y(n_9398)
);

BUFx6f_ASAP7_75t_L g9399 ( 
.A(n_8757),
.Y(n_9399)
);

AND2x2_ASAP7_75t_L g9400 ( 
.A(n_8898),
.B(n_5819),
.Y(n_9400)
);

INVx1_ASAP7_75t_L g9401 ( 
.A(n_8744),
.Y(n_9401)
);

BUFx10_ASAP7_75t_L g9402 ( 
.A(n_9159),
.Y(n_9402)
);

INVx1_ASAP7_75t_L g9403 ( 
.A(n_8746),
.Y(n_9403)
);

AND2x4_ASAP7_75t_L g9404 ( 
.A(n_9110),
.B(n_5566),
.Y(n_9404)
);

AND2x2_ASAP7_75t_L g9405 ( 
.A(n_9007),
.B(n_5827),
.Y(n_9405)
);

INVx5_ASAP7_75t_L g9406 ( 
.A(n_8762),
.Y(n_9406)
);

INVx1_ASAP7_75t_L g9407 ( 
.A(n_8752),
.Y(n_9407)
);

INVx2_ASAP7_75t_SL g9408 ( 
.A(n_8762),
.Y(n_9408)
);

BUFx6f_ASAP7_75t_L g9409 ( 
.A(n_8797),
.Y(n_9409)
);

INVx4_ASAP7_75t_L g9410 ( 
.A(n_8797),
.Y(n_9410)
);

INVx2_ASAP7_75t_L g9411 ( 
.A(n_8862),
.Y(n_9411)
);

INVx8_ASAP7_75t_L g9412 ( 
.A(n_8815),
.Y(n_9412)
);

INVx1_ASAP7_75t_L g9413 ( 
.A(n_8753),
.Y(n_9413)
);

NAND2xp5_ASAP7_75t_L g9414 ( 
.A(n_8755),
.B(n_5828),
.Y(n_9414)
);

OR2x2_ASAP7_75t_L g9415 ( 
.A(n_9002),
.B(n_5836),
.Y(n_9415)
);

NAND2xp33_ASAP7_75t_L g9416 ( 
.A(n_8674),
.B(n_5837),
.Y(n_9416)
);

AO22x2_ASAP7_75t_L g9417 ( 
.A1(n_9107),
.A2(n_5568),
.B1(n_5572),
.B2(n_5567),
.Y(n_9417)
);

AND2x4_ASAP7_75t_L g9418 ( 
.A(n_9113),
.B(n_5573),
.Y(n_9418)
);

INVx1_ASAP7_75t_L g9419 ( 
.A(n_8759),
.Y(n_9419)
);

AND2x2_ASAP7_75t_L g9420 ( 
.A(n_9153),
.B(n_5840),
.Y(n_9420)
);

NAND2xp5_ASAP7_75t_L g9421 ( 
.A(n_8760),
.B(n_5841),
.Y(n_9421)
);

AO22x1_ASAP7_75t_L g9422 ( 
.A1(n_9138),
.A2(n_5844),
.B1(n_5845),
.B2(n_5843),
.Y(n_9422)
);

BUFx2_ASAP7_75t_L g9423 ( 
.A(n_8833),
.Y(n_9423)
);

INVx1_ASAP7_75t_L g9424 ( 
.A(n_8764),
.Y(n_9424)
);

BUFx6f_ASAP7_75t_L g9425 ( 
.A(n_8815),
.Y(n_9425)
);

NOR2x1p5_ASAP7_75t_L g9426 ( 
.A(n_9064),
.B(n_5850),
.Y(n_9426)
);

INVx1_ASAP7_75t_L g9427 ( 
.A(n_8770),
.Y(n_9427)
);

INVx1_ASAP7_75t_L g9428 ( 
.A(n_8771),
.Y(n_9428)
);

INVx1_ASAP7_75t_L g9429 ( 
.A(n_8772),
.Y(n_9429)
);

NOR2xp33_ASAP7_75t_L g9430 ( 
.A(n_8688),
.B(n_5851),
.Y(n_9430)
);

INVx2_ASAP7_75t_L g9431 ( 
.A(n_8863),
.Y(n_9431)
);

AND2x6_ASAP7_75t_L g9432 ( 
.A(n_9160),
.B(n_5575),
.Y(n_9432)
);

NOR2xp33_ASAP7_75t_SL g9433 ( 
.A(n_9098),
.B(n_5857),
.Y(n_9433)
);

NAND2xp5_ASAP7_75t_L g9434 ( 
.A(n_8773),
.B(n_5858),
.Y(n_9434)
);

CKINVDCx5p33_ASAP7_75t_R g9435 ( 
.A(n_9106),
.Y(n_9435)
);

INVx2_ASAP7_75t_L g9436 ( 
.A(n_8865),
.Y(n_9436)
);

AND2x2_ASAP7_75t_L g9437 ( 
.A(n_8675),
.B(n_5859),
.Y(n_9437)
);

BUFx2_ASAP7_75t_L g9438 ( 
.A(n_8842),
.Y(n_9438)
);

INVx3_ASAP7_75t_L g9439 ( 
.A(n_8825),
.Y(n_9439)
);

INVx1_ASAP7_75t_L g9440 ( 
.A(n_8775),
.Y(n_9440)
);

INVx2_ASAP7_75t_SL g9441 ( 
.A(n_8825),
.Y(n_9441)
);

AND2x2_ASAP7_75t_L g9442 ( 
.A(n_8881),
.B(n_5860),
.Y(n_9442)
);

INVx1_ASAP7_75t_L g9443 ( 
.A(n_8777),
.Y(n_9443)
);

NOR2xp33_ASAP7_75t_L g9444 ( 
.A(n_8781),
.B(n_5861),
.Y(n_9444)
);

BUFx2_ASAP7_75t_L g9445 ( 
.A(n_9038),
.Y(n_9445)
);

OR2x6_ASAP7_75t_L g9446 ( 
.A(n_8899),
.B(n_5581),
.Y(n_9446)
);

AND2x4_ASAP7_75t_L g9447 ( 
.A(n_9113),
.B(n_5583),
.Y(n_9447)
);

NAND2xp5_ASAP7_75t_L g9448 ( 
.A(n_8783),
.B(n_5863),
.Y(n_9448)
);

AND2x4_ASAP7_75t_L g9449 ( 
.A(n_8637),
.B(n_5592),
.Y(n_9449)
);

INVx2_ASAP7_75t_L g9450 ( 
.A(n_8869),
.Y(n_9450)
);

BUFx3_ASAP7_75t_L g9451 ( 
.A(n_8852),
.Y(n_9451)
);

BUFx3_ASAP7_75t_L g9452 ( 
.A(n_8852),
.Y(n_9452)
);

INVx1_ASAP7_75t_L g9453 ( 
.A(n_8784),
.Y(n_9453)
);

INVx1_ASAP7_75t_L g9454 ( 
.A(n_8787),
.Y(n_9454)
);

NOR2xp33_ASAP7_75t_L g9455 ( 
.A(n_8715),
.B(n_8722),
.Y(n_9455)
);

BUFx2_ASAP7_75t_L g9456 ( 
.A(n_8754),
.Y(n_9456)
);

AND2x2_ASAP7_75t_L g9457 ( 
.A(n_8879),
.B(n_5867),
.Y(n_9457)
);

INVx1_ASAP7_75t_L g9458 ( 
.A(n_8789),
.Y(n_9458)
);

NAND3xp33_ASAP7_75t_L g9459 ( 
.A(n_8719),
.B(n_5871),
.C(n_5869),
.Y(n_9459)
);

INVxp67_ASAP7_75t_SL g9460 ( 
.A(n_8785),
.Y(n_9460)
);

AND2x6_ASAP7_75t_L g9461 ( 
.A(n_9108),
.B(n_5594),
.Y(n_9461)
);

INVx4_ASAP7_75t_L g9462 ( 
.A(n_9064),
.Y(n_9462)
);

INVx1_ASAP7_75t_L g9463 ( 
.A(n_8792),
.Y(n_9463)
);

AND2x4_ASAP7_75t_L g9464 ( 
.A(n_8728),
.B(n_5607),
.Y(n_9464)
);

AND2x4_ASAP7_75t_L g9465 ( 
.A(n_8779),
.B(n_5609),
.Y(n_9465)
);

INVx2_ASAP7_75t_L g9466 ( 
.A(n_8870),
.Y(n_9466)
);

INVx4_ASAP7_75t_L g9467 ( 
.A(n_8970),
.Y(n_9467)
);

NAND2xp5_ASAP7_75t_L g9468 ( 
.A(n_8633),
.B(n_5878),
.Y(n_9468)
);

CKINVDCx5p33_ASAP7_75t_R g9469 ( 
.A(n_8948),
.Y(n_9469)
);

BUFx3_ASAP7_75t_L g9470 ( 
.A(n_9137),
.Y(n_9470)
);

AND2x2_ASAP7_75t_L g9471 ( 
.A(n_9103),
.B(n_5879),
.Y(n_9471)
);

INVx3_ASAP7_75t_L g9472 ( 
.A(n_8970),
.Y(n_9472)
);

NAND2xp5_ASAP7_75t_L g9473 ( 
.A(n_8985),
.B(n_5880),
.Y(n_9473)
);

NAND2xp5_ASAP7_75t_L g9474 ( 
.A(n_8678),
.B(n_5882),
.Y(n_9474)
);

AND2x2_ASAP7_75t_L g9475 ( 
.A(n_8880),
.B(n_5884),
.Y(n_9475)
);

BUFx2_ASAP7_75t_L g9476 ( 
.A(n_8887),
.Y(n_9476)
);

INVx1_ASAP7_75t_L g9477 ( 
.A(n_8793),
.Y(n_9477)
);

AND2x4_ASAP7_75t_L g9478 ( 
.A(n_8782),
.B(n_5610),
.Y(n_9478)
);

OR2x2_ASAP7_75t_L g9479 ( 
.A(n_8696),
.B(n_5885),
.Y(n_9479)
);

INVx1_ASAP7_75t_L g9480 ( 
.A(n_8802),
.Y(n_9480)
);

INVx1_ASAP7_75t_L g9481 ( 
.A(n_8804),
.Y(n_9481)
);

AND2x2_ASAP7_75t_L g9482 ( 
.A(n_8891),
.B(n_5888),
.Y(n_9482)
);

INVx2_ASAP7_75t_L g9483 ( 
.A(n_8871),
.Y(n_9483)
);

NAND2xp5_ASAP7_75t_L g9484 ( 
.A(n_8679),
.B(n_5894),
.Y(n_9484)
);

BUFx4f_ASAP7_75t_L g9485 ( 
.A(n_9127),
.Y(n_9485)
);

NAND2xp5_ASAP7_75t_L g9486 ( 
.A(n_8655),
.B(n_5896),
.Y(n_9486)
);

AND2x6_ASAP7_75t_L g9487 ( 
.A(n_9119),
.B(n_5612),
.Y(n_9487)
);

BUFx2_ASAP7_75t_L g9488 ( 
.A(n_8895),
.Y(n_9488)
);

AND2x2_ASAP7_75t_L g9489 ( 
.A(n_9140),
.B(n_5897),
.Y(n_9489)
);

BUFx6f_ASAP7_75t_L g9490 ( 
.A(n_8980),
.Y(n_9490)
);

INVx1_ASAP7_75t_L g9491 ( 
.A(n_8807),
.Y(n_9491)
);

NOR2xp33_ASAP7_75t_L g9492 ( 
.A(n_9003),
.B(n_5898),
.Y(n_9492)
);

CKINVDCx6p67_ASAP7_75t_R g9493 ( 
.A(n_9099),
.Y(n_9493)
);

INVx1_ASAP7_75t_L g9494 ( 
.A(n_8810),
.Y(n_9494)
);

BUFx3_ASAP7_75t_L g9495 ( 
.A(n_8660),
.Y(n_9495)
);

INVx1_ASAP7_75t_L g9496 ( 
.A(n_8812),
.Y(n_9496)
);

INVx2_ASAP7_75t_L g9497 ( 
.A(n_8877),
.Y(n_9497)
);

AO22x2_ASAP7_75t_L g9498 ( 
.A1(n_8711),
.A2(n_5632),
.B1(n_5634),
.B2(n_5623),
.Y(n_9498)
);

INVx1_ASAP7_75t_L g9499 ( 
.A(n_8816),
.Y(n_9499)
);

NAND2xp5_ASAP7_75t_SL g9500 ( 
.A(n_9149),
.B(n_5899),
.Y(n_9500)
);

INVx2_ASAP7_75t_L g9501 ( 
.A(n_8817),
.Y(n_9501)
);

INVx5_ASAP7_75t_L g9502 ( 
.A(n_9127),
.Y(n_9502)
);

OR2x2_ASAP7_75t_L g9503 ( 
.A(n_8643),
.B(n_5902),
.Y(n_9503)
);

OAI22xp5_ASAP7_75t_L g9504 ( 
.A1(n_9111),
.A2(n_5904),
.B1(n_5905),
.B2(n_5903),
.Y(n_9504)
);

INVx1_ASAP7_75t_L g9505 ( 
.A(n_8818),
.Y(n_9505)
);

AND2x2_ASAP7_75t_L g9506 ( 
.A(n_9139),
.B(n_5908),
.Y(n_9506)
);

OAI22xp5_ASAP7_75t_L g9507 ( 
.A1(n_8652),
.A2(n_5911),
.B1(n_5912),
.B2(n_5909),
.Y(n_9507)
);

CKINVDCx5p33_ASAP7_75t_R g9508 ( 
.A(n_8791),
.Y(n_9508)
);

HB1xp67_ASAP7_75t_L g9509 ( 
.A(n_8786),
.Y(n_9509)
);

INVx1_ASAP7_75t_L g9510 ( 
.A(n_8822),
.Y(n_9510)
);

BUFx6f_ASAP7_75t_L g9511 ( 
.A(n_8980),
.Y(n_9511)
);

OAI22xp33_ASAP7_75t_SL g9512 ( 
.A1(n_9071),
.A2(n_5917),
.B1(n_5918),
.B2(n_5914),
.Y(n_9512)
);

INVx2_ASAP7_75t_L g9513 ( 
.A(n_8823),
.Y(n_9513)
);

AND2x4_ASAP7_75t_L g9514 ( 
.A(n_8806),
.B(n_5636),
.Y(n_9514)
);

INVx2_ASAP7_75t_L g9515 ( 
.A(n_8824),
.Y(n_9515)
);

BUFx3_ASAP7_75t_L g9516 ( 
.A(n_8813),
.Y(n_9516)
);

BUFx3_ASAP7_75t_L g9517 ( 
.A(n_8851),
.Y(n_9517)
);

INVx1_ASAP7_75t_L g9518 ( 
.A(n_8829),
.Y(n_9518)
);

AOI22xp5_ASAP7_75t_L g9519 ( 
.A1(n_9087),
.A2(n_9112),
.B1(n_9123),
.B2(n_8905),
.Y(n_9519)
);

INVx2_ASAP7_75t_L g9520 ( 
.A(n_8831),
.Y(n_9520)
);

INVx1_ASAP7_75t_L g9521 ( 
.A(n_8836),
.Y(n_9521)
);

INVx1_ASAP7_75t_L g9522 ( 
.A(n_8839),
.Y(n_9522)
);

INVx1_ASAP7_75t_L g9523 ( 
.A(n_8841),
.Y(n_9523)
);

INVxp67_ASAP7_75t_SL g9524 ( 
.A(n_8832),
.Y(n_9524)
);

OAI22xp5_ASAP7_75t_L g9525 ( 
.A1(n_8986),
.A2(n_5921),
.B1(n_5923),
.B2(n_5920),
.Y(n_9525)
);

NOR2xp33_ASAP7_75t_L g9526 ( 
.A(n_9054),
.B(n_5924),
.Y(n_9526)
);

NOR2xp33_ASAP7_75t_L g9527 ( 
.A(n_9157),
.B(n_5927),
.Y(n_9527)
);

INVx4_ASAP7_75t_L g9528 ( 
.A(n_8987),
.Y(n_9528)
);

NAND2xp5_ASAP7_75t_L g9529 ( 
.A(n_8685),
.B(n_5940),
.Y(n_9529)
);

BUFx3_ASAP7_75t_L g9530 ( 
.A(n_8885),
.Y(n_9530)
);

AND2x2_ASAP7_75t_L g9531 ( 
.A(n_8718),
.B(n_5942),
.Y(n_9531)
);

BUFx3_ASAP7_75t_L g9532 ( 
.A(n_8894),
.Y(n_9532)
);

NAND2xp5_ASAP7_75t_L g9533 ( 
.A(n_9070),
.B(n_5945),
.Y(n_9533)
);

NOR2x1p5_ASAP7_75t_L g9534 ( 
.A(n_9172),
.B(n_5949),
.Y(n_9534)
);

INVx1_ASAP7_75t_L g9535 ( 
.A(n_8843),
.Y(n_9535)
);

INVx1_ASAP7_75t_L g9536 ( 
.A(n_8844),
.Y(n_9536)
);

AND2x4_ASAP7_75t_L g9537 ( 
.A(n_8902),
.B(n_5645),
.Y(n_9537)
);

NAND2xp5_ASAP7_75t_SL g9538 ( 
.A(n_9099),
.B(n_5952),
.Y(n_9538)
);

INVx1_ASAP7_75t_L g9539 ( 
.A(n_8846),
.Y(n_9539)
);

NAND2xp5_ASAP7_75t_SL g9540 ( 
.A(n_9151),
.B(n_5955),
.Y(n_9540)
);

NOR2xp33_ASAP7_75t_L g9541 ( 
.A(n_9165),
.B(n_5958),
.Y(n_9541)
);

CKINVDCx5p33_ASAP7_75t_R g9542 ( 
.A(n_9096),
.Y(n_9542)
);

AO22x2_ASAP7_75t_L g9543 ( 
.A1(n_9162),
.A2(n_5650),
.B1(n_5651),
.B2(n_5648),
.Y(n_9543)
);

INVx1_ASAP7_75t_L g9544 ( 
.A(n_8978),
.Y(n_9544)
);

NAND2xp5_ASAP7_75t_L g9545 ( 
.A(n_8712),
.B(n_5963),
.Y(n_9545)
);

INVx2_ASAP7_75t_L g9546 ( 
.A(n_8847),
.Y(n_9546)
);

INVx1_ASAP7_75t_L g9547 ( 
.A(n_8979),
.Y(n_9547)
);

INVx8_ASAP7_75t_L g9548 ( 
.A(n_8974),
.Y(n_9548)
);

NOR2xp33_ASAP7_75t_L g9549 ( 
.A(n_8639),
.B(n_5964),
.Y(n_9549)
);

AND2x4_ASAP7_75t_L g9550 ( 
.A(n_9079),
.B(n_5653),
.Y(n_9550)
);

INVx3_ASAP7_75t_L g9551 ( 
.A(n_8987),
.Y(n_9551)
);

XOR2xp5_ASAP7_75t_L g9552 ( 
.A(n_8701),
.B(n_4336),
.Y(n_9552)
);

INVx2_ASAP7_75t_L g9553 ( 
.A(n_8848),
.Y(n_9553)
);

NOR2xp33_ASAP7_75t_L g9554 ( 
.A(n_9073),
.B(n_5965),
.Y(n_9554)
);

INVx2_ASAP7_75t_SL g9555 ( 
.A(n_9005),
.Y(n_9555)
);

XOR2xp5_ASAP7_75t_L g9556 ( 
.A(n_8748),
.B(n_4337),
.Y(n_9556)
);

AND2x6_ASAP7_75t_L g9557 ( 
.A(n_9114),
.B(n_5662),
.Y(n_9557)
);

INVx1_ASAP7_75t_L g9558 ( 
.A(n_8998),
.Y(n_9558)
);

INVx1_ASAP7_75t_L g9559 ( 
.A(n_8882),
.Y(n_9559)
);

INVx1_ASAP7_75t_L g9560 ( 
.A(n_8886),
.Y(n_9560)
);

INVx2_ASAP7_75t_L g9561 ( 
.A(n_8850),
.Y(n_9561)
);

INVx1_ASAP7_75t_L g9562 ( 
.A(n_8857),
.Y(n_9562)
);

NAND2xp5_ASAP7_75t_L g9563 ( 
.A(n_8634),
.B(n_5968),
.Y(n_9563)
);

INVx1_ASAP7_75t_L g9564 ( 
.A(n_8860),
.Y(n_9564)
);

BUFx10_ASAP7_75t_L g9565 ( 
.A(n_9104),
.Y(n_9565)
);

INVx2_ASAP7_75t_L g9566 ( 
.A(n_8864),
.Y(n_9566)
);

OR2x2_ASAP7_75t_L g9567 ( 
.A(n_8740),
.B(n_5969),
.Y(n_9567)
);

BUFx3_ASAP7_75t_L g9568 ( 
.A(n_9023),
.Y(n_9568)
);

INVx1_ASAP7_75t_L g9569 ( 
.A(n_8876),
.Y(n_9569)
);

AND2x6_ASAP7_75t_L g9570 ( 
.A(n_9117),
.B(n_5664),
.Y(n_9570)
);

BUFx3_ASAP7_75t_L g9571 ( 
.A(n_9023),
.Y(n_9571)
);

OR2x6_ASAP7_75t_L g9572 ( 
.A(n_8974),
.B(n_5667),
.Y(n_9572)
);

BUFx3_ASAP7_75t_L g9573 ( 
.A(n_9052),
.Y(n_9573)
);

INVx3_ASAP7_75t_L g9574 ( 
.A(n_9052),
.Y(n_9574)
);

BUFx6f_ASAP7_75t_L g9575 ( 
.A(n_8916),
.Y(n_9575)
);

BUFx3_ASAP7_75t_L g9576 ( 
.A(n_8955),
.Y(n_9576)
);

AOI22xp5_ASAP7_75t_L g9577 ( 
.A1(n_8855),
.A2(n_9122),
.B1(n_9066),
.B2(n_9135),
.Y(n_9577)
);

INVx3_ASAP7_75t_L g9578 ( 
.A(n_8966),
.Y(n_9578)
);

NAND2xp5_ASAP7_75t_L g9579 ( 
.A(n_8927),
.B(n_5970),
.Y(n_9579)
);

BUFx4f_ASAP7_75t_L g9580 ( 
.A(n_9150),
.Y(n_9580)
);

CKINVDCx8_ASAP7_75t_R g9581 ( 
.A(n_9145),
.Y(n_9581)
);

BUFx8_ASAP7_75t_SL g9582 ( 
.A(n_9166),
.Y(n_9582)
);

INVx4_ASAP7_75t_L g9583 ( 
.A(n_8981),
.Y(n_9583)
);

INVx2_ASAP7_75t_L g9584 ( 
.A(n_8889),
.Y(n_9584)
);

BUFx2_ASAP7_75t_L g9585 ( 
.A(n_8726),
.Y(n_9585)
);

BUFx3_ASAP7_75t_L g9586 ( 
.A(n_8977),
.Y(n_9586)
);

AND2x4_ASAP7_75t_L g9587 ( 
.A(n_9039),
.B(n_5671),
.Y(n_9587)
);

INVxp67_ASAP7_75t_SL g9588 ( 
.A(n_8835),
.Y(n_9588)
);

INVx3_ASAP7_75t_L g9589 ( 
.A(n_8976),
.Y(n_9589)
);

AND2x6_ASAP7_75t_L g9590 ( 
.A(n_9152),
.B(n_8990),
.Y(n_9590)
);

AND2x2_ASAP7_75t_L g9591 ( 
.A(n_9040),
.B(n_5971),
.Y(n_9591)
);

INVx1_ASAP7_75t_L g9592 ( 
.A(n_9036),
.Y(n_9592)
);

INVx2_ASAP7_75t_L g9593 ( 
.A(n_8892),
.Y(n_9593)
);

INVx2_ASAP7_75t_L g9594 ( 
.A(n_8896),
.Y(n_9594)
);

NAND2xp5_ASAP7_75t_SL g9595 ( 
.A(n_8788),
.B(n_5980),
.Y(n_9595)
);

INVx1_ASAP7_75t_L g9596 ( 
.A(n_9045),
.Y(n_9596)
);

BUFx6f_ASAP7_75t_L g9597 ( 
.A(n_9101),
.Y(n_9597)
);

OAI22xp5_ASAP7_75t_L g9598 ( 
.A1(n_9131),
.A2(n_5983),
.B1(n_5987),
.B2(n_5981),
.Y(n_9598)
);

INVx4_ASAP7_75t_L g9599 ( 
.A(n_8981),
.Y(n_9599)
);

OR2x2_ASAP7_75t_L g9600 ( 
.A(n_8988),
.B(n_5989),
.Y(n_9600)
);

INVx4_ASAP7_75t_L g9601 ( 
.A(n_8982),
.Y(n_9601)
);

INVx4_ASAP7_75t_L g9602 ( 
.A(n_8989),
.Y(n_9602)
);

AND2x4_ASAP7_75t_L g9603 ( 
.A(n_9046),
.B(n_5685),
.Y(n_9603)
);

INVx1_ASAP7_75t_L g9604 ( 
.A(n_8897),
.Y(n_9604)
);

BUFx4f_ASAP7_75t_L g9605 ( 
.A(n_9167),
.Y(n_9605)
);

AND2x2_ASAP7_75t_L g9606 ( 
.A(n_9041),
.B(n_5990),
.Y(n_9606)
);

INVx1_ASAP7_75t_SL g9607 ( 
.A(n_8819),
.Y(n_9607)
);

NOR2xp33_ASAP7_75t_L g9608 ( 
.A(n_8761),
.B(n_5991),
.Y(n_9608)
);

AND2x2_ASAP7_75t_L g9609 ( 
.A(n_8918),
.B(n_5992),
.Y(n_9609)
);

AO21x2_ASAP7_75t_L g9610 ( 
.A1(n_8653),
.A2(n_5697),
.B(n_5691),
.Y(n_9610)
);

INVx1_ASAP7_75t_L g9611 ( 
.A(n_8900),
.Y(n_9611)
);

INVx2_ASAP7_75t_L g9612 ( 
.A(n_8903),
.Y(n_9612)
);

INVx1_ASAP7_75t_SL g9613 ( 
.A(n_8837),
.Y(n_9613)
);

AND2x4_ASAP7_75t_L g9614 ( 
.A(n_8991),
.B(n_5703),
.Y(n_9614)
);

NOR2xp33_ASAP7_75t_SL g9615 ( 
.A(n_9173),
.B(n_5994),
.Y(n_9615)
);

INVx1_ASAP7_75t_L g9616 ( 
.A(n_8904),
.Y(n_9616)
);

OR2x6_ASAP7_75t_L g9617 ( 
.A(n_8910),
.B(n_5716),
.Y(n_9617)
);

AND2x4_ASAP7_75t_L g9618 ( 
.A(n_8992),
.B(n_5720),
.Y(n_9618)
);

INVx2_ASAP7_75t_L g9619 ( 
.A(n_8909),
.Y(n_9619)
);

BUFx3_ASAP7_75t_L g9620 ( 
.A(n_9037),
.Y(n_9620)
);

BUFx3_ASAP7_75t_L g9621 ( 
.A(n_9044),
.Y(n_9621)
);

INVx1_ASAP7_75t_L g9622 ( 
.A(n_8915),
.Y(n_9622)
);

AND2x6_ASAP7_75t_L g9623 ( 
.A(n_8999),
.B(n_5722),
.Y(n_9623)
);

NAND2xp5_ASAP7_75t_SL g9624 ( 
.A(n_9051),
.B(n_5996),
.Y(n_9624)
);

INVx2_ASAP7_75t_L g9625 ( 
.A(n_8919),
.Y(n_9625)
);

INVx1_ASAP7_75t_L g9626 ( 
.A(n_8920),
.Y(n_9626)
);

INVx2_ASAP7_75t_SL g9627 ( 
.A(n_8827),
.Y(n_9627)
);

NOR2xp33_ASAP7_75t_L g9628 ( 
.A(n_8778),
.B(n_6003),
.Y(n_9628)
);

CKINVDCx5p33_ASAP7_75t_R g9629 ( 
.A(n_8766),
.Y(n_9629)
);

AND2x4_ASAP7_75t_L g9630 ( 
.A(n_8914),
.B(n_5749),
.Y(n_9630)
);

BUFx2_ASAP7_75t_L g9631 ( 
.A(n_8925),
.Y(n_9631)
);

BUFx2_ASAP7_75t_L g9632 ( 
.A(n_8997),
.Y(n_9632)
);

INVxp67_ASAP7_75t_SL g9633 ( 
.A(n_9015),
.Y(n_9633)
);

BUFx3_ASAP7_75t_L g9634 ( 
.A(n_9018),
.Y(n_9634)
);

NOR2xp33_ASAP7_75t_L g9635 ( 
.A(n_8794),
.B(n_6010),
.Y(n_9635)
);

AND2x4_ASAP7_75t_L g9636 ( 
.A(n_9022),
.B(n_5751),
.Y(n_9636)
);

INVx1_ASAP7_75t_L g9637 ( 
.A(n_8922),
.Y(n_9637)
);

INVx2_ASAP7_75t_L g9638 ( 
.A(n_8901),
.Y(n_9638)
);

INVx1_ASAP7_75t_L g9639 ( 
.A(n_9095),
.Y(n_9639)
);

AND3x2_ASAP7_75t_L g9640 ( 
.A(n_9164),
.B(n_5756),
.C(n_5755),
.Y(n_9640)
);

INVx5_ASAP7_75t_L g9641 ( 
.A(n_9030),
.Y(n_9641)
);

INVx1_ASAP7_75t_L g9642 ( 
.A(n_8929),
.Y(n_9642)
);

BUFx10_ASAP7_75t_L g9643 ( 
.A(n_9170),
.Y(n_9643)
);

NAND2xp5_ASAP7_75t_L g9644 ( 
.A(n_8932),
.B(n_6012),
.Y(n_9644)
);

AND2x6_ASAP7_75t_L g9645 ( 
.A(n_9126),
.B(n_5770),
.Y(n_9645)
);

OR2x6_ASAP7_75t_L g9646 ( 
.A(n_9009),
.B(n_5775),
.Y(n_9646)
);

BUFx4f_ASAP7_75t_L g9647 ( 
.A(n_9030),
.Y(n_9647)
);

INVx1_ASAP7_75t_L g9648 ( 
.A(n_8933),
.Y(n_9648)
);

INVx1_ASAP7_75t_L g9649 ( 
.A(n_8937),
.Y(n_9649)
);

NAND2xp5_ASAP7_75t_SL g9650 ( 
.A(n_9121),
.B(n_6017),
.Y(n_9650)
);

INVx4_ASAP7_75t_L g9651 ( 
.A(n_9025),
.Y(n_9651)
);

INVx1_ASAP7_75t_L g9652 ( 
.A(n_8938),
.Y(n_9652)
);

INVx3_ASAP7_75t_L g9653 ( 
.A(n_9078),
.Y(n_9653)
);

NOR2x1p5_ASAP7_75t_L g9654 ( 
.A(n_9169),
.B(n_9174),
.Y(n_9654)
);

INVx2_ASAP7_75t_L g9655 ( 
.A(n_8907),
.Y(n_9655)
);

INVx2_ASAP7_75t_L g9656 ( 
.A(n_8908),
.Y(n_9656)
);

INVx1_ASAP7_75t_L g9657 ( 
.A(n_8939),
.Y(n_9657)
);

INVx2_ASAP7_75t_SL g9658 ( 
.A(n_9072),
.Y(n_9658)
);

NAND3x1_ASAP7_75t_L g9659 ( 
.A(n_8996),
.B(n_5779),
.C(n_5777),
.Y(n_9659)
);

INVx3_ASAP7_75t_L g9660 ( 
.A(n_9085),
.Y(n_9660)
);

INVx1_ASAP7_75t_L g9661 ( 
.A(n_8946),
.Y(n_9661)
);

AND2x4_ASAP7_75t_L g9662 ( 
.A(n_9057),
.B(n_5780),
.Y(n_9662)
);

NAND2xp5_ASAP7_75t_L g9663 ( 
.A(n_8950),
.B(n_6018),
.Y(n_9663)
);

INVx1_ASAP7_75t_L g9664 ( 
.A(n_8958),
.Y(n_9664)
);

NAND2xp5_ASAP7_75t_SL g9665 ( 
.A(n_9133),
.B(n_6025),
.Y(n_9665)
);

BUFx6f_ASAP7_75t_L g9666 ( 
.A(n_9062),
.Y(n_9666)
);

BUFx10_ASAP7_75t_L g9667 ( 
.A(n_9080),
.Y(n_9667)
);

INVx2_ASAP7_75t_L g9668 ( 
.A(n_8921),
.Y(n_9668)
);

BUFx4_ASAP7_75t_L g9669 ( 
.A(n_9053),
.Y(n_9669)
);

AND2x4_ASAP7_75t_L g9670 ( 
.A(n_9063),
.B(n_9067),
.Y(n_9670)
);

AOI22xp5_ASAP7_75t_L g9671 ( 
.A1(n_9030),
.A2(n_9129),
.B1(n_9128),
.B2(n_8751),
.Y(n_9671)
);

OR2x6_ASAP7_75t_L g9672 ( 
.A(n_9029),
.B(n_5781),
.Y(n_9672)
);

INVxp33_ASAP7_75t_SL g9673 ( 
.A(n_9068),
.Y(n_9673)
);

NAND2xp5_ASAP7_75t_SL g9674 ( 
.A(n_8890),
.B(n_8944),
.Y(n_9674)
);

NOR2xp33_ASAP7_75t_L g9675 ( 
.A(n_8859),
.B(n_6026),
.Y(n_9675)
);

INVx1_ASAP7_75t_L g9676 ( 
.A(n_8965),
.Y(n_9676)
);

BUFx3_ASAP7_75t_L g9677 ( 
.A(n_9076),
.Y(n_9677)
);

INVx1_ASAP7_75t_L g9678 ( 
.A(n_8969),
.Y(n_9678)
);

INVx2_ASAP7_75t_SL g9679 ( 
.A(n_9069),
.Y(n_9679)
);

INVx1_ASAP7_75t_L g9680 ( 
.A(n_8973),
.Y(n_9680)
);

INVx2_ASAP7_75t_L g9681 ( 
.A(n_8928),
.Y(n_9681)
);

INVx1_ASAP7_75t_SL g9682 ( 
.A(n_9143),
.Y(n_9682)
);

INVx1_ASAP7_75t_L g9683 ( 
.A(n_8930),
.Y(n_9683)
);

BUFx10_ASAP7_75t_L g9684 ( 
.A(n_9058),
.Y(n_9684)
);

OR2x6_ASAP7_75t_L g9685 ( 
.A(n_9086),
.B(n_5783),
.Y(n_9685)
);

NOR2xp33_ASAP7_75t_L g9686 ( 
.A(n_8934),
.B(n_6028),
.Y(n_9686)
);

NOR2xp33_ASAP7_75t_L g9687 ( 
.A(n_9272),
.B(n_8636),
.Y(n_9687)
);

INVx1_ASAP7_75t_L g9688 ( 
.A(n_9185),
.Y(n_9688)
);

INVxp67_ASAP7_75t_SL g9689 ( 
.A(n_9509),
.Y(n_9689)
);

NAND2xp5_ASAP7_75t_L g9690 ( 
.A(n_9264),
.B(n_8931),
.Y(n_9690)
);

NOR2xp33_ASAP7_75t_L g9691 ( 
.A(n_9219),
.B(n_8647),
.Y(n_9691)
);

INVx1_ASAP7_75t_L g9692 ( 
.A(n_9188),
.Y(n_9692)
);

NOR2xp33_ASAP7_75t_L g9693 ( 
.A(n_9182),
.B(n_8672),
.Y(n_9693)
);

HB1xp67_ASAP7_75t_L g9694 ( 
.A(n_9233),
.Y(n_9694)
);

NAND2xp5_ASAP7_75t_L g9695 ( 
.A(n_9196),
.B(n_8967),
.Y(n_9695)
);

NAND2xp5_ASAP7_75t_L g9696 ( 
.A(n_9309),
.B(n_9163),
.Y(n_9696)
);

NOR2xp67_ASAP7_75t_SL g9697 ( 
.A(n_9189),
.B(n_9130),
.Y(n_9697)
);

NAND2xp5_ASAP7_75t_L g9698 ( 
.A(n_9290),
.B(n_8830),
.Y(n_9698)
);

INVx2_ASAP7_75t_SL g9699 ( 
.A(n_9406),
.Y(n_9699)
);

INVx1_ASAP7_75t_L g9700 ( 
.A(n_9191),
.Y(n_9700)
);

OAI22xp5_ASAP7_75t_L g9701 ( 
.A1(n_9367),
.A2(n_9674),
.B1(n_9577),
.B2(n_9519),
.Y(n_9701)
);

AND2x6_ASAP7_75t_SL g9702 ( 
.A(n_9193),
.B(n_9175),
.Y(n_9702)
);

AOI22xp5_ASAP7_75t_L g9703 ( 
.A1(n_9209),
.A2(n_9212),
.B1(n_9210),
.B2(n_9361),
.Y(n_9703)
);

INVx1_ASAP7_75t_L g9704 ( 
.A(n_9192),
.Y(n_9704)
);

INVx1_ASAP7_75t_L g9705 ( 
.A(n_9199),
.Y(n_9705)
);

NAND2xp5_ASAP7_75t_L g9706 ( 
.A(n_9277),
.B(n_9105),
.Y(n_9706)
);

NAND2x1p5_ASAP7_75t_L g9707 ( 
.A(n_9189),
.B(n_9065),
.Y(n_9707)
);

INVx1_ASAP7_75t_L g9708 ( 
.A(n_9201),
.Y(n_9708)
);

BUFx8_ASAP7_75t_L g9709 ( 
.A(n_9495),
.Y(n_9709)
);

NOR2xp33_ASAP7_75t_L g9710 ( 
.A(n_9228),
.B(n_8945),
.Y(n_9710)
);

NOR3xp33_ASAP7_75t_L g9711 ( 
.A(n_9273),
.B(n_8947),
.C(n_8873),
.Y(n_9711)
);

NOR2xp33_ASAP7_75t_SL g9712 ( 
.A(n_9204),
.B(n_8767),
.Y(n_9712)
);

NAND2xp5_ASAP7_75t_SL g9713 ( 
.A(n_9402),
.B(n_9090),
.Y(n_9713)
);

INVx2_ASAP7_75t_L g9714 ( 
.A(n_9501),
.Y(n_9714)
);

AND2x2_ASAP7_75t_L g9715 ( 
.A(n_9237),
.B(n_9083),
.Y(n_9715)
);

A2O1A1Ixp33_ASAP7_75t_L g9716 ( 
.A1(n_9468),
.A2(n_8954),
.B(n_8926),
.C(n_8803),
.Y(n_9716)
);

OAI22xp5_ASAP7_75t_L g9717 ( 
.A1(n_9202),
.A2(n_9019),
.B1(n_9077),
.B2(n_9074),
.Y(n_9717)
);

NAND2xp5_ASAP7_75t_L g9718 ( 
.A(n_9400),
.B(n_8694),
.Y(n_9718)
);

NAND2xp5_ASAP7_75t_L g9719 ( 
.A(n_9276),
.B(n_9545),
.Y(n_9719)
);

NAND2xp5_ASAP7_75t_SL g9720 ( 
.A(n_9275),
.B(n_8790),
.Y(n_9720)
);

BUFx6f_ASAP7_75t_SL g9721 ( 
.A(n_9306),
.Y(n_9721)
);

AND2x4_ASAP7_75t_L g9722 ( 
.A(n_9180),
.B(n_9043),
.Y(n_9722)
);

NOR2x1p5_ASAP7_75t_L g9723 ( 
.A(n_9493),
.B(n_9048),
.Y(n_9723)
);

O2A1O1Ixp33_ASAP7_75t_L g9724 ( 
.A1(n_9512),
.A2(n_8739),
.B(n_8745),
.C(n_8707),
.Y(n_9724)
);

NAND2xp5_ASAP7_75t_SL g9725 ( 
.A(n_9433),
.B(n_8809),
.Y(n_9725)
);

INVx1_ASAP7_75t_L g9726 ( 
.A(n_9213),
.Y(n_9726)
);

NAND2xp5_ASAP7_75t_L g9727 ( 
.A(n_9531),
.B(n_9049),
.Y(n_9727)
);

NAND2xp5_ASAP7_75t_L g9728 ( 
.A(n_9304),
.B(n_8856),
.Y(n_9728)
);

OR2x6_ASAP7_75t_L g9729 ( 
.A(n_9412),
.B(n_9081),
.Y(n_9729)
);

INVx8_ASAP7_75t_L g9730 ( 
.A(n_9406),
.Y(n_9730)
);

BUFx5_ASAP7_75t_L g9731 ( 
.A(n_9215),
.Y(n_9731)
);

INVx1_ASAP7_75t_L g9732 ( 
.A(n_9216),
.Y(n_9732)
);

INVx2_ASAP7_75t_SL g9733 ( 
.A(n_9176),
.Y(n_9733)
);

AOI22x1_ASAP7_75t_L g9734 ( 
.A1(n_9350),
.A2(n_8993),
.B1(n_9093),
.B2(n_9034),
.Y(n_9734)
);

NAND2xp5_ASAP7_75t_SL g9735 ( 
.A(n_9374),
.B(n_8952),
.Y(n_9735)
);

INVx2_ASAP7_75t_L g9736 ( 
.A(n_9513),
.Y(n_9736)
);

AND2x2_ASAP7_75t_L g9737 ( 
.A(n_9437),
.B(n_9020),
.Y(n_9737)
);

AOI22xp33_ASAP7_75t_L g9738 ( 
.A1(n_9591),
.A2(n_8971),
.B1(n_8913),
.B2(n_8868),
.Y(n_9738)
);

INVx2_ASAP7_75t_L g9739 ( 
.A(n_9515),
.Y(n_9739)
);

INVx1_ASAP7_75t_SL g9740 ( 
.A(n_9303),
.Y(n_9740)
);

NAND2xp5_ASAP7_75t_L g9741 ( 
.A(n_9308),
.B(n_9075),
.Y(n_9741)
);

NAND2x1_ASAP7_75t_L g9742 ( 
.A(n_9183),
.B(n_9004),
.Y(n_9742)
);

NAND2x1p5_ASAP7_75t_L g9743 ( 
.A(n_9301),
.B(n_9082),
.Y(n_9743)
);

NAND2xp5_ASAP7_75t_SL g9744 ( 
.A(n_9282),
.B(n_9084),
.Y(n_9744)
);

INVx1_ASAP7_75t_L g9745 ( 
.A(n_9217),
.Y(n_9745)
);

CKINVDCx5p33_ASAP7_75t_R g9746 ( 
.A(n_9249),
.Y(n_9746)
);

INVx8_ASAP7_75t_L g9747 ( 
.A(n_9301),
.Y(n_9747)
);

NAND2xp5_ASAP7_75t_SL g9748 ( 
.A(n_9310),
.B(n_9091),
.Y(n_9748)
);

NAND2xp5_ASAP7_75t_L g9749 ( 
.A(n_9314),
.B(n_9322),
.Y(n_9749)
);

INVxp67_ASAP7_75t_L g9750 ( 
.A(n_9585),
.Y(n_9750)
);

NAND2xp5_ASAP7_75t_SL g9751 ( 
.A(n_9184),
.B(n_9092),
.Y(n_9751)
);

NAND2xp5_ASAP7_75t_L g9752 ( 
.A(n_9326),
.B(n_9097),
.Y(n_9752)
);

NAND2xp5_ASAP7_75t_L g9753 ( 
.A(n_9337),
.B(n_9144),
.Y(n_9753)
);

NAND2xp5_ASAP7_75t_SL g9754 ( 
.A(n_9455),
.B(n_8838),
.Y(n_9754)
);

NOR2xp67_ASAP7_75t_L g9755 ( 
.A(n_9542),
.B(n_9061),
.Y(n_9755)
);

AND2x6_ASAP7_75t_SL g9756 ( 
.A(n_9221),
.B(n_5786),
.Y(n_9756)
);

AND2x2_ASAP7_75t_L g9757 ( 
.A(n_9246),
.B(n_9124),
.Y(n_9757)
);

NAND2xp5_ASAP7_75t_L g9758 ( 
.A(n_9345),
.B(n_9474),
.Y(n_9758)
);

INVx2_ASAP7_75t_L g9759 ( 
.A(n_9520),
.Y(n_9759)
);

AOI21xp5_ASAP7_75t_L g9760 ( 
.A1(n_9297),
.A2(n_8924),
.B(n_9094),
.Y(n_9760)
);

INVx1_ASAP7_75t_L g9761 ( 
.A(n_9225),
.Y(n_9761)
);

INVx2_ASAP7_75t_L g9762 ( 
.A(n_9234),
.Y(n_9762)
);

INVx1_ASAP7_75t_L g9763 ( 
.A(n_9239),
.Y(n_9763)
);

INVx1_ASAP7_75t_L g9764 ( 
.A(n_9243),
.Y(n_9764)
);

OAI221xp5_ASAP7_75t_L g9765 ( 
.A1(n_9686),
.A2(n_8692),
.B1(n_9120),
.B2(n_9158),
.C(n_8957),
.Y(n_9765)
);

INVx2_ASAP7_75t_L g9766 ( 
.A(n_9244),
.Y(n_9766)
);

INVx1_ASAP7_75t_L g9767 ( 
.A(n_9252),
.Y(n_9767)
);

NAND2xp33_ASAP7_75t_L g9768 ( 
.A(n_9629),
.B(n_8686),
.Y(n_9768)
);

INVx2_ASAP7_75t_L g9769 ( 
.A(n_9270),
.Y(n_9769)
);

NOR2xp33_ASAP7_75t_L g9770 ( 
.A(n_9473),
.B(n_9141),
.Y(n_9770)
);

INVx1_ASAP7_75t_L g9771 ( 
.A(n_9285),
.Y(n_9771)
);

INVx1_ASAP7_75t_L g9772 ( 
.A(n_9293),
.Y(n_9772)
);

NAND2xp5_ASAP7_75t_SL g9773 ( 
.A(n_9613),
.B(n_9042),
.Y(n_9773)
);

OR2x6_ASAP7_75t_L g9774 ( 
.A(n_9548),
.B(n_8763),
.Y(n_9774)
);

INVxp67_ASAP7_75t_L g9775 ( 
.A(n_9214),
.Y(n_9775)
);

NAND2xp5_ASAP7_75t_SL g9776 ( 
.A(n_9186),
.B(n_6031),
.Y(n_9776)
);

AOI22xp33_ASAP7_75t_L g9777 ( 
.A1(n_9606),
.A2(n_9161),
.B1(n_5793),
.B2(n_5802),
.Y(n_9777)
);

NAND2xp5_ASAP7_75t_L g9778 ( 
.A(n_9484),
.B(n_5791),
.Y(n_9778)
);

NAND2xp5_ASAP7_75t_L g9779 ( 
.A(n_9486),
.B(n_5805),
.Y(n_9779)
);

INVx1_ASAP7_75t_L g9780 ( 
.A(n_9298),
.Y(n_9780)
);

BUFx6f_ASAP7_75t_SL g9781 ( 
.A(n_9335),
.Y(n_9781)
);

AOI22xp5_ASAP7_75t_L g9782 ( 
.A1(n_9320),
.A2(n_9527),
.B1(n_9554),
.B2(n_9526),
.Y(n_9782)
);

OAI22xp5_ASAP7_75t_L g9783 ( 
.A1(n_9300),
.A2(n_6038),
.B1(n_6040),
.B2(n_6034),
.Y(n_9783)
);

INVx4_ASAP7_75t_L g9784 ( 
.A(n_9206),
.Y(n_9784)
);

INVx2_ASAP7_75t_L g9785 ( 
.A(n_9316),
.Y(n_9785)
);

NAND2xp33_ASAP7_75t_L g9786 ( 
.A(n_9211),
.B(n_6041),
.Y(n_9786)
);

NOR2xp33_ASAP7_75t_SL g9787 ( 
.A(n_9266),
.B(n_6044),
.Y(n_9787)
);

INVxp67_ASAP7_75t_L g9788 ( 
.A(n_9232),
.Y(n_9788)
);

NAND3xp33_ASAP7_75t_SL g9789 ( 
.A(n_9671),
.B(n_6048),
.C(n_6046),
.Y(n_9789)
);

NAND2xp33_ASAP7_75t_L g9790 ( 
.A(n_9590),
.B(n_6049),
.Y(n_9790)
);

AND2x2_ASAP7_75t_L g9791 ( 
.A(n_9257),
.B(n_6052),
.Y(n_9791)
);

INVx2_ASAP7_75t_L g9792 ( 
.A(n_9321),
.Y(n_9792)
);

NAND2xp5_ASAP7_75t_L g9793 ( 
.A(n_9529),
.B(n_9223),
.Y(n_9793)
);

NAND2xp5_ASAP7_75t_SL g9794 ( 
.A(n_9456),
.B(n_6058),
.Y(n_9794)
);

INVx1_ASAP7_75t_L g9795 ( 
.A(n_9323),
.Y(n_9795)
);

INVx1_ASAP7_75t_L g9796 ( 
.A(n_9331),
.Y(n_9796)
);

NAND2xp5_ASAP7_75t_L g9797 ( 
.A(n_9235),
.B(n_5806),
.Y(n_9797)
);

OAI22xp5_ASAP7_75t_L g9798 ( 
.A1(n_9338),
.A2(n_6061),
.B1(n_6062),
.B2(n_6060),
.Y(n_9798)
);

AND2x6_ASAP7_75t_L g9799 ( 
.A(n_9682),
.B(n_5807),
.Y(n_9799)
);

NAND2xp5_ASAP7_75t_L g9800 ( 
.A(n_9236),
.B(n_5813),
.Y(n_9800)
);

NAND2xp5_ASAP7_75t_L g9801 ( 
.A(n_9250),
.B(n_5822),
.Y(n_9801)
);

INVx2_ASAP7_75t_L g9802 ( 
.A(n_9343),
.Y(n_9802)
);

NAND2xp5_ASAP7_75t_SL g9803 ( 
.A(n_9476),
.B(n_6063),
.Y(n_9803)
);

NAND2xp5_ASAP7_75t_L g9804 ( 
.A(n_9259),
.B(n_5823),
.Y(n_9804)
);

NAND2xp5_ASAP7_75t_L g9805 ( 
.A(n_9533),
.B(n_5824),
.Y(n_9805)
);

INVx2_ASAP7_75t_L g9806 ( 
.A(n_9348),
.Y(n_9806)
);

INVx3_ASAP7_75t_L g9807 ( 
.A(n_9224),
.Y(n_9807)
);

NAND2xp5_ASAP7_75t_L g9808 ( 
.A(n_9359),
.B(n_5825),
.Y(n_9808)
);

AOI22xp33_ASAP7_75t_L g9809 ( 
.A1(n_9242),
.A2(n_5832),
.B1(n_5835),
.B2(n_5831),
.Y(n_9809)
);

BUFx2_ASAP7_75t_L g9810 ( 
.A(n_9586),
.Y(n_9810)
);

AND2x6_ASAP7_75t_L g9811 ( 
.A(n_9360),
.B(n_5862),
.Y(n_9811)
);

NOR2xp33_ASAP7_75t_SL g9812 ( 
.A(n_9327),
.B(n_6064),
.Y(n_9812)
);

INVx2_ASAP7_75t_L g9813 ( 
.A(n_9362),
.Y(n_9813)
);

NOR2xp33_ASAP7_75t_L g9814 ( 
.A(n_9312),
.B(n_6073),
.Y(n_9814)
);

INVx1_ASAP7_75t_L g9815 ( 
.A(n_9363),
.Y(n_9815)
);

INVx1_ASAP7_75t_L g9816 ( 
.A(n_9377),
.Y(n_9816)
);

INVx2_ASAP7_75t_L g9817 ( 
.A(n_9380),
.Y(n_9817)
);

NAND2xp5_ASAP7_75t_L g9818 ( 
.A(n_9395),
.B(n_5866),
.Y(n_9818)
);

INVx2_ASAP7_75t_L g9819 ( 
.A(n_9397),
.Y(n_9819)
);

NOR2xp33_ASAP7_75t_L g9820 ( 
.A(n_9274),
.B(n_6076),
.Y(n_9820)
);

INVx4_ASAP7_75t_L g9821 ( 
.A(n_9178),
.Y(n_9821)
);

INVx2_ASAP7_75t_SL g9822 ( 
.A(n_9502),
.Y(n_9822)
);

BUFx3_ASAP7_75t_L g9823 ( 
.A(n_9248),
.Y(n_9823)
);

AOI22xp5_ASAP7_75t_L g9824 ( 
.A1(n_9340),
.A2(n_6093),
.B1(n_6095),
.B2(n_6090),
.Y(n_9824)
);

AND2x2_ASAP7_75t_L g9825 ( 
.A(n_9262),
.B(n_6097),
.Y(n_9825)
);

AND2x2_ASAP7_75t_L g9826 ( 
.A(n_9305),
.B(n_6103),
.Y(n_9826)
);

INVxp67_ASAP7_75t_L g9827 ( 
.A(n_9631),
.Y(n_9827)
);

O2A1O1Ixp5_ASAP7_75t_L g9828 ( 
.A1(n_9650),
.A2(n_9665),
.B(n_9258),
.C(n_9218),
.Y(n_9828)
);

NAND2xp5_ASAP7_75t_L g9829 ( 
.A(n_9401),
.B(n_5868),
.Y(n_9829)
);

NAND2xp5_ASAP7_75t_L g9830 ( 
.A(n_9403),
.B(n_9407),
.Y(n_9830)
);

INVx2_ASAP7_75t_L g9831 ( 
.A(n_9413),
.Y(n_9831)
);

INVx2_ASAP7_75t_L g9832 ( 
.A(n_9419),
.Y(n_9832)
);

NAND2xp5_ASAP7_75t_SL g9833 ( 
.A(n_9488),
.B(n_6109),
.Y(n_9833)
);

NAND2xp5_ASAP7_75t_SL g9834 ( 
.A(n_9580),
.B(n_6112),
.Y(n_9834)
);

AOI22xp5_ASAP7_75t_L g9835 ( 
.A1(n_9177),
.A2(n_6122),
.B1(n_6123),
.B2(n_6118),
.Y(n_9835)
);

INVx2_ASAP7_75t_L g9836 ( 
.A(n_9424),
.Y(n_9836)
);

BUFx5_ASAP7_75t_L g9837 ( 
.A(n_9427),
.Y(n_9837)
);

NOR2xp33_ASAP7_75t_L g9838 ( 
.A(n_9460),
.B(n_6124),
.Y(n_9838)
);

INVx3_ASAP7_75t_L g9839 ( 
.A(n_9462),
.Y(n_9839)
);

INVx2_ASAP7_75t_L g9840 ( 
.A(n_9428),
.Y(n_9840)
);

NAND2xp5_ASAP7_75t_L g9841 ( 
.A(n_9429),
.B(n_5872),
.Y(n_9841)
);

CKINVDCx5p33_ASAP7_75t_R g9842 ( 
.A(n_9435),
.Y(n_9842)
);

INVx2_ASAP7_75t_L g9843 ( 
.A(n_9440),
.Y(n_9843)
);

AOI22xp5_ASAP7_75t_L g9844 ( 
.A1(n_9608),
.A2(n_6128),
.B1(n_6130),
.B2(n_6126),
.Y(n_9844)
);

INVx1_ASAP7_75t_L g9845 ( 
.A(n_9443),
.Y(n_9845)
);

INVxp67_ASAP7_75t_SL g9846 ( 
.A(n_9524),
.Y(n_9846)
);

NAND2xp33_ASAP7_75t_L g9847 ( 
.A(n_9590),
.B(n_6131),
.Y(n_9847)
);

NAND2xp5_ASAP7_75t_SL g9848 ( 
.A(n_9555),
.B(n_6136),
.Y(n_9848)
);

AOI22xp33_ASAP7_75t_L g9849 ( 
.A1(n_9628),
.A2(n_9635),
.B1(n_9675),
.B2(n_9459),
.Y(n_9849)
);

INVx2_ASAP7_75t_L g9850 ( 
.A(n_9453),
.Y(n_9850)
);

OAI22xp5_ASAP7_75t_L g9851 ( 
.A1(n_9454),
.A2(n_6139),
.B1(n_6140),
.B2(n_6138),
.Y(n_9851)
);

NAND2xp5_ASAP7_75t_L g9852 ( 
.A(n_9457),
.B(n_5873),
.Y(n_9852)
);

NOR2xp33_ASAP7_75t_L g9853 ( 
.A(n_9588),
.B(n_6143),
.Y(n_9853)
);

INVxp33_ASAP7_75t_L g9854 ( 
.A(n_9307),
.Y(n_9854)
);

OAI21xp5_ASAP7_75t_L g9855 ( 
.A1(n_9563),
.A2(n_5876),
.B(n_5874),
.Y(n_9855)
);

NAND2xp33_ASAP7_75t_L g9856 ( 
.A(n_9654),
.B(n_6145),
.Y(n_9856)
);

INVxp67_ASAP7_75t_L g9857 ( 
.A(n_9198),
.Y(n_9857)
);

AO221x1_ASAP7_75t_L g9858 ( 
.A1(n_9498),
.A2(n_5891),
.B1(n_5892),
.B2(n_5889),
.C(n_5881),
.Y(n_9858)
);

AND2x2_ASAP7_75t_L g9859 ( 
.A(n_9324),
.B(n_6148),
.Y(n_9859)
);

AOI22xp33_ASAP7_75t_L g9860 ( 
.A1(n_9609),
.A2(n_9624),
.B1(n_9507),
.B2(n_9241),
.Y(n_9860)
);

INVx1_ASAP7_75t_L g9861 ( 
.A(n_9458),
.Y(n_9861)
);

AND2x2_ASAP7_75t_L g9862 ( 
.A(n_9325),
.B(n_9351),
.Y(n_9862)
);

NAND2xp33_ASAP7_75t_L g9863 ( 
.A(n_9666),
.B(n_6149),
.Y(n_9863)
);

INVx2_ASAP7_75t_L g9864 ( 
.A(n_9642),
.Y(n_9864)
);

BUFx6f_ASAP7_75t_L g9865 ( 
.A(n_9178),
.Y(n_9865)
);

INVxp67_ASAP7_75t_L g9866 ( 
.A(n_9334),
.Y(n_9866)
);

AOI22xp33_ASAP7_75t_L g9867 ( 
.A1(n_9289),
.A2(n_5900),
.B1(n_5907),
.B2(n_5895),
.Y(n_9867)
);

NAND2xp5_ASAP7_75t_L g9868 ( 
.A(n_9544),
.B(n_5913),
.Y(n_9868)
);

NAND2xp5_ASAP7_75t_SL g9869 ( 
.A(n_9615),
.B(n_6150),
.Y(n_9869)
);

NAND3x1_ASAP7_75t_L g9870 ( 
.A(n_9179),
.B(n_5929),
.C(n_5916),
.Y(n_9870)
);

NAND2xp5_ASAP7_75t_L g9871 ( 
.A(n_9547),
.B(n_5933),
.Y(n_9871)
);

INVx1_ASAP7_75t_L g9872 ( 
.A(n_9463),
.Y(n_9872)
);

NAND2xp5_ASAP7_75t_L g9873 ( 
.A(n_9558),
.B(n_9592),
.Y(n_9873)
);

OAI22xp33_ASAP7_75t_L g9874 ( 
.A1(n_9347),
.A2(n_6157),
.B1(n_6158),
.B2(n_6152),
.Y(n_9874)
);

AOI22xp5_ASAP7_75t_L g9875 ( 
.A1(n_9541),
.A2(n_6166),
.B1(n_6167),
.B2(n_6165),
.Y(n_9875)
);

INVx2_ASAP7_75t_L g9876 ( 
.A(n_9648),
.Y(n_9876)
);

INVx2_ASAP7_75t_SL g9877 ( 
.A(n_9502),
.Y(n_9877)
);

NAND2xp5_ASAP7_75t_L g9878 ( 
.A(n_9596),
.B(n_5935),
.Y(n_9878)
);

AND2x2_ASAP7_75t_L g9879 ( 
.A(n_9471),
.B(n_6168),
.Y(n_9879)
);

NAND2xp5_ASAP7_75t_SL g9880 ( 
.A(n_9605),
.B(n_6170),
.Y(n_9880)
);

AOI22xp33_ASAP7_75t_L g9881 ( 
.A1(n_9595),
.A2(n_5938),
.B1(n_5941),
.B2(n_5936),
.Y(n_9881)
);

AND2x2_ASAP7_75t_L g9882 ( 
.A(n_9405),
.B(n_6173),
.Y(n_9882)
);

NAND2xp5_ASAP7_75t_L g9883 ( 
.A(n_9639),
.B(n_5946),
.Y(n_9883)
);

NAND2xp5_ASAP7_75t_SL g9884 ( 
.A(n_9666),
.B(n_9670),
.Y(n_9884)
);

OR2x2_ASAP7_75t_L g9885 ( 
.A(n_9423),
.B(n_6174),
.Y(n_9885)
);

NAND2xp5_ASAP7_75t_L g9886 ( 
.A(n_9477),
.B(n_5947),
.Y(n_9886)
);

INVx1_ASAP7_75t_L g9887 ( 
.A(n_9480),
.Y(n_9887)
);

NOR2xp33_ASAP7_75t_SL g9888 ( 
.A(n_9263),
.B(n_6175),
.Y(n_9888)
);

NAND2xp5_ASAP7_75t_L g9889 ( 
.A(n_9481),
.B(n_5948),
.Y(n_9889)
);

OR2x6_ASAP7_75t_L g9890 ( 
.A(n_9269),
.B(n_9181),
.Y(n_9890)
);

NAND2xp5_ASAP7_75t_L g9891 ( 
.A(n_9491),
.B(n_5959),
.Y(n_9891)
);

NAND2xp5_ASAP7_75t_SL g9892 ( 
.A(n_9339),
.B(n_9597),
.Y(n_9892)
);

INVx1_ASAP7_75t_L g9893 ( 
.A(n_9494),
.Y(n_9893)
);

NAND2xp5_ASAP7_75t_L g9894 ( 
.A(n_9496),
.B(n_5962),
.Y(n_9894)
);

NAND2xp5_ASAP7_75t_L g9895 ( 
.A(n_9499),
.B(n_5966),
.Y(n_9895)
);

AOI22xp5_ASAP7_75t_L g9896 ( 
.A1(n_9420),
.A2(n_6178),
.B1(n_6180),
.B2(n_6176),
.Y(n_9896)
);

NOR3xp33_ASAP7_75t_L g9897 ( 
.A(n_9364),
.B(n_9416),
.C(n_9205),
.Y(n_9897)
);

INVx2_ASAP7_75t_L g9898 ( 
.A(n_9649),
.Y(n_9898)
);

NAND2xp5_ASAP7_75t_L g9899 ( 
.A(n_9505),
.B(n_5967),
.Y(n_9899)
);

NOR2xp33_ASAP7_75t_L g9900 ( 
.A(n_9353),
.B(n_6182),
.Y(n_9900)
);

INVx2_ASAP7_75t_L g9901 ( 
.A(n_9652),
.Y(n_9901)
);

AOI22xp33_ASAP7_75t_L g9902 ( 
.A1(n_9461),
.A2(n_5979),
.B1(n_5984),
.B2(n_5976),
.Y(n_9902)
);

INVx3_ASAP7_75t_L g9903 ( 
.A(n_9490),
.Y(n_9903)
);

INVx1_ASAP7_75t_L g9904 ( 
.A(n_9510),
.Y(n_9904)
);

INVx1_ASAP7_75t_L g9905 ( 
.A(n_9518),
.Y(n_9905)
);

NAND2xp5_ASAP7_75t_L g9906 ( 
.A(n_9521),
.B(n_5985),
.Y(n_9906)
);

OR2x6_ASAP7_75t_L g9907 ( 
.A(n_9583),
.B(n_5997),
.Y(n_9907)
);

NAND2xp5_ASAP7_75t_L g9908 ( 
.A(n_9522),
.B(n_9523),
.Y(n_9908)
);

NOR2xp67_ASAP7_75t_L g9909 ( 
.A(n_9599),
.B(n_4338),
.Y(n_9909)
);

INVx1_ASAP7_75t_L g9910 ( 
.A(n_9535),
.Y(n_9910)
);

INVx1_ASAP7_75t_L g9911 ( 
.A(n_9536),
.Y(n_9911)
);

NAND2xp5_ASAP7_75t_L g9912 ( 
.A(n_9539),
.B(n_5999),
.Y(n_9912)
);

NOR2xp33_ASAP7_75t_L g9913 ( 
.A(n_9373),
.B(n_6183),
.Y(n_9913)
);

INVx3_ASAP7_75t_L g9914 ( 
.A(n_9490),
.Y(n_9914)
);

NAND2xp5_ASAP7_75t_SL g9915 ( 
.A(n_9597),
.B(n_6188),
.Y(n_9915)
);

NAND2xp5_ASAP7_75t_L g9916 ( 
.A(n_9559),
.B(n_6001),
.Y(n_9916)
);

NAND2xp5_ASAP7_75t_L g9917 ( 
.A(n_9560),
.B(n_6004),
.Y(n_9917)
);

NAND2xp5_ASAP7_75t_L g9918 ( 
.A(n_9203),
.B(n_6005),
.Y(n_9918)
);

HB1xp67_ASAP7_75t_L g9919 ( 
.A(n_9267),
.Y(n_9919)
);

NAND2xp5_ASAP7_75t_SL g9920 ( 
.A(n_9311),
.B(n_6191),
.Y(n_9920)
);

AND2x2_ASAP7_75t_L g9921 ( 
.A(n_9442),
.B(n_6197),
.Y(n_9921)
);

NAND2xp33_ASAP7_75t_L g9922 ( 
.A(n_9487),
.B(n_6201),
.Y(n_9922)
);

NOR2xp33_ASAP7_75t_L g9923 ( 
.A(n_9415),
.B(n_6203),
.Y(n_9923)
);

NAND2xp5_ASAP7_75t_SL g9924 ( 
.A(n_9485),
.B(n_6208),
.Y(n_9924)
);

INVx2_ASAP7_75t_L g9925 ( 
.A(n_9657),
.Y(n_9925)
);

NAND2xp5_ASAP7_75t_SL g9926 ( 
.A(n_9469),
.B(n_6215),
.Y(n_9926)
);

AND2x2_ASAP7_75t_L g9927 ( 
.A(n_9489),
.B(n_6216),
.Y(n_9927)
);

NAND2xp5_ASAP7_75t_L g9928 ( 
.A(n_9207),
.B(n_6013),
.Y(n_9928)
);

INVx2_ASAP7_75t_L g9929 ( 
.A(n_9661),
.Y(n_9929)
);

INVxp67_ASAP7_75t_L g9930 ( 
.A(n_9438),
.Y(n_9930)
);

NAND2xp5_ASAP7_75t_L g9931 ( 
.A(n_9208),
.B(n_6014),
.Y(n_9931)
);

INVxp67_ASAP7_75t_L g9932 ( 
.A(n_9445),
.Y(n_9932)
);

INVx1_ASAP7_75t_L g9933 ( 
.A(n_9197),
.Y(n_9933)
);

NAND2xp5_ASAP7_75t_SL g9934 ( 
.A(n_9653),
.B(n_6217),
.Y(n_9934)
);

INVx2_ASAP7_75t_SL g9935 ( 
.A(n_9195),
.Y(n_9935)
);

AND2x2_ASAP7_75t_L g9936 ( 
.A(n_9475),
.B(n_6219),
.Y(n_9936)
);

AND2x2_ASAP7_75t_L g9937 ( 
.A(n_9482),
.B(n_6221),
.Y(n_9937)
);

NAND2xp5_ASAP7_75t_L g9938 ( 
.A(n_9222),
.B(n_6015),
.Y(n_9938)
);

NAND2xp5_ASAP7_75t_SL g9939 ( 
.A(n_9660),
.B(n_6222),
.Y(n_9939)
);

INVx2_ASAP7_75t_L g9940 ( 
.A(n_9664),
.Y(n_9940)
);

AND2x4_ASAP7_75t_L g9941 ( 
.A(n_9568),
.B(n_6022),
.Y(n_9941)
);

OAI22xp5_ASAP7_75t_L g9942 ( 
.A1(n_9676),
.A2(n_6226),
.B1(n_6228),
.B2(n_6225),
.Y(n_9942)
);

NAND2xp5_ASAP7_75t_L g9943 ( 
.A(n_9245),
.B(n_6023),
.Y(n_9943)
);

INVx2_ASAP7_75t_L g9944 ( 
.A(n_9678),
.Y(n_9944)
);

INVxp33_ASAP7_75t_L g9945 ( 
.A(n_9444),
.Y(n_9945)
);

NAND2xp5_ASAP7_75t_L g9946 ( 
.A(n_9253),
.B(n_6030),
.Y(n_9946)
);

INVx2_ASAP7_75t_L g9947 ( 
.A(n_9680),
.Y(n_9947)
);

NAND2xp5_ASAP7_75t_L g9948 ( 
.A(n_9260),
.B(n_6033),
.Y(n_9948)
);

NAND2xp5_ASAP7_75t_L g9949 ( 
.A(n_9546),
.B(n_6036),
.Y(n_9949)
);

NAND2xp5_ASAP7_75t_L g9950 ( 
.A(n_9553),
.B(n_6039),
.Y(n_9950)
);

NAND2xp5_ASAP7_75t_SL g9951 ( 
.A(n_9684),
.B(n_6232),
.Y(n_9951)
);

OR2x2_ASAP7_75t_L g9952 ( 
.A(n_9567),
.B(n_6233),
.Y(n_9952)
);

BUFx5_ASAP7_75t_L g9953 ( 
.A(n_9683),
.Y(n_9953)
);

NAND2x1_ASAP7_75t_L g9954 ( 
.A(n_9200),
.B(n_6043),
.Y(n_9954)
);

NAND2xp5_ASAP7_75t_L g9955 ( 
.A(n_9561),
.B(n_9566),
.Y(n_9955)
);

INVx1_ASAP7_75t_L g9956 ( 
.A(n_9265),
.Y(n_9956)
);

NAND2xp5_ASAP7_75t_SL g9957 ( 
.A(n_9479),
.B(n_6237),
.Y(n_9957)
);

NOR2xp33_ASAP7_75t_L g9958 ( 
.A(n_9227),
.B(n_6240),
.Y(n_9958)
);

INVxp67_ASAP7_75t_L g9959 ( 
.A(n_9600),
.Y(n_9959)
);

OAI221xp5_ASAP7_75t_L g9960 ( 
.A1(n_9503),
.A2(n_6057),
.B1(n_6065),
.B2(n_6053),
.C(n_6051),
.Y(n_9960)
);

NOR2xp67_ASAP7_75t_L g9961 ( 
.A(n_9601),
.B(n_4339),
.Y(n_9961)
);

NAND2xp5_ASAP7_75t_L g9962 ( 
.A(n_9584),
.B(n_6066),
.Y(n_9962)
);

BUFx8_ASAP7_75t_L g9963 ( 
.A(n_9576),
.Y(n_9963)
);

NOR2xp67_ASAP7_75t_L g9964 ( 
.A(n_9602),
.B(n_4340),
.Y(n_9964)
);

NAND2xp5_ASAP7_75t_L g9965 ( 
.A(n_9593),
.B(n_6067),
.Y(n_9965)
);

OAI22xp5_ASAP7_75t_L g9966 ( 
.A1(n_9633),
.A2(n_6245),
.B1(n_6246),
.B2(n_6242),
.Y(n_9966)
);

NAND2xp5_ASAP7_75t_L g9967 ( 
.A(n_9594),
.B(n_6070),
.Y(n_9967)
);

INVx2_ASAP7_75t_L g9968 ( 
.A(n_9278),
.Y(n_9968)
);

NAND2xp5_ASAP7_75t_L g9969 ( 
.A(n_9612),
.B(n_9619),
.Y(n_9969)
);

BUFx3_ASAP7_75t_L g9970 ( 
.A(n_9313),
.Y(n_9970)
);

NAND2xp5_ASAP7_75t_L g9971 ( 
.A(n_9625),
.B(n_6077),
.Y(n_9971)
);

BUFx3_ASAP7_75t_L g9972 ( 
.A(n_9318),
.Y(n_9972)
);

INVx2_ASAP7_75t_L g9973 ( 
.A(n_9279),
.Y(n_9973)
);

INVx2_ASAP7_75t_L g9974 ( 
.A(n_9562),
.Y(n_9974)
);

BUFx6f_ASAP7_75t_SL g9975 ( 
.A(n_9372),
.Y(n_9975)
);

NAND2xp5_ASAP7_75t_L g9976 ( 
.A(n_9564),
.B(n_6078),
.Y(n_9976)
);

NOR2xp33_ASAP7_75t_L g9977 ( 
.A(n_9607),
.B(n_6248),
.Y(n_9977)
);

INVx2_ASAP7_75t_L g9978 ( 
.A(n_9569),
.Y(n_9978)
);

INVx1_ASAP7_75t_L g9979 ( 
.A(n_9604),
.Y(n_9979)
);

NAND2xp5_ASAP7_75t_SL g9980 ( 
.A(n_9679),
.B(n_6249),
.Y(n_9980)
);

NAND2xp5_ASAP7_75t_L g9981 ( 
.A(n_9611),
.B(n_6079),
.Y(n_9981)
);

CKINVDCx5p33_ASAP7_75t_R g9982 ( 
.A(n_9508),
.Y(n_9982)
);

INVx1_ASAP7_75t_L g9983 ( 
.A(n_9616),
.Y(n_9983)
);

NAND2xp5_ASAP7_75t_L g9984 ( 
.A(n_9622),
.B(n_6088),
.Y(n_9984)
);

NOR2xp33_ASAP7_75t_L g9985 ( 
.A(n_9549),
.B(n_6252),
.Y(n_9985)
);

AND2x4_ASAP7_75t_L g9986 ( 
.A(n_9571),
.B(n_6089),
.Y(n_9986)
);

INVx2_ASAP7_75t_L g9987 ( 
.A(n_9626),
.Y(n_9987)
);

AND2x2_ASAP7_75t_L g9988 ( 
.A(n_9506),
.B(n_6254),
.Y(n_9988)
);

NAND2xp5_ASAP7_75t_L g9989 ( 
.A(n_9637),
.B(n_6094),
.Y(n_9989)
);

NAND2xp5_ASAP7_75t_L g9990 ( 
.A(n_9681),
.B(n_6096),
.Y(n_9990)
);

NOR3xp33_ASAP7_75t_L g9991 ( 
.A(n_9538),
.B(n_6101),
.C(n_6099),
.Y(n_9991)
);

NAND2xp5_ASAP7_75t_L g9992 ( 
.A(n_9381),
.B(n_6107),
.Y(n_9992)
);

OAI22xp33_ASAP7_75t_L g9993 ( 
.A1(n_9685),
.A2(n_6258),
.B1(n_6265),
.B2(n_6256),
.Y(n_9993)
);

NOR2xp33_ASAP7_75t_L g9994 ( 
.A(n_9280),
.B(n_6271),
.Y(n_9994)
);

INVx4_ASAP7_75t_L g9995 ( 
.A(n_9195),
.Y(n_9995)
);

AOI22xp33_ASAP7_75t_L g9996 ( 
.A1(n_9461),
.A2(n_6113),
.B1(n_6114),
.B2(n_6108),
.Y(n_9996)
);

INVx2_ASAP7_75t_L g9997 ( 
.A(n_9286),
.Y(n_9997)
);

NAND2xp5_ASAP7_75t_L g9998 ( 
.A(n_9383),
.B(n_6116),
.Y(n_9998)
);

NOR2xp33_ASAP7_75t_L g9999 ( 
.A(n_9492),
.B(n_6272),
.Y(n_9999)
);

NAND3xp33_ASAP7_75t_L g10000 ( 
.A(n_9430),
.B(n_9238),
.C(n_9288),
.Y(n_10000)
);

INVx2_ASAP7_75t_L g10001 ( 
.A(n_9294),
.Y(n_10001)
);

NAND2xp5_ASAP7_75t_L g10002 ( 
.A(n_9414),
.B(n_6121),
.Y(n_10002)
);

NOR2xp33_ASAP7_75t_L g10003 ( 
.A(n_9470),
.B(n_9333),
.Y(n_10003)
);

BUFx6f_ASAP7_75t_SL g10004 ( 
.A(n_9190),
.Y(n_10004)
);

INVx2_ASAP7_75t_L g10005 ( 
.A(n_9295),
.Y(n_10005)
);

AOI221xp5_ASAP7_75t_L g10006 ( 
.A1(n_9417),
.A2(n_6132),
.B1(n_6137),
.B2(n_6129),
.C(n_6125),
.Y(n_10006)
);

INVx2_ASAP7_75t_L g10007 ( 
.A(n_9296),
.Y(n_10007)
);

NAND2xp5_ASAP7_75t_L g10008 ( 
.A(n_9421),
.B(n_6141),
.Y(n_10008)
);

NAND2xp5_ASAP7_75t_L g10009 ( 
.A(n_9434),
.B(n_6144),
.Y(n_10009)
);

INVx2_ASAP7_75t_L g10010 ( 
.A(n_9299),
.Y(n_10010)
);

NOR2xp33_ASAP7_75t_L g10011 ( 
.A(n_9673),
.B(n_6273),
.Y(n_10011)
);

AOI22xp33_ASAP7_75t_L g10012 ( 
.A1(n_9662),
.A2(n_6147),
.B1(n_6154),
.B2(n_6146),
.Y(n_10012)
);

AND2x4_ASAP7_75t_L g10013 ( 
.A(n_9573),
.B(n_6155),
.Y(n_10013)
);

OA22x2_ASAP7_75t_L g10014 ( 
.A1(n_9556),
.A2(n_6276),
.B1(n_6277),
.B2(n_6274),
.Y(n_10014)
);

INVx4_ASAP7_75t_L g10015 ( 
.A(n_9231),
.Y(n_10015)
);

NAND2xp5_ASAP7_75t_L g10016 ( 
.A(n_9448),
.B(n_6159),
.Y(n_10016)
);

INVx1_ASAP7_75t_L g10017 ( 
.A(n_9281),
.Y(n_10017)
);

INVx2_ASAP7_75t_L g10018 ( 
.A(n_9302),
.Y(n_10018)
);

NAND2xp5_ASAP7_75t_L g10019 ( 
.A(n_9315),
.B(n_9317),
.Y(n_10019)
);

INVx2_ASAP7_75t_L g10020 ( 
.A(n_9328),
.Y(n_10020)
);

BUFx3_ASAP7_75t_L g10021 ( 
.A(n_9368),
.Y(n_10021)
);

NAND2xp5_ASAP7_75t_SL g10022 ( 
.A(n_9641),
.B(n_6278),
.Y(n_10022)
);

NAND2xp5_ASAP7_75t_L g10023 ( 
.A(n_9330),
.B(n_9336),
.Y(n_10023)
);

OAI22xp5_ASAP7_75t_L g10024 ( 
.A1(n_9344),
.A2(n_6285),
.B1(n_6286),
.B2(n_6279),
.Y(n_10024)
);

BUFx8_ASAP7_75t_L g10025 ( 
.A(n_9511),
.Y(n_10025)
);

AOI22xp33_ASAP7_75t_L g10026 ( 
.A1(n_9636),
.A2(n_6163),
.B1(n_6164),
.B2(n_6162),
.Y(n_10026)
);

NAND2xp5_ASAP7_75t_L g10027 ( 
.A(n_9356),
.B(n_6177),
.Y(n_10027)
);

NAND2xp5_ASAP7_75t_SL g10028 ( 
.A(n_9641),
.B(n_6289),
.Y(n_10028)
);

INVxp67_ASAP7_75t_L g10029 ( 
.A(n_9231),
.Y(n_10029)
);

AOI22xp5_ASAP7_75t_L g10030 ( 
.A1(n_9384),
.A2(n_6292),
.B1(n_6293),
.B2(n_6290),
.Y(n_10030)
);

NAND2xp5_ASAP7_75t_L g10031 ( 
.A(n_9358),
.B(n_6184),
.Y(n_10031)
);

NAND2xp5_ASAP7_75t_SL g10032 ( 
.A(n_9575),
.B(n_6294),
.Y(n_10032)
);

NAND2xp5_ASAP7_75t_SL g10033 ( 
.A(n_9575),
.B(n_6296),
.Y(n_10033)
);

AOI22xp33_ASAP7_75t_L g10034 ( 
.A1(n_9645),
.A2(n_6186),
.B1(n_6187),
.B2(n_6185),
.Y(n_10034)
);

BUFx6f_ASAP7_75t_L g10035 ( 
.A(n_9261),
.Y(n_10035)
);

INVxp67_ASAP7_75t_L g10036 ( 
.A(n_9261),
.Y(n_10036)
);

NOR2xp33_ASAP7_75t_L g10037 ( 
.A(n_9632),
.B(n_6300),
.Y(n_10037)
);

INVx2_ASAP7_75t_SL g10038 ( 
.A(n_9268),
.Y(n_10038)
);

NAND2xp5_ASAP7_75t_L g10039 ( 
.A(n_9370),
.B(n_6189),
.Y(n_10039)
);

NAND2xp5_ASAP7_75t_L g10040 ( 
.A(n_9375),
.B(n_6190),
.Y(n_10040)
);

AND2x2_ASAP7_75t_L g10041 ( 
.A(n_9646),
.B(n_6303),
.Y(n_10041)
);

INVx4_ASAP7_75t_L g10042 ( 
.A(n_9268),
.Y(n_10042)
);

INVx8_ASAP7_75t_L g10043 ( 
.A(n_9284),
.Y(n_10043)
);

INVx2_ASAP7_75t_L g10044 ( 
.A(n_9376),
.Y(n_10044)
);

NAND2xp5_ASAP7_75t_L g10045 ( 
.A(n_9385),
.B(n_6192),
.Y(n_10045)
);

O2A1O1Ixp33_ASAP7_75t_L g10046 ( 
.A1(n_9540),
.A2(n_6196),
.B(n_6199),
.C(n_6194),
.Y(n_10046)
);

NAND2xp5_ASAP7_75t_L g10047 ( 
.A(n_9386),
.B(n_9390),
.Y(n_10047)
);

NAND2xp5_ASAP7_75t_L g10048 ( 
.A(n_9391),
.B(n_6200),
.Y(n_10048)
);

AND2x6_ASAP7_75t_SL g10049 ( 
.A(n_9187),
.B(n_6206),
.Y(n_10049)
);

INVx1_ASAP7_75t_L g10050 ( 
.A(n_9394),
.Y(n_10050)
);

INVx2_ASAP7_75t_SL g10051 ( 
.A(n_9284),
.Y(n_10051)
);

INVx1_ASAP7_75t_L g10052 ( 
.A(n_9411),
.Y(n_10052)
);

NAND2xp5_ASAP7_75t_L g10053 ( 
.A(n_9431),
.B(n_6210),
.Y(n_10053)
);

INVx2_ASAP7_75t_L g10054 ( 
.A(n_9436),
.Y(n_10054)
);

INVx1_ASAP7_75t_L g10055 ( 
.A(n_9450),
.Y(n_10055)
);

AND2x2_ASAP7_75t_L g10056 ( 
.A(n_9672),
.B(n_6304),
.Y(n_10056)
);

INVx2_ASAP7_75t_L g10057 ( 
.A(n_9466),
.Y(n_10057)
);

INVx1_ASAP7_75t_L g10058 ( 
.A(n_9483),
.Y(n_10058)
);

NOR2xp33_ASAP7_75t_L g10059 ( 
.A(n_9500),
.B(n_6309),
.Y(n_10059)
);

NOR2xp33_ASAP7_75t_L g10060 ( 
.A(n_9579),
.B(n_9644),
.Y(n_10060)
);

NAND2xp5_ASAP7_75t_L g10061 ( 
.A(n_9497),
.B(n_6212),
.Y(n_10061)
);

AO22x2_ASAP7_75t_L g10062 ( 
.A1(n_9638),
.A2(n_6214),
.B1(n_6223),
.B2(n_6213),
.Y(n_10062)
);

INVx1_ASAP7_75t_L g10063 ( 
.A(n_9655),
.Y(n_10063)
);

INVx2_ASAP7_75t_L g10064 ( 
.A(n_9656),
.Y(n_10064)
);

NAND2xp5_ASAP7_75t_L g10065 ( 
.A(n_9668),
.B(n_6224),
.Y(n_10065)
);

INVx1_ASAP7_75t_L g10066 ( 
.A(n_9614),
.Y(n_10066)
);

AOI22xp33_ASAP7_75t_L g10067 ( 
.A1(n_9645),
.A2(n_6229),
.B1(n_6231),
.B2(n_6227),
.Y(n_10067)
);

NOR3xp33_ASAP7_75t_L g10068 ( 
.A(n_9354),
.B(n_6244),
.C(n_6236),
.Y(n_10068)
);

NAND2xp5_ASAP7_75t_L g10069 ( 
.A(n_9663),
.B(n_6247),
.Y(n_10069)
);

AOI22xp5_ASAP7_75t_L g10070 ( 
.A1(n_9627),
.A2(n_6312),
.B1(n_6317),
.B2(n_6311),
.Y(n_10070)
);

AOI22xp5_ASAP7_75t_L g10071 ( 
.A1(n_9220),
.A2(n_6322),
.B1(n_6324),
.B2(n_6321),
.Y(n_10071)
);

NAND2xp5_ASAP7_75t_L g10072 ( 
.A(n_9287),
.B(n_6251),
.Y(n_10072)
);

BUFx3_ASAP7_75t_L g10073 ( 
.A(n_9393),
.Y(n_10073)
);

NAND2xp5_ASAP7_75t_SL g10074 ( 
.A(n_9292),
.B(n_6326),
.Y(n_10074)
);

NAND2xp5_ASAP7_75t_L g10075 ( 
.A(n_9487),
.B(n_9578),
.Y(n_10075)
);

NAND2xp5_ASAP7_75t_L g10076 ( 
.A(n_9589),
.B(n_9658),
.Y(n_10076)
);

NOR2xp67_ASAP7_75t_L g10077 ( 
.A(n_9651),
.B(n_4341),
.Y(n_10077)
);

NAND2xp5_ASAP7_75t_SL g10078 ( 
.A(n_9292),
.B(n_6327),
.Y(n_10078)
);

O2A1O1Ixp33_ASAP7_75t_L g10079 ( 
.A1(n_9598),
.A2(n_6255),
.B(n_6259),
.C(n_6253),
.Y(n_10079)
);

AND2x4_ASAP7_75t_L g10080 ( 
.A(n_9467),
.B(n_6262),
.Y(n_10080)
);

NAND2xp5_ASAP7_75t_SL g10081 ( 
.A(n_9341),
.B(n_6331),
.Y(n_10081)
);

INVx1_ASAP7_75t_L g10082 ( 
.A(n_9618),
.Y(n_10082)
);

AND2x2_ASAP7_75t_L g10083 ( 
.A(n_9230),
.B(n_6332),
.Y(n_10083)
);

AND2x2_ASAP7_75t_L g10084 ( 
.A(n_9587),
.B(n_6339),
.Y(n_10084)
);

BUFx6f_ASAP7_75t_SL g10085 ( 
.A(n_9226),
.Y(n_10085)
);

INVx2_ASAP7_75t_SL g10086 ( 
.A(n_9341),
.Y(n_10086)
);

NAND2xp5_ASAP7_75t_L g10087 ( 
.A(n_9557),
.B(n_6266),
.Y(n_10087)
);

NOR2xp67_ASAP7_75t_L g10088 ( 
.A(n_9528),
.B(n_4342),
.Y(n_10088)
);

AOI22xp5_ASAP7_75t_L g10089 ( 
.A1(n_9659),
.A2(n_6342),
.B1(n_6343),
.B2(n_6340),
.Y(n_10089)
);

NAND2xp5_ASAP7_75t_L g10090 ( 
.A(n_9557),
.B(n_6267),
.Y(n_10090)
);

AOI22xp5_ASAP7_75t_L g10091 ( 
.A1(n_9623),
.A2(n_6351),
.B1(n_6352),
.B2(n_6349),
.Y(n_10091)
);

AND2x6_ASAP7_75t_SL g10092 ( 
.A(n_9617),
.B(n_6268),
.Y(n_10092)
);

NAND2xp5_ASAP7_75t_SL g10093 ( 
.A(n_9342),
.B(n_6359),
.Y(n_10093)
);

NAND3xp33_ASAP7_75t_L g10094 ( 
.A(n_9357),
.B(n_6366),
.C(n_6363),
.Y(n_10094)
);

NAND2xp5_ASAP7_75t_L g10095 ( 
.A(n_9570),
.B(n_6269),
.Y(n_10095)
);

A2O1A1Ixp33_ASAP7_75t_L g10096 ( 
.A1(n_9647),
.A2(n_6287),
.B(n_6302),
.C(n_6284),
.Y(n_10096)
);

NAND2xp5_ASAP7_75t_SL g10097 ( 
.A(n_9342),
.B(n_6370),
.Y(n_10097)
);

BUFx6f_ASAP7_75t_L g10098 ( 
.A(n_9352),
.Y(n_10098)
);

NAND2xp5_ASAP7_75t_L g10099 ( 
.A(n_9570),
.B(n_6305),
.Y(n_10099)
);

NAND2xp5_ASAP7_75t_SL g10100 ( 
.A(n_9352),
.B(n_6376),
.Y(n_10100)
);

O2A1O1Ixp33_ASAP7_75t_L g10101 ( 
.A1(n_9504),
.A2(n_9525),
.B(n_9404),
.C(n_9418),
.Y(n_10101)
);

NOR2xp33_ASAP7_75t_L g10102 ( 
.A(n_9581),
.B(n_6377),
.Y(n_10102)
);

NAND2xp5_ASAP7_75t_L g10103 ( 
.A(n_9603),
.B(n_6310),
.Y(n_10103)
);

NOR2xp67_ASAP7_75t_L g10104 ( 
.A(n_9472),
.B(n_4343),
.Y(n_10104)
);

BUFx3_ASAP7_75t_L g10105 ( 
.A(n_9396),
.Y(n_10105)
);

INVxp67_ASAP7_75t_L g10106 ( 
.A(n_9365),
.Y(n_10106)
);

HB1xp67_ASAP7_75t_L g10107 ( 
.A(n_9451),
.Y(n_10107)
);

AND2x6_ASAP7_75t_SL g10108 ( 
.A(n_9446),
.B(n_6315),
.Y(n_10108)
);

INVx2_ASAP7_75t_L g10109 ( 
.A(n_9550),
.Y(n_10109)
);

INVx2_ASAP7_75t_L g10110 ( 
.A(n_9677),
.Y(n_10110)
);

NAND2xp5_ASAP7_75t_SL g10111 ( 
.A(n_9365),
.B(n_6378),
.Y(n_10111)
);

AND2x2_ASAP7_75t_L g10112 ( 
.A(n_9630),
.B(n_6379),
.Y(n_10112)
);

NAND2xp5_ASAP7_75t_SL g10113 ( 
.A(n_9371),
.B(n_9399),
.Y(n_10113)
);

INVx1_ASAP7_75t_L g10114 ( 
.A(n_9449),
.Y(n_10114)
);

NAND2xp5_ASAP7_75t_L g10115 ( 
.A(n_9623),
.B(n_6316),
.Y(n_10115)
);

INVx1_ASAP7_75t_L g10116 ( 
.A(n_9464),
.Y(n_10116)
);

OR2x6_ASAP7_75t_L g10117 ( 
.A(n_9283),
.B(n_9291),
.Y(n_10117)
);

NOR2xp33_ASAP7_75t_L g10118 ( 
.A(n_9551),
.B(n_6385),
.Y(n_10118)
);

INVx1_ASAP7_75t_L g10119 ( 
.A(n_9465),
.Y(n_10119)
);

INVx2_ASAP7_75t_SL g10120 ( 
.A(n_9371),
.Y(n_10120)
);

NAND2xp5_ASAP7_75t_SL g10121 ( 
.A(n_9399),
.B(n_6387),
.Y(n_10121)
);

NAND2xp5_ASAP7_75t_L g10122 ( 
.A(n_9574),
.B(n_6318),
.Y(n_10122)
);

NAND2xp5_ASAP7_75t_SL g10123 ( 
.A(n_9409),
.B(n_6388),
.Y(n_10123)
);

INVx2_ASAP7_75t_L g10124 ( 
.A(n_9610),
.Y(n_10124)
);

NAND2xp5_ASAP7_75t_SL g10125 ( 
.A(n_9409),
.B(n_6389),
.Y(n_10125)
);

INVx1_ASAP7_75t_L g10126 ( 
.A(n_9478),
.Y(n_10126)
);

NOR2xp33_ASAP7_75t_L g10127 ( 
.A(n_9620),
.B(n_6391),
.Y(n_10127)
);

NAND2xp5_ASAP7_75t_L g10128 ( 
.A(n_9514),
.B(n_9537),
.Y(n_10128)
);

INVx2_ASAP7_75t_L g10129 ( 
.A(n_9667),
.Y(n_10129)
);

NAND2xp5_ASAP7_75t_SL g10130 ( 
.A(n_9425),
.B(n_6392),
.Y(n_10130)
);

INVx1_ASAP7_75t_SL g10131 ( 
.A(n_9669),
.Y(n_10131)
);

NAND2xp5_ASAP7_75t_SL g10132 ( 
.A(n_9425),
.B(n_6393),
.Y(n_10132)
);

INVx8_ASAP7_75t_L g10133 ( 
.A(n_9511),
.Y(n_10133)
);

NAND2xp5_ASAP7_75t_L g10134 ( 
.A(n_9621),
.B(n_6333),
.Y(n_10134)
);

NAND2xp5_ASAP7_75t_L g10135 ( 
.A(n_9634),
.B(n_6337),
.Y(n_10135)
);

NAND2xp5_ASAP7_75t_L g10136 ( 
.A(n_9229),
.B(n_6348),
.Y(n_10136)
);

NAND2xp5_ASAP7_75t_L g10137 ( 
.A(n_9229),
.B(n_6350),
.Y(n_10137)
);

OR2x2_ASAP7_75t_L g10138 ( 
.A(n_9247),
.B(n_6394),
.Y(n_10138)
);

AOI221xp5_ASAP7_75t_L g10139 ( 
.A1(n_9543),
.A2(n_9422),
.B1(n_9447),
.B2(n_9388),
.C(n_6364),
.Y(n_10139)
);

NAND2xp5_ASAP7_75t_L g10140 ( 
.A(n_9251),
.B(n_6355),
.Y(n_10140)
);

AOI22xp33_ASAP7_75t_L g10141 ( 
.A1(n_9534),
.A2(n_6367),
.B1(n_6371),
.B2(n_6360),
.Y(n_10141)
);

NOR2xp33_ASAP7_75t_L g10142 ( 
.A(n_9319),
.B(n_6395),
.Y(n_10142)
);

NAND2xp5_ASAP7_75t_SL g10143 ( 
.A(n_9643),
.B(n_6397),
.Y(n_10143)
);

AND2x2_ASAP7_75t_L g10144 ( 
.A(n_9329),
.B(n_6398),
.Y(n_10144)
);

INVx2_ASAP7_75t_L g10145 ( 
.A(n_9255),
.Y(n_10145)
);

NAND2xp5_ASAP7_75t_SL g10146 ( 
.A(n_9346),
.B(n_6401),
.Y(n_10146)
);

NOR2xp33_ASAP7_75t_L g10147 ( 
.A(n_9355),
.B(n_6402),
.Y(n_10147)
);

NAND2xp5_ASAP7_75t_SL g10148 ( 
.A(n_9366),
.B(n_6404),
.Y(n_10148)
);

NAND2xp5_ASAP7_75t_SL g10149 ( 
.A(n_9369),
.B(n_6411),
.Y(n_10149)
);

NAND2xp5_ASAP7_75t_L g10150 ( 
.A(n_9251),
.B(n_6372),
.Y(n_10150)
);

NOR2xp67_ASAP7_75t_L g10151 ( 
.A(n_9378),
.B(n_4344),
.Y(n_10151)
);

INVx1_ASAP7_75t_L g10152 ( 
.A(n_9332),
.Y(n_10152)
);

INVx1_ASAP7_75t_L g10153 ( 
.A(n_9349),
.Y(n_10153)
);

NAND2xp5_ASAP7_75t_SL g10154 ( 
.A(n_9379),
.B(n_6412),
.Y(n_10154)
);

NAND2xp5_ASAP7_75t_L g10155 ( 
.A(n_9387),
.B(n_6373),
.Y(n_10155)
);

INVx8_ASAP7_75t_L g10156 ( 
.A(n_9439),
.Y(n_10156)
);

INVx2_ASAP7_75t_L g10157 ( 
.A(n_9516),
.Y(n_10157)
);

NAND2xp5_ASAP7_75t_SL g10158 ( 
.A(n_9382),
.B(n_9389),
.Y(n_10158)
);

NAND2xp5_ASAP7_75t_SL g10159 ( 
.A(n_9392),
.B(n_6374),
.Y(n_10159)
);

NAND2xp5_ASAP7_75t_L g10160 ( 
.A(n_9387),
.B(n_6381),
.Y(n_10160)
);

INVx1_ASAP7_75t_L g10161 ( 
.A(n_9194),
.Y(n_10161)
);

NAND2xp5_ASAP7_75t_L g10162 ( 
.A(n_9432),
.B(n_6382),
.Y(n_10162)
);

INVx2_ASAP7_75t_L g10163 ( 
.A(n_9517),
.Y(n_10163)
);

NAND2xp5_ASAP7_75t_SL g10164 ( 
.A(n_9410),
.B(n_6390),
.Y(n_10164)
);

NOR2xp33_ASAP7_75t_L g10165 ( 
.A(n_9565),
.B(n_6405),
.Y(n_10165)
);

NAND2xp5_ASAP7_75t_SL g10166 ( 
.A(n_9240),
.B(n_6406),
.Y(n_10166)
);

AND2x2_ASAP7_75t_L g10167 ( 
.A(n_9552),
.B(n_6409),
.Y(n_10167)
);

INVx1_ASAP7_75t_L g10168 ( 
.A(n_9398),
.Y(n_10168)
);

INVx1_ASAP7_75t_L g10169 ( 
.A(n_9408),
.Y(n_10169)
);

AND2x2_ASAP7_75t_L g10170 ( 
.A(n_9256),
.B(n_6415),
.Y(n_10170)
);

INVx2_ASAP7_75t_L g10171 ( 
.A(n_9530),
.Y(n_10171)
);

NOR2xp33_ASAP7_75t_L g10172 ( 
.A(n_9532),
.B(n_6416),
.Y(n_10172)
);

AND2x2_ASAP7_75t_L g10173 ( 
.A(n_9426),
.B(n_6008),
.Y(n_10173)
);

NAND2xp5_ASAP7_75t_SL g10174 ( 
.A(n_9452),
.B(n_6016),
.Y(n_10174)
);

INVx2_ASAP7_75t_L g10175 ( 
.A(n_9441),
.Y(n_10175)
);

NOR2xp33_ASAP7_75t_L g10176 ( 
.A(n_9582),
.B(n_9572),
.Y(n_10176)
);

AND2x4_ASAP7_75t_L g10177 ( 
.A(n_9271),
.B(n_4345),
.Y(n_10177)
);

NAND2xp5_ASAP7_75t_L g10178 ( 
.A(n_9432),
.B(n_6027),
.Y(n_10178)
);

NAND2xp5_ASAP7_75t_L g10179 ( 
.A(n_9640),
.B(n_6050),
.Y(n_10179)
);

NOR3xp33_ASAP7_75t_L g10180 ( 
.A(n_9226),
.B(n_6059),
.C(n_6055),
.Y(n_10180)
);

NAND2xp5_ASAP7_75t_SL g10181 ( 
.A(n_9254),
.B(n_6080),
.Y(n_10181)
);

A2O1A1Ixp33_ASAP7_75t_L g10182 ( 
.A1(n_9219),
.A2(n_6098),
.B(n_6198),
.C(n_6083),
.Y(n_10182)
);

NOR2xp33_ASAP7_75t_L g10183 ( 
.A(n_9272),
.B(n_6204),
.Y(n_10183)
);

INVx2_ASAP7_75t_L g10184 ( 
.A(n_9501),
.Y(n_10184)
);

AND2x2_ASAP7_75t_L g10185 ( 
.A(n_9237),
.B(n_6207),
.Y(n_10185)
);

AND2x2_ASAP7_75t_L g10186 ( 
.A(n_9237),
.B(n_6241),
.Y(n_10186)
);

NOR2xp33_ASAP7_75t_L g10187 ( 
.A(n_9272),
.B(n_6288),
.Y(n_10187)
);

AOI21xp5_ASAP7_75t_L g10188 ( 
.A1(n_9290),
.A2(n_6325),
.B(n_6297),
.Y(n_10188)
);

INVx1_ASAP7_75t_L g10189 ( 
.A(n_9185),
.Y(n_10189)
);

INVx1_ASAP7_75t_L g10190 ( 
.A(n_9185),
.Y(n_10190)
);

INVx1_ASAP7_75t_L g10191 ( 
.A(n_9185),
.Y(n_10191)
);

NAND2xp5_ASAP7_75t_L g10192 ( 
.A(n_9272),
.B(n_6338),
.Y(n_10192)
);

AOI22xp5_ASAP7_75t_L g10193 ( 
.A1(n_9209),
.A2(n_6407),
.B1(n_6440),
.B2(n_6368),
.Y(n_10193)
);

CKINVDCx5p33_ASAP7_75t_R g10194 ( 
.A(n_9204),
.Y(n_10194)
);

NAND2xp5_ASAP7_75t_L g10195 ( 
.A(n_9272),
.B(n_6482),
.Y(n_10195)
);

NAND2xp5_ASAP7_75t_SL g10196 ( 
.A(n_9272),
.B(n_4),
.Y(n_10196)
);

INVx1_ASAP7_75t_L g10197 ( 
.A(n_9185),
.Y(n_10197)
);

BUFx4f_ASAP7_75t_L g10198 ( 
.A(n_9412),
.Y(n_10198)
);

NAND2xp5_ASAP7_75t_SL g10199 ( 
.A(n_9272),
.B(n_4),
.Y(n_10199)
);

INVx2_ASAP7_75t_SL g10200 ( 
.A(n_9406),
.Y(n_10200)
);

AND2x2_ASAP7_75t_L g10201 ( 
.A(n_9237),
.B(n_5),
.Y(n_10201)
);

NOR2xp33_ASAP7_75t_L g10202 ( 
.A(n_9272),
.B(n_5),
.Y(n_10202)
);

INVx1_ASAP7_75t_L g10203 ( 
.A(n_9185),
.Y(n_10203)
);

NAND2xp5_ASAP7_75t_L g10204 ( 
.A(n_9272),
.B(n_6),
.Y(n_10204)
);

INVx2_ASAP7_75t_L g10205 ( 
.A(n_9501),
.Y(n_10205)
);

NAND2xp5_ASAP7_75t_L g10206 ( 
.A(n_9719),
.B(n_6),
.Y(n_10206)
);

INVx1_ASAP7_75t_L g10207 ( 
.A(n_9830),
.Y(n_10207)
);

INVx1_ASAP7_75t_L g10208 ( 
.A(n_9873),
.Y(n_10208)
);

OR2x6_ASAP7_75t_L g10209 ( 
.A(n_9747),
.B(n_4346),
.Y(n_10209)
);

NAND2xp5_ASAP7_75t_L g10210 ( 
.A(n_9696),
.B(n_7),
.Y(n_10210)
);

AO22x2_ASAP7_75t_L g10211 ( 
.A1(n_9701),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_10211)
);

INVx1_ASAP7_75t_L g10212 ( 
.A(n_9908),
.Y(n_10212)
);

INVx1_ASAP7_75t_L g10213 ( 
.A(n_9762),
.Y(n_10213)
);

AND2x2_ASAP7_75t_L g10214 ( 
.A(n_9687),
.B(n_10),
.Y(n_10214)
);

AND2x2_ASAP7_75t_L g10215 ( 
.A(n_9862),
.B(n_10167),
.Y(n_10215)
);

INVx1_ASAP7_75t_L g10216 ( 
.A(n_9766),
.Y(n_10216)
);

HB1xp67_ASAP7_75t_L g10217 ( 
.A(n_9694),
.Y(n_10217)
);

OR2x6_ASAP7_75t_L g10218 ( 
.A(n_9747),
.B(n_4347),
.Y(n_10218)
);

NAND2x1p5_ASAP7_75t_L g10219 ( 
.A(n_10198),
.B(n_4349),
.Y(n_10219)
);

INVx2_ASAP7_75t_L g10220 ( 
.A(n_9769),
.Y(n_10220)
);

NAND2xp5_ASAP7_75t_L g10221 ( 
.A(n_10060),
.B(n_11),
.Y(n_10221)
);

AO22x2_ASAP7_75t_L g10222 ( 
.A1(n_9789),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_10222)
);

NOR2xp33_ASAP7_75t_L g10223 ( 
.A(n_9691),
.B(n_4350),
.Y(n_10223)
);

INVx1_ASAP7_75t_L g10224 ( 
.A(n_9785),
.Y(n_10224)
);

NOR2xp33_ASAP7_75t_L g10225 ( 
.A(n_9945),
.B(n_4351),
.Y(n_10225)
);

OAI221xp5_ASAP7_75t_L g10226 ( 
.A1(n_9849),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.C(n_17),
.Y(n_10226)
);

AND2x4_ASAP7_75t_L g10227 ( 
.A(n_9823),
.B(n_9970),
.Y(n_10227)
);

INVx1_ASAP7_75t_L g10228 ( 
.A(n_9792),
.Y(n_10228)
);

NAND2xp5_ASAP7_75t_L g10229 ( 
.A(n_9793),
.B(n_9698),
.Y(n_10229)
);

INVx1_ASAP7_75t_L g10230 ( 
.A(n_9802),
.Y(n_10230)
);

INVx1_ASAP7_75t_L g10231 ( 
.A(n_9806),
.Y(n_10231)
);

INVxp67_ASAP7_75t_L g10232 ( 
.A(n_9689),
.Y(n_10232)
);

AO22x2_ASAP7_75t_L g10233 ( 
.A1(n_9711),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_10233)
);

INVx1_ASAP7_75t_L g10234 ( 
.A(n_9813),
.Y(n_10234)
);

AND2x4_ASAP7_75t_L g10235 ( 
.A(n_9972),
.B(n_4353),
.Y(n_10235)
);

INVx1_ASAP7_75t_L g10236 ( 
.A(n_9817),
.Y(n_10236)
);

INVx1_ASAP7_75t_L g10237 ( 
.A(n_9819),
.Y(n_10237)
);

NAND2x1p5_ASAP7_75t_L g10238 ( 
.A(n_9810),
.B(n_4354),
.Y(n_10238)
);

INVxp67_ASAP7_75t_L g10239 ( 
.A(n_9919),
.Y(n_10239)
);

INVx1_ASAP7_75t_L g10240 ( 
.A(n_9831),
.Y(n_10240)
);

NAND2xp5_ASAP7_75t_L g10241 ( 
.A(n_9749),
.B(n_18),
.Y(n_10241)
);

NOR2xp33_ASAP7_75t_L g10242 ( 
.A(n_9782),
.B(n_4355),
.Y(n_10242)
);

INVx1_ASAP7_75t_L g10243 ( 
.A(n_9832),
.Y(n_10243)
);

INVx1_ASAP7_75t_L g10244 ( 
.A(n_9836),
.Y(n_10244)
);

CKINVDCx5p33_ASAP7_75t_R g10245 ( 
.A(n_10194),
.Y(n_10245)
);

INVxp67_ASAP7_75t_L g10246 ( 
.A(n_10107),
.Y(n_10246)
);

AND2x4_ASAP7_75t_L g10247 ( 
.A(n_10021),
.B(n_4356),
.Y(n_10247)
);

INVx1_ASAP7_75t_L g10248 ( 
.A(n_9840),
.Y(n_10248)
);

HB1xp67_ASAP7_75t_L g10249 ( 
.A(n_9740),
.Y(n_10249)
);

CKINVDCx11_ASAP7_75t_R g10250 ( 
.A(n_9756),
.Y(n_10250)
);

INVx1_ASAP7_75t_L g10251 ( 
.A(n_9843),
.Y(n_10251)
);

AND2x4_ASAP7_75t_L g10252 ( 
.A(n_10073),
.B(n_4357),
.Y(n_10252)
);

AND2x4_ASAP7_75t_L g10253 ( 
.A(n_10105),
.B(n_9807),
.Y(n_10253)
);

BUFx2_ASAP7_75t_L g10254 ( 
.A(n_9857),
.Y(n_10254)
);

AOI22xp5_ASAP7_75t_L g10255 ( 
.A1(n_9693),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_10255)
);

NAND2xp5_ASAP7_75t_L g10256 ( 
.A(n_9758),
.B(n_19),
.Y(n_10256)
);

INVx2_ASAP7_75t_L g10257 ( 
.A(n_9850),
.Y(n_10257)
);

INVxp67_ASAP7_75t_SL g10258 ( 
.A(n_9846),
.Y(n_10258)
);

NAND2x1p5_ASAP7_75t_L g10259 ( 
.A(n_9697),
.B(n_4358),
.Y(n_10259)
);

INVx1_ASAP7_75t_L g10260 ( 
.A(n_9864),
.Y(n_10260)
);

NAND2x1p5_ASAP7_75t_L g10261 ( 
.A(n_9784),
.B(n_4359),
.Y(n_10261)
);

NAND2x1p5_ASAP7_75t_L g10262 ( 
.A(n_9839),
.B(n_4361),
.Y(n_10262)
);

AND2x4_ASAP7_75t_L g10263 ( 
.A(n_9733),
.B(n_4362),
.Y(n_10263)
);

INVx1_ASAP7_75t_L g10264 ( 
.A(n_9876),
.Y(n_10264)
);

AO22x2_ASAP7_75t_L g10265 ( 
.A1(n_10000),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_10265)
);

OR2x6_ASAP7_75t_L g10266 ( 
.A(n_9730),
.B(n_4363),
.Y(n_10266)
);

BUFx6f_ASAP7_75t_L g10267 ( 
.A(n_9730),
.Y(n_10267)
);

INVx1_ASAP7_75t_L g10268 ( 
.A(n_9898),
.Y(n_10268)
);

INVx1_ASAP7_75t_L g10269 ( 
.A(n_9901),
.Y(n_10269)
);

INVx1_ASAP7_75t_L g10270 ( 
.A(n_9925),
.Y(n_10270)
);

NAND2xp5_ASAP7_75t_L g10271 ( 
.A(n_10183),
.B(n_22),
.Y(n_10271)
);

AND2x4_ASAP7_75t_L g10272 ( 
.A(n_10157),
.B(n_4364),
.Y(n_10272)
);

INVx1_ASAP7_75t_L g10273 ( 
.A(n_9929),
.Y(n_10273)
);

NOR2xp33_ASAP7_75t_L g10274 ( 
.A(n_9703),
.B(n_4365),
.Y(n_10274)
);

NAND2x1p5_ASAP7_75t_L g10275 ( 
.A(n_9821),
.B(n_4366),
.Y(n_10275)
);

OAI221xp5_ASAP7_75t_L g10276 ( 
.A1(n_9738),
.A2(n_9985),
.B1(n_9999),
.B2(n_9814),
.C(n_9777),
.Y(n_10276)
);

NAND2xp5_ASAP7_75t_L g10277 ( 
.A(n_10187),
.B(n_23),
.Y(n_10277)
);

INVx2_ASAP7_75t_L g10278 ( 
.A(n_9940),
.Y(n_10278)
);

NAND2xp5_ASAP7_75t_L g10279 ( 
.A(n_9690),
.B(n_23),
.Y(n_10279)
);

INVxp67_ASAP7_75t_L g10280 ( 
.A(n_9710),
.Y(n_10280)
);

AND2x2_ASAP7_75t_L g10281 ( 
.A(n_10185),
.B(n_24),
.Y(n_10281)
);

AO22x2_ASAP7_75t_L g10282 ( 
.A1(n_9725),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_10282)
);

INVx5_ASAP7_75t_L g10283 ( 
.A(n_10043),
.Y(n_10283)
);

AO22x2_ASAP7_75t_L g10284 ( 
.A1(n_9754),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_10284)
);

BUFx3_ASAP7_75t_L g10285 ( 
.A(n_10025),
.Y(n_10285)
);

NAND2x1_ASAP7_75t_L g10286 ( 
.A(n_9979),
.B(n_4367),
.Y(n_10286)
);

INVx2_ASAP7_75t_L g10287 ( 
.A(n_9944),
.Y(n_10287)
);

OAI221xp5_ASAP7_75t_L g10288 ( 
.A1(n_9765),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.C(n_32),
.Y(n_10288)
);

INVx1_ASAP7_75t_L g10289 ( 
.A(n_9947),
.Y(n_10289)
);

NAND2xp5_ASAP7_75t_L g10290 ( 
.A(n_9695),
.B(n_29),
.Y(n_10290)
);

INVx1_ASAP7_75t_L g10291 ( 
.A(n_9688),
.Y(n_10291)
);

AO22x2_ASAP7_75t_L g10292 ( 
.A1(n_9735),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_10292)
);

INVx2_ASAP7_75t_L g10293 ( 
.A(n_9714),
.Y(n_10293)
);

INVx1_ASAP7_75t_L g10294 ( 
.A(n_9692),
.Y(n_10294)
);

INVx1_ASAP7_75t_L g10295 ( 
.A(n_9700),
.Y(n_10295)
);

BUFx6f_ASAP7_75t_SL g10296 ( 
.A(n_10177),
.Y(n_10296)
);

OR2x2_ASAP7_75t_L g10297 ( 
.A(n_10204),
.B(n_33),
.Y(n_10297)
);

AOI22xp33_ASAP7_75t_L g10298 ( 
.A1(n_9855),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_10298)
);

INVx1_ASAP7_75t_L g10299 ( 
.A(n_9704),
.Y(n_10299)
);

NAND2xp5_ASAP7_75t_L g10300 ( 
.A(n_10202),
.B(n_34),
.Y(n_10300)
);

AO22x2_ASAP7_75t_L g10301 ( 
.A1(n_9751),
.A2(n_10199),
.B1(n_10196),
.B2(n_10124),
.Y(n_10301)
);

AOI22xp33_ASAP7_75t_SL g10302 ( 
.A1(n_10011),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_10302)
);

NAND2x1p5_ASAP7_75t_L g10303 ( 
.A(n_9995),
.B(n_4368),
.Y(n_10303)
);

AO22x2_ASAP7_75t_L g10304 ( 
.A1(n_9897),
.A2(n_39),
.B1(n_36),
.B2(n_37),
.Y(n_10304)
);

INVx1_ASAP7_75t_L g10305 ( 
.A(n_9705),
.Y(n_10305)
);

INVx1_ASAP7_75t_L g10306 ( 
.A(n_9708),
.Y(n_10306)
);

AND2x2_ASAP7_75t_L g10307 ( 
.A(n_10186),
.B(n_39),
.Y(n_10307)
);

NAND2xp33_ASAP7_75t_L g10308 ( 
.A(n_9860),
.B(n_40),
.Y(n_10308)
);

AND2x2_ASAP7_75t_L g10309 ( 
.A(n_9921),
.B(n_41),
.Y(n_10309)
);

AND2x2_ASAP7_75t_L g10310 ( 
.A(n_9715),
.B(n_41),
.Y(n_10310)
);

INVx1_ASAP7_75t_L g10311 ( 
.A(n_9726),
.Y(n_10311)
);

AND2x4_ASAP7_75t_L g10312 ( 
.A(n_10163),
.B(n_4369),
.Y(n_10312)
);

INVx2_ASAP7_75t_L g10313 ( 
.A(n_9736),
.Y(n_10313)
);

AOI22xp5_ASAP7_75t_L g10314 ( 
.A1(n_9770),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_10314)
);

INVxp67_ASAP7_75t_L g10315 ( 
.A(n_9977),
.Y(n_10315)
);

INVx1_ASAP7_75t_L g10316 ( 
.A(n_9732),
.Y(n_10316)
);

AOI22xp5_ASAP7_75t_L g10317 ( 
.A1(n_9900),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_10317)
);

BUFx6f_ASAP7_75t_L g10318 ( 
.A(n_9865),
.Y(n_10318)
);

AO22x2_ASAP7_75t_L g10319 ( 
.A1(n_9717),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_10319)
);

AO22x2_ASAP7_75t_L g10320 ( 
.A1(n_9706),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_10320)
);

AOI22xp5_ASAP7_75t_L g10321 ( 
.A1(n_9913),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_10321)
);

OAI221xp5_ASAP7_75t_L g10322 ( 
.A1(n_10141),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.C(n_51),
.Y(n_10322)
);

A2O1A1Ixp33_ASAP7_75t_L g10323 ( 
.A1(n_9724),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_10323)
);

NAND2xp5_ASAP7_75t_L g10324 ( 
.A(n_9728),
.B(n_9741),
.Y(n_10324)
);

INVx1_ASAP7_75t_L g10325 ( 
.A(n_9745),
.Y(n_10325)
);

INVx1_ASAP7_75t_L g10326 ( 
.A(n_9761),
.Y(n_10326)
);

AOI22xp33_ASAP7_75t_L g10327 ( 
.A1(n_9737),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_10327)
);

AND2x4_ASAP7_75t_L g10328 ( 
.A(n_10171),
.B(n_4370),
.Y(n_10328)
);

INVx1_ASAP7_75t_L g10329 ( 
.A(n_9763),
.Y(n_10329)
);

AO22x2_ASAP7_75t_L g10330 ( 
.A1(n_9720),
.A2(n_58),
.B1(n_55),
.B2(n_56),
.Y(n_10330)
);

AOI22xp5_ASAP7_75t_L g10331 ( 
.A1(n_9923),
.A2(n_59),
.B1(n_55),
.B2(n_56),
.Y(n_10331)
);

INVx1_ASAP7_75t_L g10332 ( 
.A(n_9764),
.Y(n_10332)
);

INVx1_ASAP7_75t_L g10333 ( 
.A(n_9767),
.Y(n_10333)
);

INVx1_ASAP7_75t_L g10334 ( 
.A(n_9771),
.Y(n_10334)
);

INVx1_ASAP7_75t_L g10335 ( 
.A(n_9772),
.Y(n_10335)
);

INVx1_ASAP7_75t_L g10336 ( 
.A(n_9780),
.Y(n_10336)
);

NOR2xp33_ASAP7_75t_L g10337 ( 
.A(n_9753),
.B(n_4371),
.Y(n_10337)
);

AO22x2_ASAP7_75t_L g10338 ( 
.A1(n_9892),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_10338)
);

HB1xp67_ASAP7_75t_L g10339 ( 
.A(n_9750),
.Y(n_10339)
);

INVx1_ASAP7_75t_L g10340 ( 
.A(n_9795),
.Y(n_10340)
);

INVxp67_ASAP7_75t_SL g10341 ( 
.A(n_9775),
.Y(n_10341)
);

BUFx8_ASAP7_75t_L g10342 ( 
.A(n_10085),
.Y(n_10342)
);

NOR2xp33_ASAP7_75t_L g10343 ( 
.A(n_9752),
.B(n_4372),
.Y(n_10343)
);

INVx1_ASAP7_75t_L g10344 ( 
.A(n_9796),
.Y(n_10344)
);

INVx1_ASAP7_75t_L g10345 ( 
.A(n_9815),
.Y(n_10345)
);

NAND2xp5_ASAP7_75t_SL g10346 ( 
.A(n_9718),
.B(n_60),
.Y(n_10346)
);

NAND2xp5_ASAP7_75t_L g10347 ( 
.A(n_10192),
.B(n_10195),
.Y(n_10347)
);

INVx2_ASAP7_75t_L g10348 ( 
.A(n_9739),
.Y(n_10348)
);

INVx2_ASAP7_75t_L g10349 ( 
.A(n_9759),
.Y(n_10349)
);

NOR2xp33_ASAP7_75t_R g10350 ( 
.A(n_9746),
.B(n_9842),
.Y(n_10350)
);

OAI221xp5_ASAP7_75t_L g10351 ( 
.A1(n_9994),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.C(n_64),
.Y(n_10351)
);

INVx1_ASAP7_75t_L g10352 ( 
.A(n_9816),
.Y(n_10352)
);

INVx2_ASAP7_75t_SL g10353 ( 
.A(n_10043),
.Y(n_10353)
);

INVx1_ASAP7_75t_L g10354 ( 
.A(n_9845),
.Y(n_10354)
);

INVx2_ASAP7_75t_L g10355 ( 
.A(n_10184),
.Y(n_10355)
);

BUFx3_ASAP7_75t_L g10356 ( 
.A(n_10133),
.Y(n_10356)
);

INVxp67_ASAP7_75t_SL g10357 ( 
.A(n_9788),
.Y(n_10357)
);

AO22x2_ASAP7_75t_L g10358 ( 
.A1(n_9773),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_10358)
);

INVxp67_ASAP7_75t_L g10359 ( 
.A(n_9885),
.Y(n_10359)
);

INVx2_ASAP7_75t_SL g10360 ( 
.A(n_10133),
.Y(n_10360)
);

INVx2_ASAP7_75t_SL g10361 ( 
.A(n_10156),
.Y(n_10361)
);

AO22x2_ASAP7_75t_L g10362 ( 
.A1(n_9983),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_10362)
);

INVx1_ASAP7_75t_L g10363 ( 
.A(n_9861),
.Y(n_10363)
);

INVx1_ASAP7_75t_L g10364 ( 
.A(n_9872),
.Y(n_10364)
);

OAI221xp5_ASAP7_75t_L g10365 ( 
.A1(n_9958),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.C(n_69),
.Y(n_10365)
);

A2O1A1Ixp33_ASAP7_75t_L g10366 ( 
.A1(n_9716),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_10366)
);

INVx1_ASAP7_75t_L g10367 ( 
.A(n_9887),
.Y(n_10367)
);

INVx1_ASAP7_75t_L g10368 ( 
.A(n_9893),
.Y(n_10368)
);

NAND2xp5_ASAP7_75t_L g10369 ( 
.A(n_9927),
.B(n_70),
.Y(n_10369)
);

INVx1_ASAP7_75t_L g10370 ( 
.A(n_9904),
.Y(n_10370)
);

INVx1_ASAP7_75t_L g10371 ( 
.A(n_9905),
.Y(n_10371)
);

INVx1_ASAP7_75t_L g10372 ( 
.A(n_9910),
.Y(n_10372)
);

INVx1_ASAP7_75t_L g10373 ( 
.A(n_9911),
.Y(n_10373)
);

NAND2x1p5_ASAP7_75t_L g10374 ( 
.A(n_10015),
.B(n_4373),
.Y(n_10374)
);

OAI221xp5_ASAP7_75t_L g10375 ( 
.A1(n_10139),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.C(n_74),
.Y(n_10375)
);

INVx1_ASAP7_75t_L g10376 ( 
.A(n_10189),
.Y(n_10376)
);

INVx1_ASAP7_75t_L g10377 ( 
.A(n_10190),
.Y(n_10377)
);

BUFx2_ASAP7_75t_L g10378 ( 
.A(n_9866),
.Y(n_10378)
);

NAND2x1p5_ASAP7_75t_L g10379 ( 
.A(n_10042),
.B(n_4374),
.Y(n_10379)
);

AND2x4_ASAP7_75t_L g10380 ( 
.A(n_9890),
.B(n_10110),
.Y(n_10380)
);

OAI22xp5_ASAP7_75t_L g10381 ( 
.A1(n_9959),
.A2(n_74),
.B1(n_71),
.B2(n_72),
.Y(n_10381)
);

BUFx8_ASAP7_75t_L g10382 ( 
.A(n_9721),
.Y(n_10382)
);

INVx1_ASAP7_75t_L g10383 ( 
.A(n_10191),
.Y(n_10383)
);

INVx1_ASAP7_75t_L g10384 ( 
.A(n_10197),
.Y(n_10384)
);

AND2x4_ASAP7_75t_L g10385 ( 
.A(n_9890),
.B(n_4375),
.Y(n_10385)
);

OAI22xp33_ASAP7_75t_SL g10386 ( 
.A1(n_10136),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_10386)
);

AO22x2_ASAP7_75t_L g10387 ( 
.A1(n_10203),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_10387)
);

INVx2_ASAP7_75t_L g10388 ( 
.A(n_10205),
.Y(n_10388)
);

NAND2xp5_ASAP7_75t_L g10389 ( 
.A(n_9988),
.B(n_79),
.Y(n_10389)
);

AND2x2_ASAP7_75t_L g10390 ( 
.A(n_10201),
.B(n_79),
.Y(n_10390)
);

INVx2_ASAP7_75t_L g10391 ( 
.A(n_9974),
.Y(n_10391)
);

NAND2xp5_ASAP7_75t_SL g10392 ( 
.A(n_10101),
.B(n_80),
.Y(n_10392)
);

AND2x4_ASAP7_75t_L g10393 ( 
.A(n_9903),
.B(n_4376),
.Y(n_10393)
);

AO22x2_ASAP7_75t_L g10394 ( 
.A1(n_9858),
.A2(n_9987),
.B1(n_9978),
.B2(n_9713),
.Y(n_10394)
);

AND2x2_ASAP7_75t_L g10395 ( 
.A(n_9936),
.B(n_80),
.Y(n_10395)
);

AOI22xp5_ASAP7_75t_L g10396 ( 
.A1(n_9856),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_10396)
);

NAND2x1p5_ASAP7_75t_L g10397 ( 
.A(n_9822),
.B(n_4377),
.Y(n_10397)
);

INVx1_ASAP7_75t_L g10398 ( 
.A(n_9955),
.Y(n_10398)
);

OAI22xp5_ASAP7_75t_SL g10399 ( 
.A1(n_10131),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_10399)
);

INVx1_ASAP7_75t_L g10400 ( 
.A(n_9969),
.Y(n_10400)
);

INVx1_ASAP7_75t_L g10401 ( 
.A(n_9933),
.Y(n_10401)
);

INVx1_ASAP7_75t_L g10402 ( 
.A(n_9956),
.Y(n_10402)
);

AO22x2_ASAP7_75t_L g10403 ( 
.A1(n_9742),
.A2(n_87),
.B1(n_84),
.B2(n_86),
.Y(n_10403)
);

INVx2_ASAP7_75t_L g10404 ( 
.A(n_9968),
.Y(n_10404)
);

OAI221xp5_ASAP7_75t_L g10405 ( 
.A1(n_10059),
.A2(n_87),
.B1(n_84),
.B2(n_86),
.C(n_88),
.Y(n_10405)
);

OAI221xp5_ASAP7_75t_L g10406 ( 
.A1(n_10034),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.C(n_92),
.Y(n_10406)
);

INVx1_ASAP7_75t_L g10407 ( 
.A(n_10017),
.Y(n_10407)
);

AO22x2_ASAP7_75t_L g10408 ( 
.A1(n_10188),
.A2(n_92),
.B1(n_89),
.B2(n_90),
.Y(n_10408)
);

OAI221xp5_ASAP7_75t_L g10409 ( 
.A1(n_10067),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.C(n_96),
.Y(n_10409)
);

INVx1_ASAP7_75t_L g10410 ( 
.A(n_10050),
.Y(n_10410)
);

INVxp67_ASAP7_75t_L g10411 ( 
.A(n_10037),
.Y(n_10411)
);

BUFx2_ASAP7_75t_L g10412 ( 
.A(n_9930),
.Y(n_10412)
);

INVx1_ASAP7_75t_L g10413 ( 
.A(n_10052),
.Y(n_10413)
);

INVx1_ASAP7_75t_L g10414 ( 
.A(n_10055),
.Y(n_10414)
);

NAND2xp5_ASAP7_75t_SL g10415 ( 
.A(n_9755),
.B(n_93),
.Y(n_10415)
);

AND2x4_ASAP7_75t_L g10416 ( 
.A(n_9914),
.B(n_4379),
.Y(n_10416)
);

AO22x2_ASAP7_75t_L g10417 ( 
.A1(n_9760),
.A2(n_97),
.B1(n_94),
.B2(n_95),
.Y(n_10417)
);

AOI22xp5_ASAP7_75t_L g10418 ( 
.A1(n_10102),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_10418)
);

AOI22xp5_ASAP7_75t_SL g10419 ( 
.A1(n_9799),
.A2(n_101),
.B1(n_98),
.B2(n_99),
.Y(n_10419)
);

AO22x2_ASAP7_75t_L g10420 ( 
.A1(n_10068),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_10420)
);

INVx1_ASAP7_75t_L g10421 ( 
.A(n_10058),
.Y(n_10421)
);

NAND2x1p5_ASAP7_75t_L g10422 ( 
.A(n_9877),
.B(n_4380),
.Y(n_10422)
);

NAND2xp5_ASAP7_75t_L g10423 ( 
.A(n_9805),
.B(n_102),
.Y(n_10423)
);

INVx2_ASAP7_75t_L g10424 ( 
.A(n_9973),
.Y(n_10424)
);

INVx2_ASAP7_75t_L g10425 ( 
.A(n_9997),
.Y(n_10425)
);

HB1xp67_ASAP7_75t_L g10426 ( 
.A(n_9827),
.Y(n_10426)
);

AOI22xp5_ASAP7_75t_L g10427 ( 
.A1(n_9712),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_10427)
);

INVx1_ASAP7_75t_L g10428 ( 
.A(n_10063),
.Y(n_10428)
);

OR2x6_ASAP7_75t_L g10429 ( 
.A(n_10156),
.B(n_4382),
.Y(n_10429)
);

INVx1_ASAP7_75t_L g10430 ( 
.A(n_10019),
.Y(n_10430)
);

NAND2xp5_ASAP7_75t_SL g10431 ( 
.A(n_9727),
.B(n_104),
.Y(n_10431)
);

OR2x2_ASAP7_75t_L g10432 ( 
.A(n_9852),
.B(n_105),
.Y(n_10432)
);

INVx1_ASAP7_75t_L g10433 ( 
.A(n_10023),
.Y(n_10433)
);

AND2x2_ASAP7_75t_L g10434 ( 
.A(n_9937),
.B(n_106),
.Y(n_10434)
);

INVx1_ASAP7_75t_L g10435 ( 
.A(n_10047),
.Y(n_10435)
);

NAND2x1p5_ASAP7_75t_L g10436 ( 
.A(n_9884),
.B(n_4384),
.Y(n_10436)
);

CKINVDCx5p33_ASAP7_75t_R g10437 ( 
.A(n_9982),
.Y(n_10437)
);

INVx1_ASAP7_75t_L g10438 ( 
.A(n_10001),
.Y(n_10438)
);

OR2x6_ASAP7_75t_L g10439 ( 
.A(n_10117),
.B(n_4385),
.Y(n_10439)
);

INVx2_ASAP7_75t_L g10440 ( 
.A(n_10005),
.Y(n_10440)
);

NOR2xp33_ASAP7_75t_L g10441 ( 
.A(n_9854),
.B(n_4387),
.Y(n_10441)
);

INVx1_ASAP7_75t_L g10442 ( 
.A(n_10007),
.Y(n_10442)
);

AO22x2_ASAP7_75t_L g10443 ( 
.A1(n_9869),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_10443)
);

INVx2_ASAP7_75t_L g10444 ( 
.A(n_10010),
.Y(n_10444)
);

OAI22xp5_ASAP7_75t_L g10445 ( 
.A1(n_9932),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_10445)
);

INVx3_ASAP7_75t_L g10446 ( 
.A(n_10004),
.Y(n_10446)
);

AO22x2_ASAP7_75t_L g10447 ( 
.A1(n_9991),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_10447)
);

OAI22xp5_ASAP7_75t_L g10448 ( 
.A1(n_9820),
.A2(n_114),
.B1(n_110),
.B2(n_113),
.Y(n_10448)
);

AO22x2_ASAP7_75t_L g10449 ( 
.A1(n_10181),
.A2(n_116),
.B1(n_113),
.B2(n_115),
.Y(n_10449)
);

INVx1_ASAP7_75t_SL g10450 ( 
.A(n_10175),
.Y(n_10450)
);

NOR2xp33_ASAP7_75t_L g10451 ( 
.A(n_9757),
.B(n_4389),
.Y(n_10451)
);

INVxp67_ASAP7_75t_L g10452 ( 
.A(n_10127),
.Y(n_10452)
);

INVx1_ASAP7_75t_L g10453 ( 
.A(n_10018),
.Y(n_10453)
);

INVx1_ASAP7_75t_L g10454 ( 
.A(n_10020),
.Y(n_10454)
);

INVx1_ASAP7_75t_L g10455 ( 
.A(n_10044),
.Y(n_10455)
);

INVx1_ASAP7_75t_L g10456 ( 
.A(n_10054),
.Y(n_10456)
);

NAND2xp5_ASAP7_75t_L g10457 ( 
.A(n_9778),
.B(n_9779),
.Y(n_10457)
);

INVx1_ASAP7_75t_L g10458 ( 
.A(n_10057),
.Y(n_10458)
);

AO22x2_ASAP7_75t_L g10459 ( 
.A1(n_9954),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_10459)
);

BUFx2_ASAP7_75t_L g10460 ( 
.A(n_10029),
.Y(n_10460)
);

CKINVDCx5p33_ASAP7_75t_R g10461 ( 
.A(n_9709),
.Y(n_10461)
);

INVx1_ASAP7_75t_L g10462 ( 
.A(n_10064),
.Y(n_10462)
);

INVxp67_ASAP7_75t_L g10463 ( 
.A(n_9838),
.Y(n_10463)
);

AOI22xp5_ASAP7_75t_L g10464 ( 
.A1(n_10003),
.A2(n_9882),
.B1(n_9879),
.B2(n_9791),
.Y(n_10464)
);

INVxp67_ASAP7_75t_L g10465 ( 
.A(n_9853),
.Y(n_10465)
);

INVx2_ASAP7_75t_L g10466 ( 
.A(n_9731),
.Y(n_10466)
);

INVx1_ASAP7_75t_L g10467 ( 
.A(n_10027),
.Y(n_10467)
);

INVx1_ASAP7_75t_L g10468 ( 
.A(n_10031),
.Y(n_10468)
);

INVx2_ASAP7_75t_L g10469 ( 
.A(n_9731),
.Y(n_10469)
);

NAND2xp5_ASAP7_75t_L g10470 ( 
.A(n_9797),
.B(n_117),
.Y(n_10470)
);

HB1xp67_ASAP7_75t_L g10471 ( 
.A(n_10036),
.Y(n_10471)
);

INVx1_ASAP7_75t_L g10472 ( 
.A(n_10039),
.Y(n_10472)
);

INVx4_ASAP7_75t_L g10473 ( 
.A(n_9865),
.Y(n_10473)
);

OAI221xp5_ASAP7_75t_L g10474 ( 
.A1(n_9902),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.C(n_121),
.Y(n_10474)
);

AO22x2_ASAP7_75t_L g10475 ( 
.A1(n_9744),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_10475)
);

INVx1_ASAP7_75t_L g10476 ( 
.A(n_10040),
.Y(n_10476)
);

NAND2xp5_ASAP7_75t_SL g10477 ( 
.A(n_9731),
.B(n_122),
.Y(n_10477)
);

AO22x2_ASAP7_75t_L g10478 ( 
.A1(n_9748),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_10478)
);

AO22x2_ASAP7_75t_L g10479 ( 
.A1(n_9957),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_10479)
);

NAND2x1p5_ASAP7_75t_L g10480 ( 
.A(n_9699),
.B(n_4390),
.Y(n_10480)
);

INVx1_ASAP7_75t_L g10481 ( 
.A(n_10045),
.Y(n_10481)
);

OR2x2_ASAP7_75t_L g10482 ( 
.A(n_9800),
.B(n_126),
.Y(n_10482)
);

INVx1_ASAP7_75t_L g10483 ( 
.A(n_10048),
.Y(n_10483)
);

INVx1_ASAP7_75t_L g10484 ( 
.A(n_10053),
.Y(n_10484)
);

INVx1_ASAP7_75t_L g10485 ( 
.A(n_10061),
.Y(n_10485)
);

CKINVDCx16_ASAP7_75t_R g10486 ( 
.A(n_9781),
.Y(n_10486)
);

BUFx8_ASAP7_75t_L g10487 ( 
.A(n_9975),
.Y(n_10487)
);

AOI22xp5_ASAP7_75t_L g10488 ( 
.A1(n_9825),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_10488)
);

NAND2x1p5_ASAP7_75t_L g10489 ( 
.A(n_10200),
.B(n_4392),
.Y(n_10489)
);

NAND2x1p5_ASAP7_75t_L g10490 ( 
.A(n_10035),
.B(n_4393),
.Y(n_10490)
);

AO22x2_ASAP7_75t_L g10491 ( 
.A1(n_10115),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_10491)
);

INVx1_ASAP7_75t_L g10492 ( 
.A(n_10065),
.Y(n_10492)
);

INVxp67_ASAP7_75t_L g10493 ( 
.A(n_10161),
.Y(n_10493)
);

AO22x2_ASAP7_75t_L g10494 ( 
.A1(n_9801),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_10494)
);

INVx1_ASAP7_75t_L g10495 ( 
.A(n_9918),
.Y(n_10495)
);

OA22x2_ASAP7_75t_L g10496 ( 
.A1(n_10089),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_10496)
);

OR2x2_ASAP7_75t_SL g10497 ( 
.A(n_9952),
.B(n_133),
.Y(n_10497)
);

AND2x2_ASAP7_75t_L g10498 ( 
.A(n_9826),
.B(n_134),
.Y(n_10498)
);

INVxp67_ASAP7_75t_L g10499 ( 
.A(n_10168),
.Y(n_10499)
);

INVx1_ASAP7_75t_L g10500 ( 
.A(n_9928),
.Y(n_10500)
);

NAND3xp33_ASAP7_75t_SL g10501 ( 
.A(n_9824),
.B(n_9844),
.C(n_9996),
.Y(n_10501)
);

NAND2xp5_ASAP7_75t_L g10502 ( 
.A(n_9804),
.B(n_134),
.Y(n_10502)
);

INVx1_ASAP7_75t_L g10503 ( 
.A(n_9931),
.Y(n_10503)
);

CKINVDCx5p33_ASAP7_75t_R g10504 ( 
.A(n_9963),
.Y(n_10504)
);

INVx1_ASAP7_75t_L g10505 ( 
.A(n_9938),
.Y(n_10505)
);

INVx1_ASAP7_75t_L g10506 ( 
.A(n_9943),
.Y(n_10506)
);

NAND2xp5_ASAP7_75t_L g10507 ( 
.A(n_9859),
.B(n_9992),
.Y(n_10507)
);

AO22x2_ASAP7_75t_L g10508 ( 
.A1(n_10137),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_10508)
);

NAND2xp5_ASAP7_75t_L g10509 ( 
.A(n_9998),
.B(n_135),
.Y(n_10509)
);

INVx1_ASAP7_75t_L g10510 ( 
.A(n_9946),
.Y(n_10510)
);

INVx1_ASAP7_75t_L g10511 ( 
.A(n_9948),
.Y(n_10511)
);

NAND2xp5_ASAP7_75t_L g10512 ( 
.A(n_10002),
.B(n_137),
.Y(n_10512)
);

INVx1_ASAP7_75t_L g10513 ( 
.A(n_9990),
.Y(n_10513)
);

INVx1_ASAP7_75t_L g10514 ( 
.A(n_9949),
.Y(n_10514)
);

OAI221xp5_ASAP7_75t_L g10515 ( 
.A1(n_10008),
.A2(n_10009),
.B1(n_10069),
.B2(n_10016),
.C(n_10140),
.Y(n_10515)
);

NAND2xp5_ASAP7_75t_L g10516 ( 
.A(n_10109),
.B(n_138),
.Y(n_10516)
);

INVx1_ASAP7_75t_L g10517 ( 
.A(n_9950),
.Y(n_10517)
);

OAI22xp5_ASAP7_75t_L g10518 ( 
.A1(n_9729),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_10518)
);

AO22x2_ASAP7_75t_L g10519 ( 
.A1(n_10150),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_10519)
);

INVx1_ASAP7_75t_L g10520 ( 
.A(n_9962),
.Y(n_10520)
);

INVx1_ASAP7_75t_L g10521 ( 
.A(n_9965),
.Y(n_10521)
);

AO22x2_ASAP7_75t_L g10522 ( 
.A1(n_10155),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_10522)
);

BUFx6f_ASAP7_75t_SL g10523 ( 
.A(n_9799),
.Y(n_10523)
);

OAI22xp5_ASAP7_75t_L g10524 ( 
.A1(n_9729),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_10524)
);

INVx1_ASAP7_75t_L g10525 ( 
.A(n_9967),
.Y(n_10525)
);

NAND2xp5_ASAP7_75t_L g10526 ( 
.A(n_10066),
.B(n_146),
.Y(n_10526)
);

NAND2xp5_ASAP7_75t_L g10527 ( 
.A(n_10082),
.B(n_146),
.Y(n_10527)
);

INVx2_ASAP7_75t_L g10528 ( 
.A(n_9731),
.Y(n_10528)
);

NAND2xp5_ASAP7_75t_L g10529 ( 
.A(n_10118),
.B(n_147),
.Y(n_10529)
);

OR2x2_ASAP7_75t_L g10530 ( 
.A(n_9971),
.B(n_147),
.Y(n_10530)
);

NAND2xp5_ASAP7_75t_SL g10531 ( 
.A(n_9837),
.B(n_9812),
.Y(n_10531)
);

INVx1_ASAP7_75t_L g10532 ( 
.A(n_9976),
.Y(n_10532)
);

INVx1_ASAP7_75t_L g10533 ( 
.A(n_9981),
.Y(n_10533)
);

NAND2xp5_ASAP7_75t_L g10534 ( 
.A(n_10114),
.B(n_148),
.Y(n_10534)
);

INVx1_ASAP7_75t_L g10535 ( 
.A(n_9984),
.Y(n_10535)
);

INVx1_ASAP7_75t_L g10536 ( 
.A(n_9989),
.Y(n_10536)
);

INVx2_ASAP7_75t_L g10537 ( 
.A(n_9837),
.Y(n_10537)
);

INVx1_ASAP7_75t_L g10538 ( 
.A(n_9808),
.Y(n_10538)
);

AO22x2_ASAP7_75t_L g10539 ( 
.A1(n_10160),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_10539)
);

BUFx8_ASAP7_75t_L g10540 ( 
.A(n_10035),
.Y(n_10540)
);

INVx1_ASAP7_75t_L g10541 ( 
.A(n_9818),
.Y(n_10541)
);

AO22x2_ASAP7_75t_L g10542 ( 
.A1(n_10162),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_10542)
);

INVx1_ASAP7_75t_L g10543 ( 
.A(n_9829),
.Y(n_10543)
);

INVx2_ASAP7_75t_SL g10544 ( 
.A(n_10098),
.Y(n_10544)
);

INVx2_ASAP7_75t_L g10545 ( 
.A(n_9837),
.Y(n_10545)
);

AO22x2_ASAP7_75t_L g10546 ( 
.A1(n_10180),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_10546)
);

AO22x2_ASAP7_75t_L g10547 ( 
.A1(n_10173),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_10547)
);

AO22x2_ASAP7_75t_L g10548 ( 
.A1(n_10178),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_10548)
);

NAND2x1p5_ASAP7_75t_L g10549 ( 
.A(n_10098),
.B(n_4394),
.Y(n_10549)
);

INVx1_ASAP7_75t_L g10550 ( 
.A(n_9841),
.Y(n_10550)
);

INVx1_ASAP7_75t_L g10551 ( 
.A(n_9868),
.Y(n_10551)
);

NAND2x1p5_ASAP7_75t_L g10552 ( 
.A(n_9723),
.B(n_4395),
.Y(n_10552)
);

AND2x2_ASAP7_75t_L g10553 ( 
.A(n_10014),
.B(n_157),
.Y(n_10553)
);

INVx1_ASAP7_75t_L g10554 ( 
.A(n_9871),
.Y(n_10554)
);

INVx1_ASAP7_75t_L g10555 ( 
.A(n_9878),
.Y(n_10555)
);

INVx1_ASAP7_75t_L g10556 ( 
.A(n_9883),
.Y(n_10556)
);

INVx1_ASAP7_75t_L g10557 ( 
.A(n_9886),
.Y(n_10557)
);

INVx1_ASAP7_75t_L g10558 ( 
.A(n_9889),
.Y(n_10558)
);

INVx1_ASAP7_75t_L g10559 ( 
.A(n_9891),
.Y(n_10559)
);

INVx1_ASAP7_75t_L g10560 ( 
.A(n_9894),
.Y(n_10560)
);

INVx1_ASAP7_75t_L g10561 ( 
.A(n_9895),
.Y(n_10561)
);

AO22x2_ASAP7_75t_L g10562 ( 
.A1(n_10116),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_10562)
);

AND2x2_ASAP7_75t_L g10563 ( 
.A(n_10170),
.B(n_158),
.Y(n_10563)
);

NAND2xp5_ASAP7_75t_L g10564 ( 
.A(n_10119),
.B(n_159),
.Y(n_10564)
);

NAND2x1p5_ASAP7_75t_L g10565 ( 
.A(n_10158),
.B(n_4396),
.Y(n_10565)
);

INVx1_ASAP7_75t_L g10566 ( 
.A(n_9899),
.Y(n_10566)
);

INVx1_ASAP7_75t_L g10567 ( 
.A(n_9906),
.Y(n_10567)
);

INVx2_ASAP7_75t_L g10568 ( 
.A(n_9837),
.Y(n_10568)
);

INVx1_ASAP7_75t_L g10569 ( 
.A(n_9912),
.Y(n_10569)
);

INVx1_ASAP7_75t_L g10570 ( 
.A(n_9916),
.Y(n_10570)
);

INVx2_ASAP7_75t_SL g10571 ( 
.A(n_9935),
.Y(n_10571)
);

AO22x2_ASAP7_75t_L g10572 ( 
.A1(n_10126),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_10572)
);

INVx1_ASAP7_75t_L g10573 ( 
.A(n_9917),
.Y(n_10573)
);

AOI22xp5_ASAP7_75t_L g10574 ( 
.A1(n_10142),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_10574)
);

INVx1_ASAP7_75t_L g10575 ( 
.A(n_10062),
.Y(n_10575)
);

INVx1_ASAP7_75t_L g10576 ( 
.A(n_10062),
.Y(n_10576)
);

INVx1_ASAP7_75t_L g10577 ( 
.A(n_9953),
.Y(n_10577)
);

AND2x2_ASAP7_75t_L g10578 ( 
.A(n_10084),
.B(n_163),
.Y(n_10578)
);

INVx1_ASAP7_75t_L g10579 ( 
.A(n_9953),
.Y(n_10579)
);

AO22x2_ASAP7_75t_L g10580 ( 
.A1(n_10087),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_10580)
);

INVx2_ASAP7_75t_L g10581 ( 
.A(n_9953),
.Y(n_10581)
);

AO22x2_ASAP7_75t_L g10582 ( 
.A1(n_10090),
.A2(n_167),
.B1(n_164),
.B2(n_166),
.Y(n_10582)
);

NAND2xp5_ASAP7_75t_L g10583 ( 
.A(n_10041),
.B(n_167),
.Y(n_10583)
);

INVx2_ASAP7_75t_SL g10584 ( 
.A(n_10038),
.Y(n_10584)
);

INVx1_ASAP7_75t_L g10585 ( 
.A(n_9953),
.Y(n_10585)
);

NAND2xp5_ASAP7_75t_SL g10586 ( 
.A(n_10129),
.B(n_168),
.Y(n_10586)
);

INVx1_ASAP7_75t_L g10587 ( 
.A(n_9734),
.Y(n_10587)
);

INVx1_ASAP7_75t_L g10588 ( 
.A(n_10122),
.Y(n_10588)
);

OR2x2_ASAP7_75t_L g10589 ( 
.A(n_10138),
.B(n_168),
.Y(n_10589)
);

AO22x2_ASAP7_75t_L g10590 ( 
.A1(n_10095),
.A2(n_10099),
.B1(n_10164),
.B2(n_10159),
.Y(n_10590)
);

AO22x2_ASAP7_75t_L g10591 ( 
.A1(n_9794),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_10591)
);

NAND2xp5_ASAP7_75t_L g10592 ( 
.A(n_10056),
.B(n_169),
.Y(n_10592)
);

INVxp67_ASAP7_75t_L g10593 ( 
.A(n_10169),
.Y(n_10593)
);

INVx1_ASAP7_75t_L g10594 ( 
.A(n_10182),
.Y(n_10594)
);

NAND2x1p5_ASAP7_75t_L g10595 ( 
.A(n_10113),
.B(n_4397),
.Y(n_10595)
);

INVx1_ASAP7_75t_L g10596 ( 
.A(n_10046),
.Y(n_10596)
);

INVx2_ASAP7_75t_L g10597 ( 
.A(n_10145),
.Y(n_10597)
);

INVx1_ASAP7_75t_L g10598 ( 
.A(n_9811),
.Y(n_10598)
);

AO22x2_ASAP7_75t_L g10599 ( 
.A1(n_9803),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_10599)
);

INVx1_ASAP7_75t_L g10600 ( 
.A(n_9811),
.Y(n_10600)
);

AO22x2_ASAP7_75t_L g10601 ( 
.A1(n_9833),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_10601)
);

INVx1_ASAP7_75t_L g10602 ( 
.A(n_9811),
.Y(n_10602)
);

INVxp67_ASAP7_75t_L g10603 ( 
.A(n_10134),
.Y(n_10603)
);

INVxp67_ASAP7_75t_L g10604 ( 
.A(n_10135),
.Y(n_10604)
);

AO22x2_ASAP7_75t_L g10605 ( 
.A1(n_9980),
.A2(n_176),
.B1(n_173),
.B2(n_174),
.Y(n_10605)
);

INVx2_ASAP7_75t_SL g10606 ( 
.A(n_10051),
.Y(n_10606)
);

NOR2xp33_ASAP7_75t_L g10607 ( 
.A(n_9926),
.B(n_4400),
.Y(n_10607)
);

NAND2xp5_ASAP7_75t_SL g10608 ( 
.A(n_9888),
.B(n_176),
.Y(n_10608)
);

AO22x2_ASAP7_75t_L g10609 ( 
.A1(n_9920),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_10609)
);

AOI22xp5_ASAP7_75t_L g10610 ( 
.A1(n_10147),
.A2(n_180),
.B1(n_177),
.B2(n_178),
.Y(n_10610)
);

OAI22xp5_ASAP7_75t_L g10611 ( 
.A1(n_9867),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_10611)
);

INVx1_ASAP7_75t_L g10612 ( 
.A(n_10079),
.Y(n_10612)
);

AO22x2_ASAP7_75t_L g10613 ( 
.A1(n_10074),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_10613)
);

AO22x2_ASAP7_75t_L g10614 ( 
.A1(n_10078),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_10614)
);

INVx1_ASAP7_75t_L g10615 ( 
.A(n_10072),
.Y(n_10615)
);

INVx1_ASAP7_75t_L g10616 ( 
.A(n_10152),
.Y(n_10616)
);

AO22x2_ASAP7_75t_L g10617 ( 
.A1(n_10081),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_10617)
);

OR2x2_ASAP7_75t_L g10618 ( 
.A(n_10103),
.B(n_186),
.Y(n_10618)
);

INVx1_ASAP7_75t_L g10619 ( 
.A(n_10153),
.Y(n_10619)
);

NAND2xp5_ASAP7_75t_SL g10620 ( 
.A(n_9787),
.B(n_187),
.Y(n_10620)
);

OAI221xp5_ASAP7_75t_L g10621 ( 
.A1(n_9875),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_191),
.Y(n_10621)
);

NAND2x1p5_ASAP7_75t_L g10622 ( 
.A(n_9722),
.B(n_4401),
.Y(n_10622)
);

INVx2_ASAP7_75t_L g10623 ( 
.A(n_10076),
.Y(n_10623)
);

INVx2_ASAP7_75t_L g10624 ( 
.A(n_9828),
.Y(n_10624)
);

INVx2_ASAP7_75t_L g10625 ( 
.A(n_9707),
.Y(n_10625)
);

INVx1_ASAP7_75t_L g10626 ( 
.A(n_10104),
.Y(n_10626)
);

AO22x2_ASAP7_75t_L g10627 ( 
.A1(n_10093),
.A2(n_192),
.B1(n_188),
.B2(n_190),
.Y(n_10627)
);

INVxp67_ASAP7_75t_SL g10628 ( 
.A(n_9743),
.Y(n_10628)
);

INVx2_ASAP7_75t_L g10629 ( 
.A(n_10086),
.Y(n_10629)
);

NAND2xp5_ASAP7_75t_L g10630 ( 
.A(n_9809),
.B(n_192),
.Y(n_10630)
);

NAND2xp5_ASAP7_75t_SL g10631 ( 
.A(n_10075),
.B(n_193),
.Y(n_10631)
);

AND2x2_ASAP7_75t_L g10632 ( 
.A(n_10112),
.B(n_193),
.Y(n_10632)
);

INVx1_ASAP7_75t_L g10633 ( 
.A(n_9961),
.Y(n_10633)
);

CKINVDCx5p33_ASAP7_75t_R g10634 ( 
.A(n_9702),
.Y(n_10634)
);

AND2x4_ASAP7_75t_L g10635 ( 
.A(n_10117),
.B(n_4402),
.Y(n_10635)
);

BUFx3_ASAP7_75t_L g10636 ( 
.A(n_10120),
.Y(n_10636)
);

INVx1_ASAP7_75t_L g10637 ( 
.A(n_9964),
.Y(n_10637)
);

INVx1_ASAP7_75t_L g10638 ( 
.A(n_10077),
.Y(n_10638)
);

AO22x2_ASAP7_75t_L g10639 ( 
.A1(n_10097),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_10639)
);

AOI22xp5_ASAP7_75t_L g10640 ( 
.A1(n_9922),
.A2(n_197),
.B1(n_194),
.B2(n_196),
.Y(n_10640)
);

NAND2xp5_ASAP7_75t_L g10641 ( 
.A(n_9799),
.B(n_197),
.Y(n_10641)
);

OR2x2_ASAP7_75t_SL g10642 ( 
.A(n_10128),
.B(n_198),
.Y(n_10642)
);

NAND2xp5_ASAP7_75t_L g10643 ( 
.A(n_10012),
.B(n_198),
.Y(n_10643)
);

NOR2xp33_ASAP7_75t_L g10644 ( 
.A(n_9786),
.B(n_4403),
.Y(n_10644)
);

HB1xp67_ASAP7_75t_L g10645 ( 
.A(n_10106),
.Y(n_10645)
);

NAND2xp5_ASAP7_75t_L g10646 ( 
.A(n_10083),
.B(n_199),
.Y(n_10646)
);

NAND2xp5_ASAP7_75t_L g10647 ( 
.A(n_10144),
.B(n_200),
.Y(n_10647)
);

OAI221xp5_ASAP7_75t_L g10648 ( 
.A1(n_9896),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.C(n_204),
.Y(n_10648)
);

INVx2_ASAP7_75t_SL g10649 ( 
.A(n_9941),
.Y(n_10649)
);

NAND2xp5_ASAP7_75t_L g10650 ( 
.A(n_9874),
.B(n_202),
.Y(n_10650)
);

AO22x2_ASAP7_75t_L g10651 ( 
.A1(n_10100),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_10651)
);

AND2x4_ASAP7_75t_L g10652 ( 
.A(n_9774),
.B(n_4404),
.Y(n_10652)
);

INVx1_ASAP7_75t_L g10653 ( 
.A(n_9960),
.Y(n_10653)
);

AO22x2_ASAP7_75t_L g10654 ( 
.A1(n_10111),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_10654)
);

INVx1_ASAP7_75t_L g10655 ( 
.A(n_10088),
.Y(n_10655)
);

NAND2xp33_ASAP7_75t_L g10656 ( 
.A(n_9870),
.B(n_9934),
.Y(n_10656)
);

AO22x2_ASAP7_75t_L g10657 ( 
.A1(n_10121),
.A2(n_10125),
.B1(n_10130),
.B2(n_10123),
.Y(n_10657)
);

INVx1_ASAP7_75t_L g10658 ( 
.A(n_10151),
.Y(n_10658)
);

INVxp67_ASAP7_75t_L g10659 ( 
.A(n_10172),
.Y(n_10659)
);

INVx2_ASAP7_75t_L g10660 ( 
.A(n_9774),
.Y(n_10660)
);

INVx1_ASAP7_75t_L g10661 ( 
.A(n_9939),
.Y(n_10661)
);

INVx1_ASAP7_75t_L g10662 ( 
.A(n_10174),
.Y(n_10662)
);

INVx2_ASAP7_75t_SL g10663 ( 
.A(n_9986),
.Y(n_10663)
);

INVxp67_ASAP7_75t_L g10664 ( 
.A(n_10165),
.Y(n_10664)
);

INVx1_ASAP7_75t_L g10665 ( 
.A(n_9909),
.Y(n_10665)
);

OAI221xp5_ASAP7_75t_L g10666 ( 
.A1(n_10193),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.C(n_209),
.Y(n_10666)
);

INVx1_ASAP7_75t_L g10667 ( 
.A(n_10096),
.Y(n_10667)
);

INVx2_ASAP7_75t_L g10668 ( 
.A(n_10013),
.Y(n_10668)
);

BUFx3_ASAP7_75t_L g10669 ( 
.A(n_10080),
.Y(n_10669)
);

INVx2_ASAP7_75t_L g10670 ( 
.A(n_10132),
.Y(n_10670)
);

NAND2xp5_ASAP7_75t_L g10671 ( 
.A(n_10026),
.B(n_208),
.Y(n_10671)
);

NAND2xp5_ASAP7_75t_L g10672 ( 
.A(n_9993),
.B(n_209),
.Y(n_10672)
);

NOR2xp33_ASAP7_75t_L g10673 ( 
.A(n_9834),
.B(n_4405),
.Y(n_10673)
);

BUFx8_ASAP7_75t_L g10674 ( 
.A(n_10108),
.Y(n_10674)
);

INVx2_ASAP7_75t_L g10675 ( 
.A(n_9848),
.Y(n_10675)
);

INVx1_ASAP7_75t_SL g10676 ( 
.A(n_9863),
.Y(n_10676)
);

NAND2xp5_ASAP7_75t_L g10677 ( 
.A(n_10030),
.B(n_211),
.Y(n_10677)
);

AO22x2_ASAP7_75t_L g10678 ( 
.A1(n_10032),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_10678)
);

INVx1_ASAP7_75t_L g10679 ( 
.A(n_10006),
.Y(n_10679)
);

INVx3_ASAP7_75t_L g10680 ( 
.A(n_9907),
.Y(n_10680)
);

INVx1_ASAP7_75t_L g10681 ( 
.A(n_9915),
.Y(n_10681)
);

INVx1_ASAP7_75t_L g10682 ( 
.A(n_10033),
.Y(n_10682)
);

NOR2xp33_ASAP7_75t_L g10683 ( 
.A(n_9880),
.B(n_4407),
.Y(n_10683)
);

AOI22xp5_ASAP7_75t_L g10684 ( 
.A1(n_9768),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_10684)
);

AO22x2_ASAP7_75t_L g10685 ( 
.A1(n_10022),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_10685)
);

INVx2_ASAP7_75t_L g10686 ( 
.A(n_10179),
.Y(n_10686)
);

INVx1_ASAP7_75t_L g10687 ( 
.A(n_9881),
.Y(n_10687)
);

NAND2xp5_ASAP7_75t_L g10688 ( 
.A(n_9966),
.B(n_216),
.Y(n_10688)
);

INVx1_ASAP7_75t_L g10689 ( 
.A(n_10024),
.Y(n_10689)
);

INVx1_ASAP7_75t_L g10690 ( 
.A(n_10094),
.Y(n_10690)
);

CKINVDCx5p33_ASAP7_75t_R g10691 ( 
.A(n_10049),
.Y(n_10691)
);

AO22x2_ASAP7_75t_L g10692 ( 
.A1(n_10028),
.A2(n_220),
.B1(n_217),
.B2(n_219),
.Y(n_10692)
);

AO22x2_ASAP7_75t_L g10693 ( 
.A1(n_9783),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_10693)
);

INVx1_ASAP7_75t_L g10694 ( 
.A(n_9790),
.Y(n_10694)
);

BUFx8_ASAP7_75t_L g10695 ( 
.A(n_10092),
.Y(n_10695)
);

BUFx2_ASAP7_75t_L g10696 ( 
.A(n_9907),
.Y(n_10696)
);

INVx5_ASAP7_75t_L g10697 ( 
.A(n_10176),
.Y(n_10697)
);

INVxp67_ASAP7_75t_L g10698 ( 
.A(n_9776),
.Y(n_10698)
);

INVx3_ASAP7_75t_L g10699 ( 
.A(n_9847),
.Y(n_10699)
);

INVx2_ASAP7_75t_L g10700 ( 
.A(n_10166),
.Y(n_10700)
);

INVxp67_ASAP7_75t_L g10701 ( 
.A(n_9951),
.Y(n_10701)
);

INVx1_ASAP7_75t_L g10702 ( 
.A(n_9798),
.Y(n_10702)
);

INVxp67_ASAP7_75t_L g10703 ( 
.A(n_9924),
.Y(n_10703)
);

AO22x2_ASAP7_75t_L g10704 ( 
.A1(n_9851),
.A2(n_224),
.B1(n_221),
.B2(n_223),
.Y(n_10704)
);

INVx1_ASAP7_75t_L g10705 ( 
.A(n_9942),
.Y(n_10705)
);

NAND2x1p5_ASAP7_75t_L g10706 ( 
.A(n_10143),
.B(n_4408),
.Y(n_10706)
);

INVx1_ASAP7_75t_L g10707 ( 
.A(n_10146),
.Y(n_10707)
);

INVx1_ASAP7_75t_L g10708 ( 
.A(n_10148),
.Y(n_10708)
);

CKINVDCx16_ASAP7_75t_R g10709 ( 
.A(n_10070),
.Y(n_10709)
);

NAND2xp5_ASAP7_75t_L g10710 ( 
.A(n_9835),
.B(n_223),
.Y(n_10710)
);

INVx1_ASAP7_75t_L g10711 ( 
.A(n_10149),
.Y(n_10711)
);

BUFx8_ASAP7_75t_L g10712 ( 
.A(n_10154),
.Y(n_10712)
);

INVx1_ASAP7_75t_L g10713 ( 
.A(n_10071),
.Y(n_10713)
);

INVx1_ASAP7_75t_L g10714 ( 
.A(n_10091),
.Y(n_10714)
);

BUFx8_ASAP7_75t_L g10715 ( 
.A(n_10085),
.Y(n_10715)
);

AND2x2_ASAP7_75t_L g10716 ( 
.A(n_9687),
.B(n_224),
.Y(n_10716)
);

INVxp33_ASAP7_75t_SL g10717 ( 
.A(n_10194),
.Y(n_10717)
);

INVx1_ASAP7_75t_L g10718 ( 
.A(n_9830),
.Y(n_10718)
);

AO22x2_ASAP7_75t_L g10719 ( 
.A1(n_9701),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_10719)
);

CKINVDCx5p33_ASAP7_75t_R g10720 ( 
.A(n_10194),
.Y(n_10720)
);

INVx1_ASAP7_75t_L g10721 ( 
.A(n_9830),
.Y(n_10721)
);

AO22x2_ASAP7_75t_L g10722 ( 
.A1(n_9701),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_10722)
);

NAND2xp5_ASAP7_75t_L g10723 ( 
.A(n_9719),
.B(n_228),
.Y(n_10723)
);

INVx1_ASAP7_75t_L g10724 ( 
.A(n_9830),
.Y(n_10724)
);

NAND2x1p5_ASAP7_75t_L g10725 ( 
.A(n_10198),
.B(n_4410),
.Y(n_10725)
);

CKINVDCx20_ASAP7_75t_R g10726 ( 
.A(n_10194),
.Y(n_10726)
);

AND2x2_ASAP7_75t_L g10727 ( 
.A(n_9687),
.B(n_229),
.Y(n_10727)
);

INVx1_ASAP7_75t_L g10728 ( 
.A(n_9830),
.Y(n_10728)
);

AO22x2_ASAP7_75t_L g10729 ( 
.A1(n_9701),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_10729)
);

INVxp67_ASAP7_75t_L g10730 ( 
.A(n_9694),
.Y(n_10730)
);

INVx1_ASAP7_75t_L g10731 ( 
.A(n_9830),
.Y(n_10731)
);

INVx2_ASAP7_75t_L g10732 ( 
.A(n_9762),
.Y(n_10732)
);

AO22x2_ASAP7_75t_L g10733 ( 
.A1(n_9701),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_10733)
);

OAI221xp5_ASAP7_75t_L g10734 ( 
.A1(n_9849),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.C(n_236),
.Y(n_10734)
);

INVxp67_ASAP7_75t_L g10735 ( 
.A(n_9694),
.Y(n_10735)
);

OAI221xp5_ASAP7_75t_L g10736 ( 
.A1(n_9849),
.A2(n_238),
.B1(n_234),
.B2(n_237),
.C(n_239),
.Y(n_10736)
);

NAND2x1p5_ASAP7_75t_L g10737 ( 
.A(n_10198),
.B(n_4411),
.Y(n_10737)
);

NAND2xp5_ASAP7_75t_L g10738 ( 
.A(n_9719),
.B(n_237),
.Y(n_10738)
);

INVx2_ASAP7_75t_L g10739 ( 
.A(n_9762),
.Y(n_10739)
);

NOR2xp33_ASAP7_75t_L g10740 ( 
.A(n_9691),
.B(n_4412),
.Y(n_10740)
);

BUFx6f_ASAP7_75t_SL g10741 ( 
.A(n_9733),
.Y(n_10741)
);

INVx1_ASAP7_75t_L g10742 ( 
.A(n_9830),
.Y(n_10742)
);

INVx1_ASAP7_75t_L g10743 ( 
.A(n_9830),
.Y(n_10743)
);

INVx1_ASAP7_75t_L g10744 ( 
.A(n_9830),
.Y(n_10744)
);

INVxp67_ASAP7_75t_L g10745 ( 
.A(n_9694),
.Y(n_10745)
);

NAND2xp5_ASAP7_75t_L g10746 ( 
.A(n_9719),
.B(n_238),
.Y(n_10746)
);

AND2x4_ASAP7_75t_L g10747 ( 
.A(n_9823),
.B(n_4413),
.Y(n_10747)
);

BUFx6f_ASAP7_75t_SL g10748 ( 
.A(n_9733),
.Y(n_10748)
);

CKINVDCx5p33_ASAP7_75t_R g10749 ( 
.A(n_10194),
.Y(n_10749)
);

INVx2_ASAP7_75t_L g10750 ( 
.A(n_9762),
.Y(n_10750)
);

INVx2_ASAP7_75t_L g10751 ( 
.A(n_9762),
.Y(n_10751)
);

INVx1_ASAP7_75t_L g10752 ( 
.A(n_9830),
.Y(n_10752)
);

NAND2xp5_ASAP7_75t_L g10753 ( 
.A(n_9719),
.B(n_239),
.Y(n_10753)
);

NAND2xp5_ASAP7_75t_L g10754 ( 
.A(n_9719),
.B(n_240),
.Y(n_10754)
);

INVx2_ASAP7_75t_L g10755 ( 
.A(n_9762),
.Y(n_10755)
);

CKINVDCx20_ASAP7_75t_R g10756 ( 
.A(n_10194),
.Y(n_10756)
);

INVx1_ASAP7_75t_L g10757 ( 
.A(n_9830),
.Y(n_10757)
);

NAND2xp5_ASAP7_75t_L g10758 ( 
.A(n_9719),
.B(n_240),
.Y(n_10758)
);

NAND2xp5_ASAP7_75t_L g10759 ( 
.A(n_9719),
.B(n_241),
.Y(n_10759)
);

OAI221xp5_ASAP7_75t_L g10760 ( 
.A1(n_9849),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.C(n_244),
.Y(n_10760)
);

NAND2xp5_ASAP7_75t_L g10761 ( 
.A(n_9719),
.B(n_242),
.Y(n_10761)
);

AND2x4_ASAP7_75t_L g10762 ( 
.A(n_9823),
.B(n_4414),
.Y(n_10762)
);

AO22x1_ASAP7_75t_L g10763 ( 
.A1(n_9691),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_10763)
);

NAND2xp5_ASAP7_75t_L g10764 ( 
.A(n_9719),
.B(n_245),
.Y(n_10764)
);

AO22x2_ASAP7_75t_L g10765 ( 
.A1(n_9701),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_10765)
);

INVxp67_ASAP7_75t_L g10766 ( 
.A(n_9694),
.Y(n_10766)
);

OA22x2_ASAP7_75t_L g10767 ( 
.A1(n_9782),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_10767)
);

HB1xp67_ASAP7_75t_L g10768 ( 
.A(n_9694),
.Y(n_10768)
);

AO22x2_ASAP7_75t_L g10769 ( 
.A1(n_9701),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_10769)
);

NAND2xp5_ASAP7_75t_L g10770 ( 
.A(n_9719),
.B(n_251),
.Y(n_10770)
);

NAND2xp5_ASAP7_75t_L g10771 ( 
.A(n_9719),
.B(n_253),
.Y(n_10771)
);

AO22x2_ASAP7_75t_L g10772 ( 
.A1(n_9701),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_10772)
);

INVxp67_ASAP7_75t_SL g10773 ( 
.A(n_9846),
.Y(n_10773)
);

INVx1_ASAP7_75t_L g10774 ( 
.A(n_9830),
.Y(n_10774)
);

NAND2xp5_ASAP7_75t_L g10775 ( 
.A(n_9719),
.B(n_256),
.Y(n_10775)
);

AND2x4_ASAP7_75t_L g10776 ( 
.A(n_9823),
.B(n_4415),
.Y(n_10776)
);

NAND2xp5_ASAP7_75t_L g10777 ( 
.A(n_9719),
.B(n_257),
.Y(n_10777)
);

AOI22xp5_ASAP7_75t_L g10778 ( 
.A1(n_9691),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_10778)
);

INVx1_ASAP7_75t_L g10779 ( 
.A(n_9830),
.Y(n_10779)
);

CKINVDCx20_ASAP7_75t_R g10780 ( 
.A(n_10194),
.Y(n_10780)
);

CKINVDCx5p33_ASAP7_75t_R g10781 ( 
.A(n_10194),
.Y(n_10781)
);

INVx1_ASAP7_75t_L g10782 ( 
.A(n_9830),
.Y(n_10782)
);

AOI22xp5_ASAP7_75t_L g10783 ( 
.A1(n_9691),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_10783)
);

INVx1_ASAP7_75t_L g10784 ( 
.A(n_9830),
.Y(n_10784)
);

INVx1_ASAP7_75t_L g10785 ( 
.A(n_9830),
.Y(n_10785)
);

INVx1_ASAP7_75t_L g10786 ( 
.A(n_9830),
.Y(n_10786)
);

AO22x2_ASAP7_75t_L g10787 ( 
.A1(n_9701),
.A2(n_263),
.B1(n_260),
.B2(n_262),
.Y(n_10787)
);

INVxp67_ASAP7_75t_L g10788 ( 
.A(n_9694),
.Y(n_10788)
);

CKINVDCx5p33_ASAP7_75t_R g10789 ( 
.A(n_10194),
.Y(n_10789)
);

INVx2_ASAP7_75t_L g10790 ( 
.A(n_9762),
.Y(n_10790)
);

INVx2_ASAP7_75t_L g10791 ( 
.A(n_9762),
.Y(n_10791)
);

HB1xp67_ASAP7_75t_L g10792 ( 
.A(n_9694),
.Y(n_10792)
);

NAND2xp5_ASAP7_75t_SL g10793 ( 
.A(n_9782),
.B(n_262),
.Y(n_10793)
);

CKINVDCx5p33_ASAP7_75t_R g10794 ( 
.A(n_10194),
.Y(n_10794)
);

HB1xp67_ASAP7_75t_L g10795 ( 
.A(n_9694),
.Y(n_10795)
);

AND2x2_ASAP7_75t_SL g10796 ( 
.A(n_9691),
.B(n_264),
.Y(n_10796)
);

INVx1_ASAP7_75t_L g10797 ( 
.A(n_9830),
.Y(n_10797)
);

AO22x2_ASAP7_75t_L g10798 ( 
.A1(n_9701),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_10798)
);

NAND2xp5_ASAP7_75t_L g10799 ( 
.A(n_9719),
.B(n_265),
.Y(n_10799)
);

INVx1_ASAP7_75t_L g10800 ( 
.A(n_9830),
.Y(n_10800)
);

INVxp67_ASAP7_75t_L g10801 ( 
.A(n_9694),
.Y(n_10801)
);

INVx1_ASAP7_75t_L g10802 ( 
.A(n_9830),
.Y(n_10802)
);

INVx1_ASAP7_75t_L g10803 ( 
.A(n_9830),
.Y(n_10803)
);

BUFx8_ASAP7_75t_L g10804 ( 
.A(n_10085),
.Y(n_10804)
);

AND2x6_ASAP7_75t_L g10805 ( 
.A(n_9737),
.B(n_4416),
.Y(n_10805)
);

INVx1_ASAP7_75t_L g10806 ( 
.A(n_9830),
.Y(n_10806)
);

AO22x2_ASAP7_75t_L g10807 ( 
.A1(n_9701),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_10807)
);

INVx1_ASAP7_75t_L g10808 ( 
.A(n_9830),
.Y(n_10808)
);

AND2x4_ASAP7_75t_L g10809 ( 
.A(n_9823),
.B(n_4417),
.Y(n_10809)
);

INVx2_ASAP7_75t_SL g10810 ( 
.A(n_9730),
.Y(n_10810)
);

INVx1_ASAP7_75t_L g10811 ( 
.A(n_9830),
.Y(n_10811)
);

AOI22xp5_ASAP7_75t_L g10812 ( 
.A1(n_9691),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_10812)
);

AO22x2_ASAP7_75t_L g10813 ( 
.A1(n_9701),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_10813)
);

INVx1_ASAP7_75t_L g10814 ( 
.A(n_9830),
.Y(n_10814)
);

OAI22xp5_ASAP7_75t_L g10815 ( 
.A1(n_9691),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_10815)
);

INVx1_ASAP7_75t_L g10816 ( 
.A(n_9830),
.Y(n_10816)
);

OAI22xp5_ASAP7_75t_L g10817 ( 
.A1(n_9691),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_10817)
);

INVx1_ASAP7_75t_L g10818 ( 
.A(n_9830),
.Y(n_10818)
);

INVx1_ASAP7_75t_L g10819 ( 
.A(n_9830),
.Y(n_10819)
);

AO22x2_ASAP7_75t_L g10820 ( 
.A1(n_9701),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_10820)
);

HB1xp67_ASAP7_75t_L g10821 ( 
.A(n_9694),
.Y(n_10821)
);

INVx1_ASAP7_75t_L g10822 ( 
.A(n_9830),
.Y(n_10822)
);

INVx1_ASAP7_75t_L g10823 ( 
.A(n_9830),
.Y(n_10823)
);

AOI21xp5_ASAP7_75t_L g10824 ( 
.A1(n_10324),
.A2(n_4419),
.B(n_4418),
.Y(n_10824)
);

AOI21xp5_ASAP7_75t_L g10825 ( 
.A1(n_10229),
.A2(n_4421),
.B(n_4420),
.Y(n_10825)
);

NOR3xp33_ASAP7_75t_L g10826 ( 
.A(n_10276),
.B(n_10501),
.C(n_10288),
.Y(n_10826)
);

NAND2xp5_ASAP7_75t_L g10827 ( 
.A(n_10532),
.B(n_276),
.Y(n_10827)
);

OAI21xp5_ASAP7_75t_L g10828 ( 
.A1(n_10515),
.A2(n_277),
.B(n_278),
.Y(n_10828)
);

INVx1_ASAP7_75t_L g10829 ( 
.A(n_10291),
.Y(n_10829)
);

NAND2xp5_ASAP7_75t_L g10830 ( 
.A(n_10533),
.B(n_277),
.Y(n_10830)
);

AOI22xp33_ASAP7_75t_L g10831 ( 
.A1(n_10308),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_10831)
);

AOI21x1_ASAP7_75t_L g10832 ( 
.A1(n_10392),
.A2(n_4424),
.B(n_4423),
.Y(n_10832)
);

INVx2_ASAP7_75t_L g10833 ( 
.A(n_10220),
.Y(n_10833)
);

INVx1_ASAP7_75t_L g10834 ( 
.A(n_10294),
.Y(n_10834)
);

AOI21xp5_ASAP7_75t_L g10835 ( 
.A1(n_10624),
.A2(n_4427),
.B(n_4426),
.Y(n_10835)
);

O2A1O1Ixp33_ASAP7_75t_L g10836 ( 
.A1(n_10323),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_10836)
);

AOI21xp5_ASAP7_75t_L g10837 ( 
.A1(n_10457),
.A2(n_4430),
.B(n_4428),
.Y(n_10837)
);

OAI22xp5_ASAP7_75t_L g10838 ( 
.A1(n_10280),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_10838)
);

AOI21xp5_ASAP7_75t_L g10839 ( 
.A1(n_10347),
.A2(n_10242),
.B(n_10531),
.Y(n_10839)
);

O2A1O1Ixp33_ASAP7_75t_L g10840 ( 
.A1(n_10366),
.A2(n_285),
.B(n_282),
.C(n_284),
.Y(n_10840)
);

NAND2xp5_ASAP7_75t_L g10841 ( 
.A(n_10535),
.B(n_285),
.Y(n_10841)
);

AOI21xp5_ASAP7_75t_L g10842 ( 
.A1(n_10274),
.A2(n_4432),
.B(n_4431),
.Y(n_10842)
);

AOI21xp5_ASAP7_75t_L g10843 ( 
.A1(n_10258),
.A2(n_4434),
.B(n_4433),
.Y(n_10843)
);

NAND2xp5_ASAP7_75t_L g10844 ( 
.A(n_10536),
.B(n_286),
.Y(n_10844)
);

NAND2xp5_ASAP7_75t_L g10845 ( 
.A(n_10538),
.B(n_286),
.Y(n_10845)
);

AND2x6_ASAP7_75t_L g10846 ( 
.A(n_10598),
.B(n_4435),
.Y(n_10846)
);

A2O1A1Ixp33_ASAP7_75t_L g10847 ( 
.A1(n_10740),
.A2(n_289),
.B(n_287),
.C(n_288),
.Y(n_10847)
);

AND2x4_ASAP7_75t_L g10848 ( 
.A(n_10380),
.B(n_4437),
.Y(n_10848)
);

OAI22xp5_ASAP7_75t_L g10849 ( 
.A1(n_10411),
.A2(n_290),
.B1(n_287),
.B2(n_288),
.Y(n_10849)
);

NAND2xp5_ASAP7_75t_SL g10850 ( 
.A(n_10541),
.B(n_4438),
.Y(n_10850)
);

AOI21xp5_ASAP7_75t_L g10851 ( 
.A1(n_10773),
.A2(n_4441),
.B(n_4439),
.Y(n_10851)
);

INVxp67_ASAP7_75t_L g10852 ( 
.A(n_10217),
.Y(n_10852)
);

BUFx4f_ASAP7_75t_L g10853 ( 
.A(n_10267),
.Y(n_10853)
);

O2A1O1Ixp33_ASAP7_75t_L g10854 ( 
.A1(n_10793),
.A2(n_292),
.B(n_290),
.C(n_291),
.Y(n_10854)
);

AOI21xp5_ASAP7_75t_L g10855 ( 
.A1(n_10337),
.A2(n_10343),
.B(n_10644),
.Y(n_10855)
);

INVx1_ASAP7_75t_SL g10856 ( 
.A(n_10215),
.Y(n_10856)
);

AND2x4_ASAP7_75t_L g10857 ( 
.A(n_10446),
.B(n_4442),
.Y(n_10857)
);

NOR2xp33_ASAP7_75t_SL g10858 ( 
.A(n_10717),
.B(n_4443),
.Y(n_10858)
);

AND2x2_ASAP7_75t_L g10859 ( 
.A(n_10310),
.B(n_10623),
.Y(n_10859)
);

AOI21xp5_ASAP7_75t_L g10860 ( 
.A1(n_10207),
.A2(n_4446),
.B(n_4445),
.Y(n_10860)
);

AOI21xp5_ASAP7_75t_L g10861 ( 
.A1(n_10208),
.A2(n_4448),
.B(n_4447),
.Y(n_10861)
);

AOI21xp5_ASAP7_75t_L g10862 ( 
.A1(n_10212),
.A2(n_4450),
.B(n_4449),
.Y(n_10862)
);

NAND2xp5_ASAP7_75t_L g10863 ( 
.A(n_10543),
.B(n_291),
.Y(n_10863)
);

NAND2xp5_ASAP7_75t_SL g10864 ( 
.A(n_10550),
.B(n_4451),
.Y(n_10864)
);

NAND2xp5_ASAP7_75t_L g10865 ( 
.A(n_10551),
.B(n_292),
.Y(n_10865)
);

INVx1_ASAP7_75t_L g10866 ( 
.A(n_10295),
.Y(n_10866)
);

NAND2xp5_ASAP7_75t_L g10867 ( 
.A(n_10554),
.B(n_293),
.Y(n_10867)
);

AOI21xp5_ASAP7_75t_L g10868 ( 
.A1(n_10718),
.A2(n_4453),
.B(n_4452),
.Y(n_10868)
);

AOI21xp5_ASAP7_75t_L g10869 ( 
.A1(n_10721),
.A2(n_4455),
.B(n_4454),
.Y(n_10869)
);

NAND2xp5_ASAP7_75t_L g10870 ( 
.A(n_10555),
.B(n_10556),
.Y(n_10870)
);

NOR2xp33_ASAP7_75t_L g10871 ( 
.A(n_10315),
.B(n_4456),
.Y(n_10871)
);

AO22x1_ASAP7_75t_L g10872 ( 
.A1(n_10223),
.A2(n_10805),
.B1(n_10695),
.B2(n_10674),
.Y(n_10872)
);

OAI22xp5_ASAP7_75t_L g10873 ( 
.A1(n_10463),
.A2(n_297),
.B1(n_293),
.B2(n_294),
.Y(n_10873)
);

AOI21xp5_ASAP7_75t_L g10874 ( 
.A1(n_10724),
.A2(n_4459),
.B(n_4457),
.Y(n_10874)
);

BUFx2_ASAP7_75t_L g10875 ( 
.A(n_10249),
.Y(n_10875)
);

AOI21xp5_ASAP7_75t_L g10876 ( 
.A1(n_10728),
.A2(n_4462),
.B(n_4461),
.Y(n_10876)
);

O2A1O1Ixp33_ASAP7_75t_L g10877 ( 
.A1(n_10300),
.A2(n_298),
.B(n_294),
.C(n_297),
.Y(n_10877)
);

AOI22xp33_ASAP7_75t_L g10878 ( 
.A1(n_10796),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_10878)
);

BUFx12f_ASAP7_75t_L g10879 ( 
.A(n_10382),
.Y(n_10879)
);

AOI22xp5_ASAP7_75t_L g10880 ( 
.A1(n_10709),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_10880)
);

AOI21x1_ASAP7_75t_L g10881 ( 
.A1(n_10587),
.A2(n_4464),
.B(n_4463),
.Y(n_10881)
);

NAND2xp5_ASAP7_75t_L g10882 ( 
.A(n_10557),
.B(n_301),
.Y(n_10882)
);

AOI21xp5_ASAP7_75t_L g10883 ( 
.A1(n_10731),
.A2(n_4469),
.B(n_4468),
.Y(n_10883)
);

INVx1_ASAP7_75t_SL g10884 ( 
.A(n_10254),
.Y(n_10884)
);

OAI22xp5_ASAP7_75t_L g10885 ( 
.A1(n_10465),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_10885)
);

OAI21xp33_ASAP7_75t_L g10886 ( 
.A1(n_10653),
.A2(n_302),
.B(n_304),
.Y(n_10886)
);

INVx3_ASAP7_75t_L g10887 ( 
.A(n_10227),
.Y(n_10887)
);

AOI21xp5_ASAP7_75t_L g10888 ( 
.A1(n_10742),
.A2(n_4471),
.B(n_4470),
.Y(n_10888)
);

AOI21xp5_ASAP7_75t_L g10889 ( 
.A1(n_10743),
.A2(n_4473),
.B(n_4472),
.Y(n_10889)
);

AOI21xp5_ASAP7_75t_L g10890 ( 
.A1(n_10744),
.A2(n_4478),
.B(n_4477),
.Y(n_10890)
);

INVx2_ASAP7_75t_L g10891 ( 
.A(n_10257),
.Y(n_10891)
);

INVxp67_ASAP7_75t_L g10892 ( 
.A(n_10768),
.Y(n_10892)
);

O2A1O1Ixp33_ASAP7_75t_L g10893 ( 
.A1(n_10221),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_10893)
);

OAI22xp5_ASAP7_75t_L g10894 ( 
.A1(n_10659),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.Y(n_10894)
);

OAI22xp5_ASAP7_75t_L g10895 ( 
.A1(n_10464),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_10895)
);

NOR2xp33_ASAP7_75t_L g10896 ( 
.A(n_10452),
.B(n_4479),
.Y(n_10896)
);

AOI21xp5_ASAP7_75t_L g10897 ( 
.A1(n_10752),
.A2(n_4481),
.B(n_4480),
.Y(n_10897)
);

NAND2xp5_ASAP7_75t_L g10898 ( 
.A(n_10558),
.B(n_310),
.Y(n_10898)
);

NAND2xp5_ASAP7_75t_L g10899 ( 
.A(n_10559),
.B(n_311),
.Y(n_10899)
);

NAND2xp5_ASAP7_75t_SL g10900 ( 
.A(n_10560),
.B(n_4482),
.Y(n_10900)
);

AND2x2_ASAP7_75t_L g10901 ( 
.A(n_10281),
.B(n_4483),
.Y(n_10901)
);

NAND2xp33_ASAP7_75t_SL g10902 ( 
.A(n_10350),
.B(n_311),
.Y(n_10902)
);

INVx2_ASAP7_75t_L g10903 ( 
.A(n_10278),
.Y(n_10903)
);

A2O1A1Ixp33_ASAP7_75t_L g10904 ( 
.A1(n_10679),
.A2(n_10612),
.B(n_10713),
.C(n_10290),
.Y(n_10904)
);

BUFx6f_ASAP7_75t_L g10905 ( 
.A(n_10318),
.Y(n_10905)
);

AOI21xp5_ASAP7_75t_L g10906 ( 
.A1(n_10757),
.A2(n_4487),
.B(n_4484),
.Y(n_10906)
);

BUFx2_ASAP7_75t_L g10907 ( 
.A(n_10792),
.Y(n_10907)
);

AND2x4_ASAP7_75t_L g10908 ( 
.A(n_10660),
.B(n_4488),
.Y(n_10908)
);

NAND2x1p5_ASAP7_75t_L g10909 ( 
.A(n_10283),
.B(n_4489),
.Y(n_10909)
);

AOI21xp5_ASAP7_75t_L g10910 ( 
.A1(n_10774),
.A2(n_4491),
.B(n_4490),
.Y(n_10910)
);

AOI21x1_ASAP7_75t_L g10911 ( 
.A1(n_10301),
.A2(n_4493),
.B(n_4492),
.Y(n_10911)
);

INVx1_ASAP7_75t_L g10912 ( 
.A(n_10299),
.Y(n_10912)
);

AOI21xp5_ASAP7_75t_L g10913 ( 
.A1(n_10779),
.A2(n_4498),
.B(n_4494),
.Y(n_10913)
);

NAND2xp5_ASAP7_75t_L g10914 ( 
.A(n_10561),
.B(n_312),
.Y(n_10914)
);

OAI21xp33_ASAP7_75t_L g10915 ( 
.A1(n_10317),
.A2(n_313),
.B(n_314),
.Y(n_10915)
);

NAND2xp5_ASAP7_75t_L g10916 ( 
.A(n_10566),
.B(n_10567),
.Y(n_10916)
);

INVx1_ASAP7_75t_L g10917 ( 
.A(n_10305),
.Y(n_10917)
);

AOI21xp5_ASAP7_75t_L g10918 ( 
.A1(n_10782),
.A2(n_4500),
.B(n_4499),
.Y(n_10918)
);

CKINVDCx8_ASAP7_75t_R g10919 ( 
.A(n_10283),
.Y(n_10919)
);

NAND2xp5_ASAP7_75t_SL g10920 ( 
.A(n_10569),
.B(n_10570),
.Y(n_10920)
);

NAND2xp5_ASAP7_75t_L g10921 ( 
.A(n_10573),
.B(n_313),
.Y(n_10921)
);

AOI21xp5_ASAP7_75t_L g10922 ( 
.A1(n_10784),
.A2(n_4502),
.B(n_4501),
.Y(n_10922)
);

NAND2xp5_ASAP7_75t_L g10923 ( 
.A(n_10785),
.B(n_314),
.Y(n_10923)
);

BUFx2_ASAP7_75t_L g10924 ( 
.A(n_10795),
.Y(n_10924)
);

OAI21xp5_ASAP7_75t_L g10925 ( 
.A1(n_10603),
.A2(n_315),
.B(n_316),
.Y(n_10925)
);

INVx2_ASAP7_75t_L g10926 ( 
.A(n_10287),
.Y(n_10926)
);

NAND2xp5_ASAP7_75t_L g10927 ( 
.A(n_10786),
.B(n_315),
.Y(n_10927)
);

OAI22xp5_ASAP7_75t_SL g10928 ( 
.A1(n_10497),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_10928)
);

AOI21x1_ASAP7_75t_L g10929 ( 
.A1(n_10477),
.A2(n_10394),
.B(n_10594),
.Y(n_10929)
);

OAI21xp5_ASAP7_75t_L g10930 ( 
.A1(n_10604),
.A2(n_317),
.B(n_318),
.Y(n_10930)
);

AOI21xp5_ASAP7_75t_L g10931 ( 
.A1(n_10797),
.A2(n_4504),
.B(n_4503),
.Y(n_10931)
);

AOI21xp5_ASAP7_75t_L g10932 ( 
.A1(n_10800),
.A2(n_4506),
.B(n_4505),
.Y(n_10932)
);

OAI22xp5_ASAP7_75t_L g10933 ( 
.A1(n_10664),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_10933)
);

AOI21xp5_ASAP7_75t_L g10934 ( 
.A1(n_10802),
.A2(n_4509),
.B(n_4508),
.Y(n_10934)
);

O2A1O1Ixp33_ASAP7_75t_L g10935 ( 
.A1(n_10365),
.A2(n_322),
.B(n_320),
.C(n_321),
.Y(n_10935)
);

NAND2xp5_ASAP7_75t_L g10936 ( 
.A(n_10803),
.B(n_322),
.Y(n_10936)
);

NAND2xp5_ASAP7_75t_L g10937 ( 
.A(n_10806),
.B(n_323),
.Y(n_10937)
);

AOI21xp5_ASAP7_75t_L g10938 ( 
.A1(n_10808),
.A2(n_4511),
.B(n_4510),
.Y(n_10938)
);

AOI21xp5_ASAP7_75t_L g10939 ( 
.A1(n_10811),
.A2(n_4514),
.B(n_4513),
.Y(n_10939)
);

AOI22x1_ASAP7_75t_L g10940 ( 
.A1(n_10211),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_10940)
);

OAI22xp5_ASAP7_75t_L g10941 ( 
.A1(n_10507),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_10941)
);

AOI21xp5_ASAP7_75t_L g10942 ( 
.A1(n_10814),
.A2(n_4517),
.B(n_4515),
.Y(n_10942)
);

NAND2xp5_ASAP7_75t_L g10943 ( 
.A(n_10816),
.B(n_326),
.Y(n_10943)
);

BUFx6f_ASAP7_75t_L g10944 ( 
.A(n_10318),
.Y(n_10944)
);

AOI21xp5_ASAP7_75t_L g10945 ( 
.A1(n_10818),
.A2(n_10822),
.B(n_10819),
.Y(n_10945)
);

AOI21xp5_ASAP7_75t_L g10946 ( 
.A1(n_10823),
.A2(n_4519),
.B(n_4518),
.Y(n_10946)
);

NOR2xp33_ASAP7_75t_L g10947 ( 
.A(n_10451),
.B(n_4520),
.Y(n_10947)
);

INVx1_ASAP7_75t_L g10948 ( 
.A(n_10306),
.Y(n_10948)
);

HB1xp67_ASAP7_75t_L g10949 ( 
.A(n_10821),
.Y(n_10949)
);

AOI21xp5_ASAP7_75t_L g10950 ( 
.A1(n_10694),
.A2(n_4523),
.B(n_4521),
.Y(n_10950)
);

INVx1_ASAP7_75t_L g10951 ( 
.A(n_10311),
.Y(n_10951)
);

AOI21xp5_ASAP7_75t_L g10952 ( 
.A1(n_10577),
.A2(n_4525),
.B(n_4524),
.Y(n_10952)
);

AOI21xp5_ASAP7_75t_L g10953 ( 
.A1(n_10579),
.A2(n_4527),
.B(n_4526),
.Y(n_10953)
);

INVx1_ASAP7_75t_SL g10954 ( 
.A(n_10378),
.Y(n_10954)
);

AOI21xp5_ASAP7_75t_L g10955 ( 
.A1(n_10585),
.A2(n_4530),
.B(n_4528),
.Y(n_10955)
);

AOI21xp5_ASAP7_75t_L g10956 ( 
.A1(n_10467),
.A2(n_4533),
.B(n_4532),
.Y(n_10956)
);

AOI21xp5_ASAP7_75t_L g10957 ( 
.A1(n_10468),
.A2(n_4536),
.B(n_4534),
.Y(n_10957)
);

NAND2xp5_ASAP7_75t_L g10958 ( 
.A(n_10514),
.B(n_327),
.Y(n_10958)
);

HB1xp67_ASAP7_75t_L g10959 ( 
.A(n_10232),
.Y(n_10959)
);

AOI21xp5_ASAP7_75t_L g10960 ( 
.A1(n_10472),
.A2(n_4538),
.B(n_4537),
.Y(n_10960)
);

NAND2xp5_ASAP7_75t_L g10961 ( 
.A(n_10517),
.B(n_10520),
.Y(n_10961)
);

BUFx2_ASAP7_75t_L g10962 ( 
.A(n_10730),
.Y(n_10962)
);

BUFx3_ASAP7_75t_L g10963 ( 
.A(n_10540),
.Y(n_10963)
);

O2A1O1Ixp33_ASAP7_75t_L g10964 ( 
.A1(n_10351),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_10964)
);

OAI21xp5_ASAP7_75t_L g10965 ( 
.A1(n_10529),
.A2(n_328),
.B(n_329),
.Y(n_10965)
);

O2A1O1Ixp33_ASAP7_75t_SL g10966 ( 
.A1(n_10650),
.A2(n_332),
.B(n_330),
.C(n_331),
.Y(n_10966)
);

INVx1_ASAP7_75t_L g10967 ( 
.A(n_10316),
.Y(n_10967)
);

A2O1A1Ixp33_ASAP7_75t_L g10968 ( 
.A1(n_10714),
.A2(n_334),
.B(n_332),
.C(n_333),
.Y(n_10968)
);

AOI21xp5_ASAP7_75t_L g10969 ( 
.A1(n_10476),
.A2(n_10483),
.B(n_10481),
.Y(n_10969)
);

AOI21xp5_ASAP7_75t_L g10970 ( 
.A1(n_10484),
.A2(n_4540),
.B(n_4539),
.Y(n_10970)
);

NAND2xp5_ASAP7_75t_L g10971 ( 
.A(n_10521),
.B(n_333),
.Y(n_10971)
);

AOI21xp33_ASAP7_75t_L g10972 ( 
.A1(n_10690),
.A2(n_334),
.B(n_335),
.Y(n_10972)
);

NAND2xp5_ASAP7_75t_L g10973 ( 
.A(n_10525),
.B(n_335),
.Y(n_10973)
);

NAND2xp5_ASAP7_75t_L g10974 ( 
.A(n_10398),
.B(n_336),
.Y(n_10974)
);

AOI21xp5_ASAP7_75t_L g10975 ( 
.A1(n_10485),
.A2(n_4542),
.B(n_4541),
.Y(n_10975)
);

NAND2xp5_ASAP7_75t_SL g10976 ( 
.A(n_10699),
.B(n_4543),
.Y(n_10976)
);

A2O1A1Ixp33_ASAP7_75t_L g10977 ( 
.A1(n_10271),
.A2(n_339),
.B(n_337),
.C(n_338),
.Y(n_10977)
);

AOI21xp5_ASAP7_75t_L g10978 ( 
.A1(n_10492),
.A2(n_4545),
.B(n_4544),
.Y(n_10978)
);

INVxp67_ASAP7_75t_L g10979 ( 
.A(n_10339),
.Y(n_10979)
);

AOI21xp5_ASAP7_75t_L g10980 ( 
.A1(n_10495),
.A2(n_10503),
.B(n_10500),
.Y(n_10980)
);

BUFx2_ASAP7_75t_L g10981 ( 
.A(n_10735),
.Y(n_10981)
);

AOI21x1_ASAP7_75t_L g10982 ( 
.A1(n_10590),
.A2(n_4547),
.B(n_4546),
.Y(n_10982)
);

A2O1A1Ixp33_ASAP7_75t_L g10983 ( 
.A1(n_10277),
.A2(n_341),
.B(n_339),
.C(n_340),
.Y(n_10983)
);

INVx1_ASAP7_75t_SL g10984 ( 
.A(n_10412),
.Y(n_10984)
);

NAND2xp5_ASAP7_75t_L g10985 ( 
.A(n_10400),
.B(n_341),
.Y(n_10985)
);

AOI21xp5_ASAP7_75t_L g10986 ( 
.A1(n_10505),
.A2(n_4552),
.B(n_4549),
.Y(n_10986)
);

NAND2xp5_ASAP7_75t_SL g10987 ( 
.A(n_10506),
.B(n_4554),
.Y(n_10987)
);

NAND2x1_ASAP7_75t_L g10988 ( 
.A(n_10466),
.B(n_4556),
.Y(n_10988)
);

NAND2xp5_ASAP7_75t_L g10989 ( 
.A(n_10510),
.B(n_10511),
.Y(n_10989)
);

AOI21xp5_ASAP7_75t_L g10990 ( 
.A1(n_10513),
.A2(n_4558),
.B(n_4557),
.Y(n_10990)
);

BUFx6f_ASAP7_75t_L g10991 ( 
.A(n_10253),
.Y(n_10991)
);

OAI21xp5_ASAP7_75t_L g10992 ( 
.A1(n_10588),
.A2(n_342),
.B(n_343),
.Y(n_10992)
);

OR2x6_ASAP7_75t_L g10993 ( 
.A(n_10439),
.B(n_4559),
.Y(n_10993)
);

AOI21x1_ASAP7_75t_L g10994 ( 
.A1(n_10596),
.A2(n_4565),
.B(n_4561),
.Y(n_10994)
);

A2O1A1Ixp33_ASAP7_75t_L g10995 ( 
.A1(n_10241),
.A2(n_345),
.B(n_342),
.C(n_344),
.Y(n_10995)
);

AOI21xp5_ASAP7_75t_L g10996 ( 
.A1(n_10417),
.A2(n_4567),
.B(n_4566),
.Y(n_10996)
);

NOR2xp33_ASAP7_75t_L g10997 ( 
.A(n_10359),
.B(n_4569),
.Y(n_10997)
);

AOI21xp5_ASAP7_75t_L g10998 ( 
.A1(n_10615),
.A2(n_4571),
.B(n_4570),
.Y(n_10998)
);

AOI21xp5_ASAP7_75t_L g10999 ( 
.A1(n_10430),
.A2(n_4573),
.B(n_4572),
.Y(n_10999)
);

NAND2xp5_ASAP7_75t_L g11000 ( 
.A(n_10433),
.B(n_344),
.Y(n_11000)
);

AOI21xp5_ASAP7_75t_L g11001 ( 
.A1(n_10435),
.A2(n_4576),
.B(n_4575),
.Y(n_11001)
);

A2O1A1Ixp33_ASAP7_75t_L g11002 ( 
.A1(n_10256),
.A2(n_347),
.B(n_345),
.C(n_346),
.Y(n_11002)
);

AOI21xp5_ASAP7_75t_L g11003 ( 
.A1(n_10581),
.A2(n_10528),
.B(n_10469),
.Y(n_11003)
);

INVx3_ASAP7_75t_L g11004 ( 
.A(n_10473),
.Y(n_11004)
);

INVx2_ASAP7_75t_L g11005 ( 
.A(n_10391),
.Y(n_11005)
);

INVx2_ASAP7_75t_L g11006 ( 
.A(n_10732),
.Y(n_11006)
);

AOI21xp5_ASAP7_75t_L g11007 ( 
.A1(n_10537),
.A2(n_4578),
.B(n_4577),
.Y(n_11007)
);

INVx3_ASAP7_75t_L g11008 ( 
.A(n_10356),
.Y(n_11008)
);

NAND2xp33_ASAP7_75t_L g11009 ( 
.A(n_10676),
.B(n_347),
.Y(n_11009)
);

INVx1_ASAP7_75t_L g11010 ( 
.A(n_10325),
.Y(n_11010)
);

INVx1_ASAP7_75t_L g11011 ( 
.A(n_10326),
.Y(n_11011)
);

AOI21xp5_ASAP7_75t_L g11012 ( 
.A1(n_10545),
.A2(n_4581),
.B(n_4579),
.Y(n_11012)
);

OAI22xp5_ASAP7_75t_L g11013 ( 
.A1(n_10698),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_11013)
);

NAND2xp5_ASAP7_75t_L g11014 ( 
.A(n_10210),
.B(n_10279),
.Y(n_11014)
);

HB1xp67_ASAP7_75t_L g11015 ( 
.A(n_10341),
.Y(n_11015)
);

AOI22xp5_ASAP7_75t_L g11016 ( 
.A1(n_10656),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_11016)
);

BUFx2_ASAP7_75t_L g11017 ( 
.A(n_10745),
.Y(n_11017)
);

INVx2_ASAP7_75t_L g11018 ( 
.A(n_10739),
.Y(n_11018)
);

A2O1A1Ixp33_ASAP7_75t_L g11019 ( 
.A1(n_10206),
.A2(n_10738),
.B(n_10746),
.C(n_10723),
.Y(n_11019)
);

NAND2xp5_ASAP7_75t_L g11020 ( 
.A(n_10346),
.B(n_352),
.Y(n_11020)
);

AOI22xp33_ASAP7_75t_L g11021 ( 
.A1(n_10621),
.A2(n_10648),
.B1(n_10405),
.B2(n_10226),
.Y(n_11021)
);

AO21x1_ASAP7_75t_L g11022 ( 
.A1(n_10386),
.A2(n_352),
.B(n_353),
.Y(n_11022)
);

NOR2xp33_ASAP7_75t_L g11023 ( 
.A(n_10703),
.B(n_4582),
.Y(n_11023)
);

AOI21xp5_ASAP7_75t_L g11024 ( 
.A1(n_10568),
.A2(n_4584),
.B(n_4583),
.Y(n_11024)
);

INVx2_ASAP7_75t_SL g11025 ( 
.A(n_10267),
.Y(n_11025)
);

NAND2xp5_ASAP7_75t_L g11026 ( 
.A(n_10766),
.B(n_353),
.Y(n_11026)
);

NOR2xp67_ASAP7_75t_L g11027 ( 
.A(n_10697),
.B(n_4585),
.Y(n_11027)
);

NAND2xp5_ASAP7_75t_L g11028 ( 
.A(n_10788),
.B(n_354),
.Y(n_11028)
);

AND2x4_ASAP7_75t_L g11029 ( 
.A(n_10460),
.B(n_4586),
.Y(n_11029)
);

NAND2xp5_ASAP7_75t_L g11030 ( 
.A(n_10801),
.B(n_354),
.Y(n_11030)
);

NOR2xp33_ASAP7_75t_L g11031 ( 
.A(n_10701),
.B(n_4587),
.Y(n_11031)
);

AOI21xp5_ASAP7_75t_L g11032 ( 
.A1(n_10626),
.A2(n_4589),
.B(n_4588),
.Y(n_11032)
);

AOI221xp5_ASAP7_75t_SL g11033 ( 
.A1(n_10815),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.C(n_358),
.Y(n_11033)
);

AOI21xp5_ASAP7_75t_L g11034 ( 
.A1(n_10820),
.A2(n_10722),
.B(n_10719),
.Y(n_11034)
);

AND2x2_ASAP7_75t_L g11035 ( 
.A(n_10307),
.B(n_4590),
.Y(n_11035)
);

NAND2xp5_ASAP7_75t_L g11036 ( 
.A(n_10753),
.B(n_355),
.Y(n_11036)
);

OAI21xp33_ASAP7_75t_L g11037 ( 
.A1(n_10321),
.A2(n_356),
.B(n_357),
.Y(n_11037)
);

A2O1A1Ixp33_ASAP7_75t_L g11038 ( 
.A1(n_10754),
.A2(n_361),
.B(n_359),
.C(n_360),
.Y(n_11038)
);

NAND2xp5_ASAP7_75t_L g11039 ( 
.A(n_10758),
.B(n_359),
.Y(n_11039)
);

AOI21xp5_ASAP7_75t_L g11040 ( 
.A1(n_10729),
.A2(n_4592),
.B(n_4591),
.Y(n_11040)
);

OAI21xp5_ASAP7_75t_L g11041 ( 
.A1(n_10710),
.A2(n_360),
.B(n_361),
.Y(n_11041)
);

AND3x2_ASAP7_75t_L g11042 ( 
.A(n_10696),
.B(n_363),
.C(n_364),
.Y(n_11042)
);

AOI21xp33_ASAP7_75t_L g11043 ( 
.A1(n_10689),
.A2(n_363),
.B(n_365),
.Y(n_11043)
);

NAND2x1_ASAP7_75t_L g11044 ( 
.A(n_10633),
.B(n_4594),
.Y(n_11044)
);

O2A1O1Ixp33_ASAP7_75t_L g11045 ( 
.A1(n_10608),
.A2(n_367),
.B(n_365),
.C(n_366),
.Y(n_11045)
);

BUFx2_ASAP7_75t_L g11046 ( 
.A(n_10426),
.Y(n_11046)
);

AOI21xp5_ASAP7_75t_L g11047 ( 
.A1(n_10733),
.A2(n_4597),
.B(n_4596),
.Y(n_11047)
);

BUFx4f_ASAP7_75t_L g11048 ( 
.A(n_10552),
.Y(n_11048)
);

NOR2xp33_ASAP7_75t_L g11049 ( 
.A(n_10225),
.B(n_4598),
.Y(n_11049)
);

NOR2xp33_ASAP7_75t_L g11050 ( 
.A(n_10437),
.B(n_4600),
.Y(n_11050)
);

INVx4_ASAP7_75t_L g11051 ( 
.A(n_10245),
.Y(n_11051)
);

AOI21xp5_ASAP7_75t_L g11052 ( 
.A1(n_10765),
.A2(n_4602),
.B(n_4601),
.Y(n_11052)
);

INVxp67_ASAP7_75t_L g11053 ( 
.A(n_10471),
.Y(n_11053)
);

INVx1_ASAP7_75t_L g11054 ( 
.A(n_10329),
.Y(n_11054)
);

INVx1_ASAP7_75t_L g11055 ( 
.A(n_10332),
.Y(n_11055)
);

OAI22xp5_ASAP7_75t_L g11056 ( 
.A1(n_10255),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_11056)
);

AOI21xp5_ASAP7_75t_L g11057 ( 
.A1(n_10769),
.A2(n_10787),
.B(n_10772),
.Y(n_11057)
);

INVx1_ASAP7_75t_L g11058 ( 
.A(n_10333),
.Y(n_11058)
);

INVx1_ASAP7_75t_L g11059 ( 
.A(n_10334),
.Y(n_11059)
);

HB1xp67_ASAP7_75t_L g11060 ( 
.A(n_10357),
.Y(n_11060)
);

BUFx3_ASAP7_75t_L g11061 ( 
.A(n_10636),
.Y(n_11061)
);

NAND2xp5_ASAP7_75t_L g11062 ( 
.A(n_10759),
.B(n_369),
.Y(n_11062)
);

AOI21xp5_ASAP7_75t_L g11063 ( 
.A1(n_10798),
.A2(n_4605),
.B(n_4603),
.Y(n_11063)
);

INVx2_ASAP7_75t_L g11064 ( 
.A(n_10750),
.Y(n_11064)
);

AOI21xp5_ASAP7_75t_L g11065 ( 
.A1(n_10807),
.A2(n_4607),
.B(n_4606),
.Y(n_11065)
);

AOI21xp5_ASAP7_75t_L g11066 ( 
.A1(n_10813),
.A2(n_4610),
.B(n_4608),
.Y(n_11066)
);

INVx1_ASAP7_75t_SL g11067 ( 
.A(n_10450),
.Y(n_11067)
);

INVx1_ASAP7_75t_L g11068 ( 
.A(n_10335),
.Y(n_11068)
);

NAND2xp5_ASAP7_75t_L g11069 ( 
.A(n_10761),
.B(n_369),
.Y(n_11069)
);

AOI21xp5_ASAP7_75t_L g11070 ( 
.A1(n_10637),
.A2(n_4615),
.B(n_4614),
.Y(n_11070)
);

NAND2xp5_ASAP7_75t_L g11071 ( 
.A(n_10764),
.B(n_370),
.Y(n_11071)
);

NAND2xp5_ASAP7_75t_L g11072 ( 
.A(n_10770),
.B(n_371),
.Y(n_11072)
);

INVx1_ASAP7_75t_L g11073 ( 
.A(n_10336),
.Y(n_11073)
);

NAND2xp5_ASAP7_75t_L g11074 ( 
.A(n_10771),
.B(n_372),
.Y(n_11074)
);

O2A1O1Ixp33_ASAP7_75t_L g11075 ( 
.A1(n_10620),
.A2(n_374),
.B(n_372),
.C(n_373),
.Y(n_11075)
);

AOI21xp5_ASAP7_75t_L g11076 ( 
.A1(n_10638),
.A2(n_10658),
.B(n_10655),
.Y(n_11076)
);

AOI21xp5_ASAP7_75t_L g11077 ( 
.A1(n_10439),
.A2(n_10667),
.B(n_10286),
.Y(n_11077)
);

AOI21xp5_ASAP7_75t_L g11078 ( 
.A1(n_10665),
.A2(n_4617),
.B(n_4616),
.Y(n_11078)
);

OR2x6_ASAP7_75t_L g11079 ( 
.A(n_10209),
.B(n_10218),
.Y(n_11079)
);

NAND2xp5_ASAP7_75t_L g11080 ( 
.A(n_10775),
.B(n_373),
.Y(n_11080)
);

OAI22xp5_ASAP7_75t_L g11081 ( 
.A1(n_10778),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_11081)
);

INVx2_ASAP7_75t_L g11082 ( 
.A(n_10751),
.Y(n_11082)
);

NAND2xp5_ASAP7_75t_L g11083 ( 
.A(n_10777),
.B(n_376),
.Y(n_11083)
);

NOR2xp67_ASAP7_75t_L g11084 ( 
.A(n_10697),
.B(n_4618),
.Y(n_11084)
);

AOI21xp5_ASAP7_75t_L g11085 ( 
.A1(n_10702),
.A2(n_4621),
.B(n_4620),
.Y(n_11085)
);

NOR2xp33_ASAP7_75t_L g11086 ( 
.A(n_10720),
.B(n_10749),
.Y(n_11086)
);

CKINVDCx5p33_ASAP7_75t_R g11087 ( 
.A(n_10781),
.Y(n_11087)
);

AOI21xp5_ASAP7_75t_L g11088 ( 
.A1(n_10705),
.A2(n_4623),
.B(n_4622),
.Y(n_11088)
);

OAI21xp5_ASAP7_75t_L g11089 ( 
.A1(n_10677),
.A2(n_377),
.B(n_378),
.Y(n_11089)
);

NAND2xp5_ASAP7_75t_SL g11090 ( 
.A(n_10600),
.B(n_4624),
.Y(n_11090)
);

NAND2xp5_ASAP7_75t_SL g11091 ( 
.A(n_10602),
.B(n_4625),
.Y(n_11091)
);

INVxp67_ASAP7_75t_SL g11092 ( 
.A(n_10755),
.Y(n_11092)
);

OAI22xp5_ASAP7_75t_L g11093 ( 
.A1(n_10783),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_11093)
);

OAI321xp33_ASAP7_75t_L g11094 ( 
.A1(n_10734),
.A2(n_381),
.A3(n_383),
.B1(n_379),
.B2(n_380),
.C(n_382),
.Y(n_11094)
);

AOI21xp5_ASAP7_75t_L g11095 ( 
.A1(n_10736),
.A2(n_10760),
.B(n_10259),
.Y(n_11095)
);

AOI21xp5_ASAP7_75t_L g11096 ( 
.A1(n_10673),
.A2(n_4627),
.B(n_4626),
.Y(n_11096)
);

AOI21x1_ASAP7_75t_L g11097 ( 
.A1(n_10657),
.A2(n_4629),
.B(n_4628),
.Y(n_11097)
);

NAND2xp5_ASAP7_75t_L g11098 ( 
.A(n_10799),
.B(n_380),
.Y(n_11098)
);

NOR2xp67_ASAP7_75t_L g11099 ( 
.A(n_10686),
.B(n_4630),
.Y(n_11099)
);

AOI21xp5_ASAP7_75t_L g11100 ( 
.A1(n_10683),
.A2(n_4632),
.B(n_4631),
.Y(n_11100)
);

AOI21xp5_ASAP7_75t_L g11101 ( 
.A1(n_10431),
.A2(n_4634),
.B(n_4633),
.Y(n_11101)
);

AOI22xp5_ASAP7_75t_L g11102 ( 
.A1(n_10607),
.A2(n_384),
.B1(n_381),
.B2(n_382),
.Y(n_11102)
);

AOI21xp5_ASAP7_75t_L g11103 ( 
.A1(n_10763),
.A2(n_4637),
.B(n_4635),
.Y(n_11103)
);

INVx1_ASAP7_75t_L g11104 ( 
.A(n_10340),
.Y(n_11104)
);

AOI21xp5_ASAP7_75t_L g11105 ( 
.A1(n_10298),
.A2(n_4639),
.B(n_4638),
.Y(n_11105)
);

AND2x2_ASAP7_75t_L g11106 ( 
.A(n_10553),
.B(n_4640),
.Y(n_11106)
);

INVx2_ASAP7_75t_L g11107 ( 
.A(n_10790),
.Y(n_11107)
);

INVx1_ASAP7_75t_L g11108 ( 
.A(n_10344),
.Y(n_11108)
);

AOI22x1_ASAP7_75t_L g11109 ( 
.A1(n_10282),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_11109)
);

BUFx3_ASAP7_75t_L g11110 ( 
.A(n_10544),
.Y(n_11110)
);

HB1xp67_ASAP7_75t_L g11111 ( 
.A(n_10345),
.Y(n_11111)
);

NOR2xp33_ASAP7_75t_L g11112 ( 
.A(n_10789),
.B(n_4643),
.Y(n_11112)
);

OAI21xp33_ASAP7_75t_L g11113 ( 
.A1(n_10331),
.A2(n_386),
.B(n_387),
.Y(n_11113)
);

INVx2_ASAP7_75t_L g11114 ( 
.A(n_10791),
.Y(n_11114)
);

NOR2xp33_ASAP7_75t_L g11115 ( 
.A(n_10794),
.B(n_10634),
.Y(n_11115)
);

NAND2xp5_ASAP7_75t_L g11116 ( 
.A(n_10438),
.B(n_387),
.Y(n_11116)
);

NOR2xp33_ASAP7_75t_L g11117 ( 
.A(n_10675),
.B(n_4644),
.Y(n_11117)
);

AOI21xp5_ASAP7_75t_L g11118 ( 
.A1(n_10403),
.A2(n_4646),
.B(n_4645),
.Y(n_11118)
);

AOI21x1_ASAP7_75t_L g11119 ( 
.A1(n_10575),
.A2(n_4650),
.B(n_4649),
.Y(n_11119)
);

AOI21xp5_ASAP7_75t_L g11120 ( 
.A1(n_10319),
.A2(n_4652),
.B(n_4651),
.Y(n_11120)
);

NAND2xp5_ASAP7_75t_L g11121 ( 
.A(n_10442),
.B(n_388),
.Y(n_11121)
);

O2A1O1Ixp5_ASAP7_75t_L g11122 ( 
.A1(n_10415),
.A2(n_390),
.B(n_388),
.C(n_389),
.Y(n_11122)
);

INVx1_ASAP7_75t_L g11123 ( 
.A(n_10352),
.Y(n_11123)
);

NAND2x1p5_ASAP7_75t_L g11124 ( 
.A(n_10285),
.B(n_4653),
.Y(n_11124)
);

NAND2xp5_ASAP7_75t_L g11125 ( 
.A(n_10453),
.B(n_389),
.Y(n_11125)
);

INVx2_ASAP7_75t_L g11126 ( 
.A(n_10293),
.Y(n_11126)
);

BUFx6f_ASAP7_75t_L g11127 ( 
.A(n_10669),
.Y(n_11127)
);

AOI21xp5_ASAP7_75t_L g11128 ( 
.A1(n_10630),
.A2(n_4657),
.B(n_4654),
.Y(n_11128)
);

AOI21xp5_ASAP7_75t_L g11129 ( 
.A1(n_10661),
.A2(n_4659),
.B(n_4658),
.Y(n_11129)
);

INVx2_ASAP7_75t_SL g11130 ( 
.A(n_10353),
.Y(n_11130)
);

NAND2xp5_ASAP7_75t_L g11131 ( 
.A(n_10454),
.B(n_390),
.Y(n_11131)
);

INVx1_ASAP7_75t_SL g11132 ( 
.A(n_10645),
.Y(n_11132)
);

INVx2_ASAP7_75t_L g11133 ( 
.A(n_10313),
.Y(n_11133)
);

BUFx6f_ASAP7_75t_L g11134 ( 
.A(n_10360),
.Y(n_11134)
);

NAND3xp33_ASAP7_75t_L g11135 ( 
.A(n_10574),
.B(n_391),
.C(n_392),
.Y(n_11135)
);

AOI21xp5_ASAP7_75t_L g11136 ( 
.A1(n_10436),
.A2(n_10262),
.B(n_10408),
.Y(n_11136)
);

O2A1O1Ixp33_ASAP7_75t_L g11137 ( 
.A1(n_10375),
.A2(n_393),
.B(n_391),
.C(n_392),
.Y(n_11137)
);

AOI21xp5_ASAP7_75t_L g11138 ( 
.A1(n_10322),
.A2(n_4661),
.B(n_4660),
.Y(n_11138)
);

OAI21xp5_ASAP7_75t_L g11139 ( 
.A1(n_10423),
.A2(n_393),
.B(n_394),
.Y(n_11139)
);

NAND2xp5_ASAP7_75t_L g11140 ( 
.A(n_10455),
.B(n_394),
.Y(n_11140)
);

OAI22xp5_ASAP7_75t_L g11141 ( 
.A1(n_10812),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_11141)
);

OAI21x1_ASAP7_75t_L g11142 ( 
.A1(n_10354),
.A2(n_4663),
.B(n_4662),
.Y(n_11142)
);

BUFx12f_ASAP7_75t_L g11143 ( 
.A(n_10487),
.Y(n_11143)
);

INVx2_ASAP7_75t_SL g11144 ( 
.A(n_10571),
.Y(n_11144)
);

NAND2xp5_ASAP7_75t_SL g11145 ( 
.A(n_10707),
.B(n_4664),
.Y(n_11145)
);

INVx2_ASAP7_75t_L g11146 ( 
.A(n_10348),
.Y(n_11146)
);

INVxp33_ASAP7_75t_SL g11147 ( 
.A(n_10461),
.Y(n_11147)
);

AOI21xp5_ASAP7_75t_L g11148 ( 
.A1(n_10622),
.A2(n_4668),
.B(n_4665),
.Y(n_11148)
);

INVx3_ASAP7_75t_L g11149 ( 
.A(n_10741),
.Y(n_11149)
);

AOI21xp5_ASAP7_75t_L g11150 ( 
.A1(n_10565),
.A2(n_4671),
.B(n_4670),
.Y(n_11150)
);

NOR2xp33_ASAP7_75t_L g11151 ( 
.A(n_10708),
.B(n_10711),
.Y(n_11151)
);

OAI22xp5_ASAP7_75t_L g11152 ( 
.A1(n_10427),
.A2(n_398),
.B1(n_395),
.B2(n_397),
.Y(n_11152)
);

NAND2xp5_ASAP7_75t_L g11153 ( 
.A(n_10456),
.B(n_10458),
.Y(n_11153)
);

INVx1_ASAP7_75t_L g11154 ( 
.A(n_10363),
.Y(n_11154)
);

INVx2_ASAP7_75t_L g11155 ( 
.A(n_10349),
.Y(n_11155)
);

BUFx3_ASAP7_75t_L g11156 ( 
.A(n_10726),
.Y(n_11156)
);

OA22x2_ASAP7_75t_L g11157 ( 
.A1(n_10418),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_11157)
);

AOI21xp5_ASAP7_75t_L g11158 ( 
.A1(n_10238),
.A2(n_4673),
.B(n_4672),
.Y(n_11158)
);

AOI21xp5_ASAP7_75t_L g11159 ( 
.A1(n_10406),
.A2(n_4675),
.B(n_4674),
.Y(n_11159)
);

AOI21xp5_ASAP7_75t_L g11160 ( 
.A1(n_10409),
.A2(n_4678),
.B(n_4677),
.Y(n_11160)
);

INVx2_ASAP7_75t_L g11161 ( 
.A(n_10355),
.Y(n_11161)
);

NAND2xp5_ASAP7_75t_L g11162 ( 
.A(n_10462),
.B(n_399),
.Y(n_11162)
);

INVx1_ASAP7_75t_L g11163 ( 
.A(n_10364),
.Y(n_11163)
);

NAND2xp5_ASAP7_75t_L g11164 ( 
.A(n_10388),
.B(n_401),
.Y(n_11164)
);

NAND2xp5_ASAP7_75t_L g11165 ( 
.A(n_10213),
.B(n_401),
.Y(n_11165)
);

NOR3xp33_ASAP7_75t_L g11166 ( 
.A(n_10666),
.B(n_402),
.C(n_403),
.Y(n_11166)
);

AO21x1_ASAP7_75t_L g11167 ( 
.A1(n_10448),
.A2(n_402),
.B(n_403),
.Y(n_11167)
);

INVx1_ASAP7_75t_L g11168 ( 
.A(n_10367),
.Y(n_11168)
);

A2O1A1Ixp33_ASAP7_75t_L g11169 ( 
.A1(n_10470),
.A2(n_406),
.B(n_404),
.C(n_405),
.Y(n_11169)
);

NAND2xp5_ASAP7_75t_L g11170 ( 
.A(n_10216),
.B(n_406),
.Y(n_11170)
);

NAND2xp5_ASAP7_75t_L g11171 ( 
.A(n_10224),
.B(n_407),
.Y(n_11171)
);

AOI21xp5_ASAP7_75t_L g11172 ( 
.A1(n_10474),
.A2(n_4680),
.B(n_4679),
.Y(n_11172)
);

OAI21xp5_ASAP7_75t_L g11173 ( 
.A1(n_10502),
.A2(n_407),
.B(n_408),
.Y(n_11173)
);

OAI21xp5_ASAP7_75t_L g11174 ( 
.A1(n_10509),
.A2(n_408),
.B(n_409),
.Y(n_11174)
);

OAI22xp5_ASAP7_75t_L g11175 ( 
.A1(n_10688),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_11175)
);

NAND2xp5_ASAP7_75t_L g11176 ( 
.A(n_10228),
.B(n_410),
.Y(n_11176)
);

A2O1A1Ixp33_ASAP7_75t_L g11177 ( 
.A1(n_10512),
.A2(n_413),
.B(n_411),
.C(n_412),
.Y(n_11177)
);

NAND2xp5_ASAP7_75t_L g11178 ( 
.A(n_10230),
.B(n_413),
.Y(n_11178)
);

A2O1A1Ixp33_ASAP7_75t_L g11179 ( 
.A1(n_10396),
.A2(n_416),
.B(n_414),
.C(n_415),
.Y(n_11179)
);

NAND2xp5_ASAP7_75t_L g11180 ( 
.A(n_10231),
.B(n_415),
.Y(n_11180)
);

AOI21xp5_ASAP7_75t_L g11181 ( 
.A1(n_10767),
.A2(n_4683),
.B(n_4682),
.Y(n_11181)
);

NAND2xp5_ASAP7_75t_L g11182 ( 
.A(n_10234),
.B(n_416),
.Y(n_11182)
);

NAND2xp5_ASAP7_75t_L g11183 ( 
.A(n_10236),
.B(n_417),
.Y(n_11183)
);

AOI21x1_ASAP7_75t_L g11184 ( 
.A1(n_10576),
.A2(n_4685),
.B(n_4684),
.Y(n_11184)
);

OAI22xp5_ASAP7_75t_L g11185 ( 
.A1(n_10672),
.A2(n_419),
.B1(n_417),
.B2(n_418),
.Y(n_11185)
);

HB1xp67_ASAP7_75t_L g11186 ( 
.A(n_10368),
.Y(n_11186)
);

AOI21xp5_ASAP7_75t_L g11187 ( 
.A1(n_10237),
.A2(n_4688),
.B(n_4687),
.Y(n_11187)
);

NAND2xp5_ASAP7_75t_SL g11188 ( 
.A(n_10681),
.B(n_4689),
.Y(n_11188)
);

INVx1_ASAP7_75t_L g11189 ( 
.A(n_10370),
.Y(n_11189)
);

A2O1A1Ixp33_ASAP7_75t_L g11190 ( 
.A1(n_10640),
.A2(n_420),
.B(n_418),
.C(n_419),
.Y(n_11190)
);

AOI22xp33_ASAP7_75t_L g11191 ( 
.A1(n_10214),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_11191)
);

AOI21xp5_ASAP7_75t_L g11192 ( 
.A1(n_10240),
.A2(n_4691),
.B(n_4690),
.Y(n_11192)
);

OAI21xp5_ASAP7_75t_L g11193 ( 
.A1(n_10671),
.A2(n_421),
.B(n_422),
.Y(n_11193)
);

AOI21xp5_ASAP7_75t_L g11194 ( 
.A1(n_10243),
.A2(n_4693),
.B(n_4692),
.Y(n_11194)
);

AOI21xp5_ASAP7_75t_L g11195 ( 
.A1(n_10244),
.A2(n_4695),
.B(n_4694),
.Y(n_11195)
);

INVx3_ASAP7_75t_L g11196 ( 
.A(n_10748),
.Y(n_11196)
);

OAI321xp33_ASAP7_75t_L g11197 ( 
.A1(n_10817),
.A2(n_425),
.A3(n_427),
.B1(n_423),
.B2(n_424),
.C(n_426),
.Y(n_11197)
);

O2A1O1Ixp33_ASAP7_75t_L g11198 ( 
.A1(n_10631),
.A2(n_10586),
.B(n_10381),
.C(n_10445),
.Y(n_11198)
);

NOR2xp33_ASAP7_75t_L g11199 ( 
.A(n_10756),
.B(n_4696),
.Y(n_11199)
);

AOI21xp5_ASAP7_75t_L g11200 ( 
.A1(n_10248),
.A2(n_4698),
.B(n_4697),
.Y(n_11200)
);

INVx2_ASAP7_75t_L g11201 ( 
.A(n_10404),
.Y(n_11201)
);

AO32x1_ASAP7_75t_L g11202 ( 
.A1(n_10611),
.A2(n_426),
.A3(n_424),
.B1(n_425),
.B2(n_427),
.Y(n_11202)
);

AOI22xp5_ASAP7_75t_L g11203 ( 
.A1(n_10805),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.Y(n_11203)
);

AOI21xp5_ASAP7_75t_L g11204 ( 
.A1(n_10251),
.A2(n_4701),
.B(n_4699),
.Y(n_11204)
);

AND2x2_ASAP7_75t_L g11205 ( 
.A(n_10390),
.B(n_4703),
.Y(n_11205)
);

BUFx12f_ASAP7_75t_L g11206 ( 
.A(n_10504),
.Y(n_11206)
);

A2O1A1Ixp33_ASAP7_75t_L g11207 ( 
.A1(n_10610),
.A2(n_430),
.B(n_428),
.C(n_429),
.Y(n_11207)
);

AND2x2_ASAP7_75t_L g11208 ( 
.A(n_10716),
.B(n_4704),
.Y(n_11208)
);

OAI21xp5_ASAP7_75t_L g11209 ( 
.A1(n_10643),
.A2(n_431),
.B(n_432),
.Y(n_11209)
);

OR2x2_ASAP7_75t_L g11210 ( 
.A(n_10297),
.B(n_431),
.Y(n_11210)
);

INVx8_ASAP7_75t_L g11211 ( 
.A(n_10296),
.Y(n_11211)
);

AOI21xp5_ASAP7_75t_L g11212 ( 
.A1(n_10260),
.A2(n_4706),
.B(n_4705),
.Y(n_11212)
);

OAI21xp5_ASAP7_75t_L g11213 ( 
.A1(n_10314),
.A2(n_432),
.B(n_434),
.Y(n_11213)
);

BUFx12f_ASAP7_75t_L g11214 ( 
.A(n_10342),
.Y(n_11214)
);

NAND2xp5_ASAP7_75t_SL g11215 ( 
.A(n_10682),
.B(n_4707),
.Y(n_11215)
);

INVx2_ASAP7_75t_L g11216 ( 
.A(n_10424),
.Y(n_11216)
);

O2A1O1Ixp33_ASAP7_75t_L g11217 ( 
.A1(n_10641),
.A2(n_10727),
.B(n_10518),
.C(n_10524),
.Y(n_11217)
);

AOI21x1_ASAP7_75t_L g11218 ( 
.A1(n_10371),
.A2(n_4709),
.B(n_4708),
.Y(n_11218)
);

NAND2xp5_ASAP7_75t_L g11219 ( 
.A(n_10264),
.B(n_434),
.Y(n_11219)
);

AOI21xp5_ASAP7_75t_L g11220 ( 
.A1(n_10268),
.A2(n_4712),
.B(n_4711),
.Y(n_11220)
);

NAND2xp5_ASAP7_75t_L g11221 ( 
.A(n_10269),
.B(n_10270),
.Y(n_11221)
);

O2A1O1Ixp5_ASAP7_75t_L g11222 ( 
.A1(n_10687),
.A2(n_437),
.B(n_435),
.C(n_436),
.Y(n_11222)
);

NAND2xp5_ASAP7_75t_L g11223 ( 
.A(n_10273),
.B(n_435),
.Y(n_11223)
);

A2O1A1Ixp33_ASAP7_75t_L g11224 ( 
.A1(n_10488),
.A2(n_439),
.B(n_436),
.C(n_438),
.Y(n_11224)
);

AOI21xp5_ASAP7_75t_L g11225 ( 
.A1(n_10289),
.A2(n_4715),
.B(n_4713),
.Y(n_11225)
);

AND2x2_ASAP7_75t_L g11226 ( 
.A(n_10222),
.B(n_4716),
.Y(n_11226)
);

NAND2xp5_ASAP7_75t_L g11227 ( 
.A(n_10425),
.B(n_438),
.Y(n_11227)
);

OAI22xp5_ASAP7_75t_L g11228 ( 
.A1(n_10628),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_11228)
);

AOI21xp5_ASAP7_75t_L g11229 ( 
.A1(n_10706),
.A2(n_4719),
.B(n_4717),
.Y(n_11229)
);

INVx1_ASAP7_75t_L g11230 ( 
.A(n_10372),
.Y(n_11230)
);

AO21x1_ASAP7_75t_L g11231 ( 
.A1(n_10684),
.A2(n_440),
.B(n_441),
.Y(n_11231)
);

AOI21xp5_ASAP7_75t_L g11232 ( 
.A1(n_10595),
.A2(n_4721),
.B(n_4720),
.Y(n_11232)
);

NOR2x1p5_ASAP7_75t_SL g11233 ( 
.A(n_10440),
.B(n_4722),
.Y(n_11233)
);

NAND2xp5_ASAP7_75t_L g11234 ( 
.A(n_10444),
.B(n_442),
.Y(n_11234)
);

OAI21xp33_ASAP7_75t_L g11235 ( 
.A1(n_10302),
.A2(n_10327),
.B(n_10233),
.Y(n_11235)
);

NAND2xp5_ASAP7_75t_L g11236 ( 
.A(n_10401),
.B(n_443),
.Y(n_11236)
);

INVx2_ASAP7_75t_L g11237 ( 
.A(n_10402),
.Y(n_11237)
);

O2A1O1Ixp33_ASAP7_75t_L g11238 ( 
.A1(n_10583),
.A2(n_445),
.B(n_443),
.C(n_444),
.Y(n_11238)
);

NAND2xp5_ASAP7_75t_L g11239 ( 
.A(n_10407),
.B(n_445),
.Y(n_11239)
);

BUFx6f_ASAP7_75t_L g11240 ( 
.A(n_10361),
.Y(n_11240)
);

OR2x6_ASAP7_75t_L g11241 ( 
.A(n_10209),
.B(n_4723),
.Y(n_11241)
);

NOR2xp33_ASAP7_75t_L g11242 ( 
.A(n_10780),
.B(n_4725),
.Y(n_11242)
);

NOR2xp33_ASAP7_75t_SL g11243 ( 
.A(n_10486),
.B(n_4726),
.Y(n_11243)
);

AOI21xp33_ASAP7_75t_L g11244 ( 
.A1(n_10670),
.A2(n_446),
.B(n_447),
.Y(n_11244)
);

INVxp67_ASAP7_75t_SL g11245 ( 
.A(n_10410),
.Y(n_11245)
);

HB1xp67_ASAP7_75t_L g11246 ( 
.A(n_10373),
.Y(n_11246)
);

INVx2_ASAP7_75t_L g11247 ( 
.A(n_10413),
.Y(n_11247)
);

AND2x2_ASAP7_75t_L g11248 ( 
.A(n_10309),
.B(n_4727),
.Y(n_11248)
);

NAND2xp5_ASAP7_75t_SL g11249 ( 
.A(n_10625),
.B(n_4728),
.Y(n_11249)
);

NAND2xp5_ASAP7_75t_L g11250 ( 
.A(n_10414),
.B(n_446),
.Y(n_11250)
);

A2O1A1Ixp33_ASAP7_75t_L g11251 ( 
.A1(n_10419),
.A2(n_449),
.B(n_447),
.C(n_448),
.Y(n_11251)
);

INVx1_ASAP7_75t_L g11252 ( 
.A(n_10376),
.Y(n_11252)
);

NAND2xp5_ASAP7_75t_L g11253 ( 
.A(n_10421),
.B(n_448),
.Y(n_11253)
);

NAND2xp5_ASAP7_75t_L g11254 ( 
.A(n_10428),
.B(n_450),
.Y(n_11254)
);

NAND2xp5_ASAP7_75t_L g11255 ( 
.A(n_10482),
.B(n_10377),
.Y(n_11255)
);

INVx1_ASAP7_75t_L g11256 ( 
.A(n_10383),
.Y(n_11256)
);

AOI21xp5_ASAP7_75t_L g11257 ( 
.A1(n_10275),
.A2(n_4731),
.B(n_4730),
.Y(n_11257)
);

NAND2xp5_ASAP7_75t_L g11258 ( 
.A(n_10384),
.B(n_450),
.Y(n_11258)
);

INVx2_ASAP7_75t_L g11259 ( 
.A(n_10597),
.Y(n_11259)
);

AOI21xp5_ASAP7_75t_L g11260 ( 
.A1(n_10303),
.A2(n_4733),
.B(n_4732),
.Y(n_11260)
);

INVx1_ASAP7_75t_L g11261 ( 
.A(n_10616),
.Y(n_11261)
);

AOI21x1_ASAP7_75t_L g11262 ( 
.A1(n_10304),
.A2(n_4735),
.B(n_4734),
.Y(n_11262)
);

INVxp67_ASAP7_75t_L g11263 ( 
.A(n_10629),
.Y(n_11263)
);

AOI22xp5_ASAP7_75t_L g11264 ( 
.A1(n_10805),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_11264)
);

INVx3_ASAP7_75t_L g11265 ( 
.A(n_10584),
.Y(n_11265)
);

INVx2_ASAP7_75t_L g11266 ( 
.A(n_10619),
.Y(n_11266)
);

NAND2xp5_ASAP7_75t_L g11267 ( 
.A(n_10530),
.B(n_452),
.Y(n_11267)
);

NAND2xp5_ASAP7_75t_L g11268 ( 
.A(n_10432),
.B(n_453),
.Y(n_11268)
);

NAND2x1p5_ASAP7_75t_L g11269 ( 
.A(n_10385),
.B(n_4736),
.Y(n_11269)
);

NAND3xp33_ASAP7_75t_L g11270 ( 
.A(n_10592),
.B(n_454),
.C(n_455),
.Y(n_11270)
);

INVx1_ASAP7_75t_L g11271 ( 
.A(n_10493),
.Y(n_11271)
);

AOI21xp5_ASAP7_75t_L g11272 ( 
.A1(n_10374),
.A2(n_4739),
.B(n_4737),
.Y(n_11272)
);

INVx1_ASAP7_75t_L g11273 ( 
.A(n_10499),
.Y(n_11273)
);

A2O1A1Ixp33_ASAP7_75t_L g11274 ( 
.A1(n_10369),
.A2(n_456),
.B(n_454),
.C(n_455),
.Y(n_11274)
);

AOI21xp5_ASAP7_75t_L g11275 ( 
.A1(n_10379),
.A2(n_4741),
.B(n_4740),
.Y(n_11275)
);

NAND2xp5_ASAP7_75t_L g11276 ( 
.A(n_10239),
.B(n_457),
.Y(n_11276)
);

AOI21xp5_ASAP7_75t_L g11277 ( 
.A1(n_10429),
.A2(n_4743),
.B(n_4742),
.Y(n_11277)
);

AND2x2_ASAP7_75t_L g11278 ( 
.A(n_10395),
.B(n_4744),
.Y(n_11278)
);

NAND2xp5_ASAP7_75t_SL g11279 ( 
.A(n_10662),
.B(n_4747),
.Y(n_11279)
);

NAND2xp5_ASAP7_75t_L g11280 ( 
.A(n_10246),
.B(n_458),
.Y(n_11280)
);

AOI22xp33_ASAP7_75t_L g11281 ( 
.A1(n_10496),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_11281)
);

NAND2xp5_ASAP7_75t_L g11282 ( 
.A(n_10700),
.B(n_459),
.Y(n_11282)
);

AOI22x1_ASAP7_75t_L g11283 ( 
.A1(n_10330),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_11283)
);

NAND2xp5_ASAP7_75t_L g11284 ( 
.A(n_10593),
.B(n_10494),
.Y(n_11284)
);

INVx4_ASAP7_75t_L g11285 ( 
.A(n_10429),
.Y(n_11285)
);

NAND2xp5_ASAP7_75t_SL g11286 ( 
.A(n_10680),
.B(n_4748),
.Y(n_11286)
);

INVx2_ASAP7_75t_L g11287 ( 
.A(n_10272),
.Y(n_11287)
);

AOI21xp5_ASAP7_75t_L g11288 ( 
.A1(n_10261),
.A2(n_4751),
.B(n_4750),
.Y(n_11288)
);

AOI22xp33_ASAP7_75t_L g11289 ( 
.A1(n_10265),
.A2(n_464),
.B1(n_461),
.B2(n_463),
.Y(n_11289)
);

O2A1O1Ixp33_ASAP7_75t_L g11290 ( 
.A1(n_10389),
.A2(n_466),
.B(n_464),
.C(n_465),
.Y(n_11290)
);

AOI21xp5_ASAP7_75t_L g11291 ( 
.A1(n_10635),
.A2(n_4753),
.B(n_4752),
.Y(n_11291)
);

OAI22xp5_ASAP7_75t_L g11292 ( 
.A1(n_10642),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_11292)
);

NOR2xp33_ASAP7_75t_L g11293 ( 
.A(n_10649),
.B(n_4754),
.Y(n_11293)
);

AOI21xp5_ASAP7_75t_L g11294 ( 
.A1(n_10362),
.A2(n_4758),
.B(n_4757),
.Y(n_11294)
);

NOR2xp67_ASAP7_75t_L g11295 ( 
.A(n_10810),
.B(n_4759),
.Y(n_11295)
);

OAI22xp5_ASAP7_75t_L g11296 ( 
.A1(n_10668),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_11296)
);

NOR2xp33_ASAP7_75t_L g11297 ( 
.A(n_10663),
.B(n_4760),
.Y(n_11297)
);

AND2x2_ASAP7_75t_L g11298 ( 
.A(n_10434),
.B(n_4761),
.Y(n_11298)
);

OAI22xp5_ASAP7_75t_L g11299 ( 
.A1(n_10547),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.Y(n_11299)
);

AOI21xp5_ASAP7_75t_L g11300 ( 
.A1(n_10387),
.A2(n_4763),
.B(n_4762),
.Y(n_11300)
);

BUFx2_ASAP7_75t_L g11301 ( 
.A(n_10606),
.Y(n_11301)
);

AOI21xp5_ASAP7_75t_L g11302 ( 
.A1(n_10490),
.A2(n_4765),
.B(n_4764),
.Y(n_11302)
);

AOI21xp5_ASAP7_75t_L g11303 ( 
.A1(n_10549),
.A2(n_4767),
.B(n_4766),
.Y(n_11303)
);

AOI21xp5_ASAP7_75t_L g11304 ( 
.A1(n_10218),
.A2(n_4770),
.B(n_4768),
.Y(n_11304)
);

NAND2xp5_ASAP7_75t_L g11305 ( 
.A(n_10420),
.B(n_470),
.Y(n_11305)
);

HB1xp67_ASAP7_75t_L g11306 ( 
.A(n_10516),
.Y(n_11306)
);

AND2x2_ASAP7_75t_L g11307 ( 
.A(n_10498),
.B(n_4775),
.Y(n_11307)
);

NAND2xp5_ASAP7_75t_L g11308 ( 
.A(n_10447),
.B(n_471),
.Y(n_11308)
);

NOR2xp33_ASAP7_75t_L g11309 ( 
.A(n_10441),
.B(n_4776),
.Y(n_11309)
);

BUFx4f_ASAP7_75t_L g11310 ( 
.A(n_10266),
.Y(n_11310)
);

AOI21xp5_ASAP7_75t_L g11311 ( 
.A1(n_10266),
.A2(n_4778),
.B(n_4777),
.Y(n_11311)
);

OAI22xp5_ASAP7_75t_L g11312 ( 
.A1(n_10647),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_11312)
);

OAI21xp33_ASAP7_75t_L g11313 ( 
.A1(n_10479),
.A2(n_472),
.B(n_473),
.Y(n_11313)
);

AOI22xp5_ASAP7_75t_L g11314 ( 
.A1(n_10523),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.Y(n_11314)
);

AOI21xp5_ASAP7_75t_L g11315 ( 
.A1(n_10284),
.A2(n_4780),
.B(n_4779),
.Y(n_11315)
);

O2A1O1Ixp33_ASAP7_75t_L g11316 ( 
.A1(n_10646),
.A2(n_477),
.B(n_475),
.C(n_476),
.Y(n_11316)
);

INVx1_ASAP7_75t_L g11317 ( 
.A(n_10320),
.Y(n_11317)
);

INVx5_ASAP7_75t_L g11318 ( 
.A(n_10652),
.Y(n_11318)
);

INVx1_ASAP7_75t_L g11319 ( 
.A(n_10475),
.Y(n_11319)
);

INVx4_ASAP7_75t_L g11320 ( 
.A(n_10393),
.Y(n_11320)
);

AOI21xp5_ASAP7_75t_L g11321 ( 
.A1(n_10292),
.A2(n_4782),
.B(n_4781),
.Y(n_11321)
);

AOI21x1_ASAP7_75t_L g11322 ( 
.A1(n_10459),
.A2(n_4785),
.B(n_4783),
.Y(n_11322)
);

BUFx8_ASAP7_75t_L g11323 ( 
.A(n_10578),
.Y(n_11323)
);

NAND2xp5_ASAP7_75t_L g11324 ( 
.A(n_10618),
.B(n_477),
.Y(n_11324)
);

NAND2x1_ASAP7_75t_L g11325 ( 
.A(n_10312),
.B(n_4786),
.Y(n_11325)
);

INVx3_ASAP7_75t_L g11326 ( 
.A(n_10416),
.Y(n_11326)
);

AOI21xp5_ASAP7_75t_L g11327 ( 
.A1(n_10693),
.A2(n_4790),
.B(n_4789),
.Y(n_11327)
);

O2A1O1Ixp33_ASAP7_75t_L g11328 ( 
.A1(n_10589),
.A2(n_480),
.B(n_478),
.C(n_479),
.Y(n_11328)
);

AOI21xp5_ASAP7_75t_L g11329 ( 
.A1(n_10704),
.A2(n_4792),
.B(n_4791),
.Y(n_11329)
);

AOI21x1_ASAP7_75t_L g11330 ( 
.A1(n_10338),
.A2(n_10358),
.B(n_10478),
.Y(n_11330)
);

NAND3xp33_ASAP7_75t_L g11331 ( 
.A(n_10526),
.B(n_478),
.C(n_479),
.Y(n_11331)
);

O2A1O1Ixp33_ASAP7_75t_L g11332 ( 
.A1(n_10527),
.A2(n_482),
.B(n_480),
.C(n_481),
.Y(n_11332)
);

NAND2xp5_ASAP7_75t_L g11333 ( 
.A(n_10443),
.B(n_481),
.Y(n_11333)
);

INVx1_ASAP7_75t_L g11334 ( 
.A(n_10534),
.Y(n_11334)
);

NAND2xp5_ASAP7_75t_L g11335 ( 
.A(n_10609),
.B(n_483),
.Y(n_11335)
);

BUFx6f_ASAP7_75t_L g11336 ( 
.A(n_10235),
.Y(n_11336)
);

AOI21xp5_ASAP7_75t_L g11337 ( 
.A1(n_10397),
.A2(n_4794),
.B(n_4793),
.Y(n_11337)
);

AND2x2_ASAP7_75t_L g11338 ( 
.A(n_10563),
.B(n_4795),
.Y(n_11338)
);

NOR2x1_ASAP7_75t_L g11339 ( 
.A(n_10564),
.B(n_483),
.Y(n_11339)
);

AOI21xp5_ASAP7_75t_L g11340 ( 
.A1(n_10422),
.A2(n_4799),
.B(n_4796),
.Y(n_11340)
);

NAND2xp5_ASAP7_75t_L g11341 ( 
.A(n_10605),
.B(n_10449),
.Y(n_11341)
);

BUFx2_ASAP7_75t_L g11342 ( 
.A(n_10247),
.Y(n_11342)
);

OAI321xp33_ASAP7_75t_L g11343 ( 
.A1(n_10399),
.A2(n_486),
.A3(n_488),
.B1(n_484),
.B2(n_485),
.C(n_487),
.Y(n_11343)
);

O2A1O1Ixp33_ASAP7_75t_L g11344 ( 
.A1(n_10632),
.A2(n_488),
.B(n_484),
.C(n_486),
.Y(n_11344)
);

NAND2xp5_ASAP7_75t_L g11345 ( 
.A(n_10678),
.B(n_489),
.Y(n_11345)
);

INVxp67_ASAP7_75t_L g11346 ( 
.A(n_10328),
.Y(n_11346)
);

AOI22xp33_ASAP7_75t_L g11347 ( 
.A1(n_10591),
.A2(n_10599),
.B1(n_10601),
.B2(n_10613),
.Y(n_11347)
);

BUFx6f_ASAP7_75t_L g11348 ( 
.A(n_10252),
.Y(n_11348)
);

NAND2xp5_ASAP7_75t_L g11349 ( 
.A(n_10614),
.B(n_489),
.Y(n_11349)
);

AOI21xp5_ASAP7_75t_L g11350 ( 
.A1(n_10480),
.A2(n_4802),
.B(n_4801),
.Y(n_11350)
);

OAI21xp5_ASAP7_75t_L g11351 ( 
.A1(n_10489),
.A2(n_490),
.B(n_491),
.Y(n_11351)
);

NOR2xp33_ASAP7_75t_L g11352 ( 
.A(n_10691),
.B(n_4804),
.Y(n_11352)
);

A2O1A1Ixp33_ASAP7_75t_L g11353 ( 
.A1(n_10263),
.A2(n_493),
.B(n_491),
.C(n_492),
.Y(n_11353)
);

OAI22xp5_ASAP7_75t_L g11354 ( 
.A1(n_10562),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_11354)
);

O2A1O1Ixp33_ASAP7_75t_L g11355 ( 
.A1(n_10219),
.A2(n_497),
.B(n_495),
.C(n_496),
.Y(n_11355)
);

INVx2_ASAP7_75t_L g11356 ( 
.A(n_10572),
.Y(n_11356)
);

NOR2xp33_ASAP7_75t_L g11357 ( 
.A(n_10250),
.B(n_4805),
.Y(n_11357)
);

NAND2x1_ASAP7_75t_L g11358 ( 
.A(n_10747),
.B(n_4806),
.Y(n_11358)
);

O2A1O1Ixp33_ASAP7_75t_L g11359 ( 
.A1(n_10725),
.A2(n_497),
.B(n_495),
.C(n_496),
.Y(n_11359)
);

NAND2xp5_ASAP7_75t_L g11360 ( 
.A(n_10617),
.B(n_498),
.Y(n_11360)
);

AOI21x1_ASAP7_75t_L g11361 ( 
.A1(n_10546),
.A2(n_4809),
.B(n_4808),
.Y(n_11361)
);

OAI21xp5_ASAP7_75t_L g11362 ( 
.A1(n_10737),
.A2(n_499),
.B(n_500),
.Y(n_11362)
);

INVx1_ASAP7_75t_L g11363 ( 
.A(n_10548),
.Y(n_11363)
);

AOI21xp5_ASAP7_75t_L g11364 ( 
.A1(n_10491),
.A2(n_4812),
.B(n_4811),
.Y(n_11364)
);

OAI22xp5_ASAP7_75t_L g11365 ( 
.A1(n_10627),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.Y(n_11365)
);

AOI21xp5_ASAP7_75t_L g11366 ( 
.A1(n_10508),
.A2(n_4815),
.B(n_4813),
.Y(n_11366)
);

NAND2xp5_ASAP7_75t_L g11367 ( 
.A(n_10639),
.B(n_501),
.Y(n_11367)
);

INVx3_ASAP7_75t_L g11368 ( 
.A(n_10762),
.Y(n_11368)
);

AND2x2_ASAP7_75t_SL g11369 ( 
.A(n_10776),
.B(n_502),
.Y(n_11369)
);

INVx1_ASAP7_75t_L g11370 ( 
.A(n_10580),
.Y(n_11370)
);

O2A1O1Ixp33_ASAP7_75t_L g11371 ( 
.A1(n_10809),
.A2(n_505),
.B(n_503),
.C(n_504),
.Y(n_11371)
);

A2O1A1Ixp33_ASAP7_75t_L g11372 ( 
.A1(n_10651),
.A2(n_506),
.B(n_503),
.C(n_505),
.Y(n_11372)
);

AO21x1_ASAP7_75t_L g11373 ( 
.A1(n_10582),
.A2(n_506),
.B(n_507),
.Y(n_11373)
);

AOI21xp5_ASAP7_75t_L g11374 ( 
.A1(n_10519),
.A2(n_10539),
.B(n_10522),
.Y(n_11374)
);

AOI21xp5_ASAP7_75t_L g11375 ( 
.A1(n_10542),
.A2(n_4817),
.B(n_4816),
.Y(n_11375)
);

INVxp67_ASAP7_75t_SL g11376 ( 
.A(n_10712),
.Y(n_11376)
);

AOI21xp5_ASAP7_75t_L g11377 ( 
.A1(n_10654),
.A2(n_10692),
.B(n_10685),
.Y(n_11377)
);

NAND2xp5_ASAP7_75t_L g11378 ( 
.A(n_10715),
.B(n_507),
.Y(n_11378)
);

NOR2xp33_ASAP7_75t_L g11379 ( 
.A(n_10804),
.B(n_4818),
.Y(n_11379)
);

A2O1A1Ixp33_ASAP7_75t_L g11380 ( 
.A1(n_10276),
.A2(n_510),
.B(n_508),
.C(n_509),
.Y(n_11380)
);

OAI22xp5_ASAP7_75t_L g11381 ( 
.A1(n_10276),
.A2(n_512),
.B1(n_508),
.B2(n_511),
.Y(n_11381)
);

AOI21xp5_ASAP7_75t_L g11382 ( 
.A1(n_10324),
.A2(n_4821),
.B(n_4820),
.Y(n_11382)
);

AND2x2_ASAP7_75t_SL g11383 ( 
.A(n_10308),
.B(n_511),
.Y(n_11383)
);

NAND2xp5_ASAP7_75t_L g11384 ( 
.A(n_10229),
.B(n_513),
.Y(n_11384)
);

NOR2xp33_ASAP7_75t_L g11385 ( 
.A(n_10276),
.B(n_4822),
.Y(n_11385)
);

NOR2xp33_ASAP7_75t_SL g11386 ( 
.A(n_10717),
.B(n_4824),
.Y(n_11386)
);

AND2x2_ASAP7_75t_L g11387 ( 
.A(n_10310),
.B(n_4825),
.Y(n_11387)
);

OAI22xp5_ASAP7_75t_L g11388 ( 
.A1(n_10276),
.A2(n_515),
.B1(n_513),
.B2(n_514),
.Y(n_11388)
);

INVx1_ASAP7_75t_SL g11389 ( 
.A(n_10215),
.Y(n_11389)
);

AND2x4_ASAP7_75t_L g11390 ( 
.A(n_10380),
.B(n_4826),
.Y(n_11390)
);

NOR2xp33_ASAP7_75t_L g11391 ( 
.A(n_10276),
.B(n_4827),
.Y(n_11391)
);

NOR2xp33_ASAP7_75t_L g11392 ( 
.A(n_10276),
.B(n_4828),
.Y(n_11392)
);

AOI21xp5_ASAP7_75t_L g11393 ( 
.A1(n_10324),
.A2(n_4831),
.B(n_4830),
.Y(n_11393)
);

NOR2xp33_ASAP7_75t_L g11394 ( 
.A(n_10276),
.B(n_4832),
.Y(n_11394)
);

OAI22xp5_ASAP7_75t_L g11395 ( 
.A1(n_10276),
.A2(n_516),
.B1(n_514),
.B2(n_515),
.Y(n_11395)
);

OAI21xp5_ASAP7_75t_L g11396 ( 
.A1(n_10276),
.A2(n_516),
.B(n_517),
.Y(n_11396)
);

INVxp67_ASAP7_75t_L g11397 ( 
.A(n_10217),
.Y(n_11397)
);

BUFx6f_ASAP7_75t_L g11398 ( 
.A(n_10318),
.Y(n_11398)
);

NOR2xp33_ASAP7_75t_L g11399 ( 
.A(n_10276),
.B(n_4834),
.Y(n_11399)
);

NOR2xp33_ASAP7_75t_L g11400 ( 
.A(n_10276),
.B(n_4835),
.Y(n_11400)
);

AOI22xp5_ASAP7_75t_L g11401 ( 
.A1(n_10276),
.A2(n_519),
.B1(n_517),
.B2(n_518),
.Y(n_11401)
);

AOI21xp5_ASAP7_75t_L g11402 ( 
.A1(n_10324),
.A2(n_4837),
.B(n_4836),
.Y(n_11402)
);

AOI21xp5_ASAP7_75t_L g11403 ( 
.A1(n_10324),
.A2(n_4840),
.B(n_4839),
.Y(n_11403)
);

AOI21xp5_ASAP7_75t_L g11404 ( 
.A1(n_10324),
.A2(n_4842),
.B(n_4841),
.Y(n_11404)
);

NAND2xp5_ASAP7_75t_L g11405 ( 
.A(n_10229),
.B(n_519),
.Y(n_11405)
);

INVx3_ASAP7_75t_L g11406 ( 
.A(n_10227),
.Y(n_11406)
);

NAND2xp5_ASAP7_75t_L g11407 ( 
.A(n_10229),
.B(n_520),
.Y(n_11407)
);

NAND2xp5_ASAP7_75t_SL g11408 ( 
.A(n_10229),
.B(n_4843),
.Y(n_11408)
);

AOI21xp5_ASAP7_75t_L g11409 ( 
.A1(n_10324),
.A2(n_4845),
.B(n_4844),
.Y(n_11409)
);

INVx1_ASAP7_75t_L g11410 ( 
.A(n_10291),
.Y(n_11410)
);

NAND2xp5_ASAP7_75t_L g11411 ( 
.A(n_10229),
.B(n_521),
.Y(n_11411)
);

OAI21xp5_ASAP7_75t_L g11412 ( 
.A1(n_10276),
.A2(n_521),
.B(n_522),
.Y(n_11412)
);

INVx1_ASAP7_75t_SL g11413 ( 
.A(n_10215),
.Y(n_11413)
);

INVx1_ASAP7_75t_L g11414 ( 
.A(n_10291),
.Y(n_11414)
);

NAND2xp5_ASAP7_75t_SL g11415 ( 
.A(n_10229),
.B(n_4846),
.Y(n_11415)
);

AOI21xp5_ASAP7_75t_L g11416 ( 
.A1(n_10324),
.A2(n_4849),
.B(n_4847),
.Y(n_11416)
);

NAND2xp5_ASAP7_75t_L g11417 ( 
.A(n_10229),
.B(n_522),
.Y(n_11417)
);

OAI21xp5_ASAP7_75t_L g11418 ( 
.A1(n_10276),
.A2(n_523),
.B(n_524),
.Y(n_11418)
);

AND2x2_ASAP7_75t_L g11419 ( 
.A(n_10310),
.B(n_4850),
.Y(n_11419)
);

INVx1_ASAP7_75t_L g11420 ( 
.A(n_10291),
.Y(n_11420)
);

AOI21xp5_ASAP7_75t_L g11421 ( 
.A1(n_10324),
.A2(n_4852),
.B(n_4851),
.Y(n_11421)
);

AOI21xp5_ASAP7_75t_L g11422 ( 
.A1(n_10324),
.A2(n_4854),
.B(n_4853),
.Y(n_11422)
);

NOR2xp67_ASAP7_75t_L g11423 ( 
.A(n_10280),
.B(n_4855),
.Y(n_11423)
);

A2O1A1Ixp33_ASAP7_75t_L g11424 ( 
.A1(n_10276),
.A2(n_525),
.B(n_523),
.C(n_524),
.Y(n_11424)
);

INVx2_ASAP7_75t_L g11425 ( 
.A(n_10220),
.Y(n_11425)
);

OAI21xp33_ASAP7_75t_SL g11426 ( 
.A1(n_10242),
.A2(n_525),
.B(n_526),
.Y(n_11426)
);

AO32x2_ASAP7_75t_L g11427 ( 
.A1(n_10815),
.A2(n_528),
.A3(n_526),
.B1(n_527),
.B2(n_529),
.Y(n_11427)
);

NAND2xp5_ASAP7_75t_SL g11428 ( 
.A(n_10229),
.B(n_4856),
.Y(n_11428)
);

AOI21xp5_ASAP7_75t_L g11429 ( 
.A1(n_10324),
.A2(n_4858),
.B(n_4857),
.Y(n_11429)
);

AOI21x1_ASAP7_75t_L g11430 ( 
.A1(n_10392),
.A2(n_4860),
.B(n_4859),
.Y(n_11430)
);

NOR2xp67_ASAP7_75t_L g11431 ( 
.A(n_10280),
.B(n_4861),
.Y(n_11431)
);

AOI21xp5_ASAP7_75t_L g11432 ( 
.A1(n_10324),
.A2(n_4863),
.B(n_4862),
.Y(n_11432)
);

OAI22xp5_ASAP7_75t_L g11433 ( 
.A1(n_10276),
.A2(n_530),
.B1(n_527),
.B2(n_529),
.Y(n_11433)
);

NAND2xp5_ASAP7_75t_SL g11434 ( 
.A(n_10229),
.B(n_4864),
.Y(n_11434)
);

NAND2xp5_ASAP7_75t_L g11435 ( 
.A(n_10229),
.B(n_530),
.Y(n_11435)
);

AOI21xp5_ASAP7_75t_L g11436 ( 
.A1(n_10324),
.A2(n_4866),
.B(n_4865),
.Y(n_11436)
);

AOI21xp5_ASAP7_75t_L g11437 ( 
.A1(n_10324),
.A2(n_4869),
.B(n_4867),
.Y(n_11437)
);

OAI21xp5_ASAP7_75t_L g11438 ( 
.A1(n_10276),
.A2(n_531),
.B(n_532),
.Y(n_11438)
);

HB1xp67_ASAP7_75t_L g11439 ( 
.A(n_10217),
.Y(n_11439)
);

NOR3xp33_ASAP7_75t_L g11440 ( 
.A(n_10276),
.B(n_531),
.C(n_532),
.Y(n_11440)
);

INVx1_ASAP7_75t_L g11441 ( 
.A(n_10291),
.Y(n_11441)
);

OAI22xp5_ASAP7_75t_L g11442 ( 
.A1(n_10276),
.A2(n_535),
.B1(n_533),
.B2(n_534),
.Y(n_11442)
);

INVx2_ASAP7_75t_L g11443 ( 
.A(n_10220),
.Y(n_11443)
);

OAI21xp5_ASAP7_75t_L g11444 ( 
.A1(n_10276),
.A2(n_533),
.B(n_534),
.Y(n_11444)
);

INVx1_ASAP7_75t_L g11445 ( 
.A(n_10291),
.Y(n_11445)
);

AND2x2_ASAP7_75t_L g11446 ( 
.A(n_10310),
.B(n_4870),
.Y(n_11446)
);

NOR2x1p5_ASAP7_75t_L g11447 ( 
.A(n_10699),
.B(n_4871),
.Y(n_11447)
);

BUFx12f_ASAP7_75t_L g11448 ( 
.A(n_10382),
.Y(n_11448)
);

AND2x2_ASAP7_75t_L g11449 ( 
.A(n_10310),
.B(n_4872),
.Y(n_11449)
);

HB1xp67_ASAP7_75t_L g11450 ( 
.A(n_10217),
.Y(n_11450)
);

CKINVDCx5p33_ASAP7_75t_R g11451 ( 
.A(n_10350),
.Y(n_11451)
);

INVx2_ASAP7_75t_L g11452 ( 
.A(n_10220),
.Y(n_11452)
);

NAND2xp5_ASAP7_75t_L g11453 ( 
.A(n_10229),
.B(n_535),
.Y(n_11453)
);

INVx2_ASAP7_75t_L g11454 ( 
.A(n_10220),
.Y(n_11454)
);

CKINVDCx8_ASAP7_75t_R g11455 ( 
.A(n_10283),
.Y(n_11455)
);

AND2x2_ASAP7_75t_L g11456 ( 
.A(n_10310),
.B(n_4873),
.Y(n_11456)
);

NAND2xp5_ASAP7_75t_SL g11457 ( 
.A(n_10229),
.B(n_4874),
.Y(n_11457)
);

INVx1_ASAP7_75t_L g11458 ( 
.A(n_10291),
.Y(n_11458)
);

OAI21xp5_ASAP7_75t_L g11459 ( 
.A1(n_10276),
.A2(n_536),
.B(n_537),
.Y(n_11459)
);

BUFx6f_ASAP7_75t_L g11460 ( 
.A(n_10318),
.Y(n_11460)
);

NAND2xp5_ASAP7_75t_L g11461 ( 
.A(n_10229),
.B(n_536),
.Y(n_11461)
);

NAND2xp5_ASAP7_75t_SL g11462 ( 
.A(n_10229),
.B(n_4875),
.Y(n_11462)
);

OAI21xp5_ASAP7_75t_L g11463 ( 
.A1(n_10276),
.A2(n_537),
.B(n_539),
.Y(n_11463)
);

NOR2xp33_ASAP7_75t_SL g11464 ( 
.A(n_10717),
.B(n_4876),
.Y(n_11464)
);

NAND2xp5_ASAP7_75t_L g11465 ( 
.A(n_10229),
.B(n_539),
.Y(n_11465)
);

NAND2xp5_ASAP7_75t_L g11466 ( 
.A(n_10229),
.B(n_540),
.Y(n_11466)
);

NOR3xp33_ASAP7_75t_L g11467 ( 
.A(n_10276),
.B(n_540),
.C(n_541),
.Y(n_11467)
);

NAND2xp5_ASAP7_75t_SL g11468 ( 
.A(n_10229),
.B(n_4877),
.Y(n_11468)
);

AOI22xp5_ASAP7_75t_L g11469 ( 
.A1(n_10276),
.A2(n_543),
.B1(n_541),
.B2(n_542),
.Y(n_11469)
);

AOI21xp5_ASAP7_75t_L g11470 ( 
.A1(n_10324),
.A2(n_4879),
.B(n_4878),
.Y(n_11470)
);

CKINVDCx10_ASAP7_75t_R g11471 ( 
.A(n_10296),
.Y(n_11471)
);

INVx1_ASAP7_75t_L g11472 ( 
.A(n_10291),
.Y(n_11472)
);

AOI21xp5_ASAP7_75t_L g11473 ( 
.A1(n_10324),
.A2(n_4883),
.B(n_4881),
.Y(n_11473)
);

INVx2_ASAP7_75t_L g11474 ( 
.A(n_10220),
.Y(n_11474)
);

AOI21xp5_ASAP7_75t_L g11475 ( 
.A1(n_10324),
.A2(n_4886),
.B(n_4885),
.Y(n_11475)
);

CKINVDCx5p33_ASAP7_75t_R g11476 ( 
.A(n_10350),
.Y(n_11476)
);

AOI21xp5_ASAP7_75t_L g11477 ( 
.A1(n_10324),
.A2(n_4889),
.B(n_4887),
.Y(n_11477)
);

NAND2xp5_ASAP7_75t_L g11478 ( 
.A(n_10229),
.B(n_543),
.Y(n_11478)
);

AOI21x1_ASAP7_75t_L g11479 ( 
.A1(n_10392),
.A2(n_4892),
.B(n_4890),
.Y(n_11479)
);

OAI21xp5_ASAP7_75t_L g11480 ( 
.A1(n_10276),
.A2(n_544),
.B(n_546),
.Y(n_11480)
);

NAND2xp5_ASAP7_75t_SL g11481 ( 
.A(n_10229),
.B(n_4893),
.Y(n_11481)
);

BUFx12f_ASAP7_75t_L g11482 ( 
.A(n_10382),
.Y(n_11482)
);

NAND2xp5_ASAP7_75t_L g11483 ( 
.A(n_10229),
.B(n_544),
.Y(n_11483)
);

NOR2xp33_ASAP7_75t_L g11484 ( 
.A(n_10276),
.B(n_4894),
.Y(n_11484)
);

NOR2xp33_ASAP7_75t_L g11485 ( 
.A(n_10276),
.B(n_4895),
.Y(n_11485)
);

AND2x2_ASAP7_75t_L g11486 ( 
.A(n_10310),
.B(n_4896),
.Y(n_11486)
);

AOI21xp5_ASAP7_75t_L g11487 ( 
.A1(n_10324),
.A2(n_4901),
.B(n_4898),
.Y(n_11487)
);

NAND2xp5_ASAP7_75t_L g11488 ( 
.A(n_10229),
.B(n_546),
.Y(n_11488)
);

AOI21xp33_ASAP7_75t_L g11489 ( 
.A1(n_10276),
.A2(n_547),
.B(n_548),
.Y(n_11489)
);

NAND2xp5_ASAP7_75t_L g11490 ( 
.A(n_10229),
.B(n_547),
.Y(n_11490)
);

OAI22xp5_ASAP7_75t_L g11491 ( 
.A1(n_10276),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.Y(n_11491)
);

BUFx6f_ASAP7_75t_L g11492 ( 
.A(n_10318),
.Y(n_11492)
);

OAI21xp5_ASAP7_75t_L g11493 ( 
.A1(n_10276),
.A2(n_549),
.B(n_550),
.Y(n_11493)
);

AOI21xp5_ASAP7_75t_L g11494 ( 
.A1(n_10324),
.A2(n_4903),
.B(n_4902),
.Y(n_11494)
);

INVx1_ASAP7_75t_L g11495 ( 
.A(n_10291),
.Y(n_11495)
);

NAND2xp5_ASAP7_75t_L g11496 ( 
.A(n_10229),
.B(n_551),
.Y(n_11496)
);

AOI21x1_ASAP7_75t_L g11497 ( 
.A1(n_10392),
.A2(n_4905),
.B(n_4904),
.Y(n_11497)
);

AOI21x1_ASAP7_75t_L g11498 ( 
.A1(n_10392),
.A2(n_4907),
.B(n_4906),
.Y(n_11498)
);

INVx2_ASAP7_75t_SL g11499 ( 
.A(n_10540),
.Y(n_11499)
);

AOI21x1_ASAP7_75t_L g11500 ( 
.A1(n_10392),
.A2(n_4909),
.B(n_4908),
.Y(n_11500)
);

NOR3xp33_ASAP7_75t_L g11501 ( 
.A(n_10276),
.B(n_551),
.C(n_552),
.Y(n_11501)
);

NOR2xp33_ASAP7_75t_L g11502 ( 
.A(n_10276),
.B(n_4910),
.Y(n_11502)
);

HB1xp67_ASAP7_75t_L g11503 ( 
.A(n_10217),
.Y(n_11503)
);

OAI21xp5_ASAP7_75t_L g11504 ( 
.A1(n_10276),
.A2(n_553),
.B(n_554),
.Y(n_11504)
);

OAI22xp5_ASAP7_75t_L g11505 ( 
.A1(n_10276),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.Y(n_11505)
);

NAND2xp5_ASAP7_75t_L g11506 ( 
.A(n_10229),
.B(n_555),
.Y(n_11506)
);

AOI21xp5_ASAP7_75t_L g11507 ( 
.A1(n_10324),
.A2(n_4913),
.B(n_4912),
.Y(n_11507)
);

AND2x4_ASAP7_75t_L g11508 ( 
.A(n_10380),
.B(n_4914),
.Y(n_11508)
);

NAND2xp5_ASAP7_75t_L g11509 ( 
.A(n_10229),
.B(n_556),
.Y(n_11509)
);

INVx2_ASAP7_75t_L g11510 ( 
.A(n_10220),
.Y(n_11510)
);

INVx1_ASAP7_75t_L g11511 ( 
.A(n_10291),
.Y(n_11511)
);

AOI21xp5_ASAP7_75t_L g11512 ( 
.A1(n_10324),
.A2(n_4916),
.B(n_4915),
.Y(n_11512)
);

BUFx4f_ASAP7_75t_L g11513 ( 
.A(n_10267),
.Y(n_11513)
);

INVx1_ASAP7_75t_L g11514 ( 
.A(n_10291),
.Y(n_11514)
);

AOI21xp5_ASAP7_75t_L g11515 ( 
.A1(n_10324),
.A2(n_4918),
.B(n_4917),
.Y(n_11515)
);

AOI21xp5_ASAP7_75t_L g11516 ( 
.A1(n_10324),
.A2(n_4920),
.B(n_4919),
.Y(n_11516)
);

AOI222xp33_ASAP7_75t_L g11517 ( 
.A1(n_10276),
.A2(n_558),
.B1(n_560),
.B2(n_556),
.C1(n_557),
.C2(n_559),
.Y(n_11517)
);

A2O1A1Ixp33_ASAP7_75t_L g11518 ( 
.A1(n_10276),
.A2(n_559),
.B(n_557),
.C(n_558),
.Y(n_11518)
);

AOI21xp5_ASAP7_75t_L g11519 ( 
.A1(n_10324),
.A2(n_4922),
.B(n_4921),
.Y(n_11519)
);

BUFx2_ASAP7_75t_L g11520 ( 
.A(n_10249),
.Y(n_11520)
);

AOI21xp5_ASAP7_75t_L g11521 ( 
.A1(n_10324),
.A2(n_4924),
.B(n_4923),
.Y(n_11521)
);

OAI21x1_ASAP7_75t_L g11522 ( 
.A1(n_10587),
.A2(n_4926),
.B(n_4925),
.Y(n_11522)
);

OAI21xp5_ASAP7_75t_L g11523 ( 
.A1(n_10276),
.A2(n_560),
.B(n_561),
.Y(n_11523)
);

AOI21xp5_ASAP7_75t_L g11524 ( 
.A1(n_10324),
.A2(n_4928),
.B(n_4927),
.Y(n_11524)
);

AOI22xp33_ASAP7_75t_L g11525 ( 
.A1(n_10276),
.A2(n_563),
.B1(n_561),
.B2(n_562),
.Y(n_11525)
);

BUFx8_ASAP7_75t_L g11526 ( 
.A(n_10523),
.Y(n_11526)
);

O2A1O1Ixp33_ASAP7_75t_L g11527 ( 
.A1(n_10276),
.A2(n_564),
.B(n_562),
.C(n_563),
.Y(n_11527)
);

NAND2xp5_ASAP7_75t_L g11528 ( 
.A(n_10229),
.B(n_564),
.Y(n_11528)
);

AND2x4_ASAP7_75t_L g11529 ( 
.A(n_10380),
.B(n_4929),
.Y(n_11529)
);

NAND2xp5_ASAP7_75t_L g11530 ( 
.A(n_10229),
.B(n_565),
.Y(n_11530)
);

BUFx6f_ASAP7_75t_L g11531 ( 
.A(n_10318),
.Y(n_11531)
);

INVx2_ASAP7_75t_L g11532 ( 
.A(n_10220),
.Y(n_11532)
);

NAND2xp5_ASAP7_75t_SL g11533 ( 
.A(n_10229),
.B(n_4930),
.Y(n_11533)
);

O2A1O1Ixp33_ASAP7_75t_L g11534 ( 
.A1(n_10276),
.A2(n_568),
.B(n_566),
.C(n_567),
.Y(n_11534)
);

OAI22xp5_ASAP7_75t_L g11535 ( 
.A1(n_10276),
.A2(n_569),
.B1(n_566),
.B2(n_568),
.Y(n_11535)
);

AOI21xp5_ASAP7_75t_L g11536 ( 
.A1(n_10324),
.A2(n_4932),
.B(n_4931),
.Y(n_11536)
);

AOI22xp5_ASAP7_75t_L g11537 ( 
.A1(n_10276),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_11537)
);

AOI21xp5_ASAP7_75t_L g11538 ( 
.A1(n_10324),
.A2(n_4934),
.B(n_4933),
.Y(n_11538)
);

A2O1A1Ixp33_ASAP7_75t_L g11539 ( 
.A1(n_10276),
.A2(n_574),
.B(n_572),
.C(n_573),
.Y(n_11539)
);

OR2x2_ASAP7_75t_L g11540 ( 
.A(n_10217),
.B(n_572),
.Y(n_11540)
);

AND2x2_ASAP7_75t_L g11541 ( 
.A(n_10310),
.B(n_4935),
.Y(n_11541)
);

INVx2_ASAP7_75t_L g11542 ( 
.A(n_10220),
.Y(n_11542)
);

AOI21xp5_ASAP7_75t_L g11543 ( 
.A1(n_10324),
.A2(n_4937),
.B(n_4936),
.Y(n_11543)
);

INVx2_ASAP7_75t_L g11544 ( 
.A(n_10220),
.Y(n_11544)
);

NAND2xp5_ASAP7_75t_L g11545 ( 
.A(n_10229),
.B(n_573),
.Y(n_11545)
);

INVx2_ASAP7_75t_L g11546 ( 
.A(n_10220),
.Y(n_11546)
);

NAND2xp5_ASAP7_75t_SL g11547 ( 
.A(n_10229),
.B(n_4938),
.Y(n_11547)
);

OAI22xp5_ASAP7_75t_L g11548 ( 
.A1(n_10276),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_11548)
);

AOI22xp5_ASAP7_75t_L g11549 ( 
.A1(n_10276),
.A2(n_578),
.B1(n_575),
.B2(n_577),
.Y(n_11549)
);

O2A1O1Ixp33_ASAP7_75t_L g11550 ( 
.A1(n_10276),
.A2(n_581),
.B(n_579),
.C(n_580),
.Y(n_11550)
);

NAND2xp5_ASAP7_75t_SL g11551 ( 
.A(n_10229),
.B(n_4939),
.Y(n_11551)
);

OAI22x1_ASAP7_75t_L g11552 ( 
.A1(n_10255),
.A2(n_581),
.B1(n_579),
.B2(n_580),
.Y(n_11552)
);

INVx1_ASAP7_75t_L g11553 ( 
.A(n_10291),
.Y(n_11553)
);

A2O1A1Ixp33_ASAP7_75t_L g11554 ( 
.A1(n_10276),
.A2(n_584),
.B(n_582),
.C(n_583),
.Y(n_11554)
);

O2A1O1Ixp33_ASAP7_75t_L g11555 ( 
.A1(n_10276),
.A2(n_584),
.B(n_582),
.C(n_583),
.Y(n_11555)
);

NAND2xp5_ASAP7_75t_L g11556 ( 
.A(n_10229),
.B(n_585),
.Y(n_11556)
);

AOI21xp5_ASAP7_75t_L g11557 ( 
.A1(n_10324),
.A2(n_4942),
.B(n_4940),
.Y(n_11557)
);

AOI21xp5_ASAP7_75t_L g11558 ( 
.A1(n_10324),
.A2(n_4944),
.B(n_4943),
.Y(n_11558)
);

INVx11_ASAP7_75t_L g11559 ( 
.A(n_10540),
.Y(n_11559)
);

INVx2_ASAP7_75t_L g11560 ( 
.A(n_10220),
.Y(n_11560)
);

AOI21xp5_ASAP7_75t_L g11561 ( 
.A1(n_10324),
.A2(n_4946),
.B(n_4945),
.Y(n_11561)
);

NAND2xp5_ASAP7_75t_L g11562 ( 
.A(n_10229),
.B(n_585),
.Y(n_11562)
);

NAND2xp5_ASAP7_75t_SL g11563 ( 
.A(n_10229),
.B(n_4947),
.Y(n_11563)
);

INVx2_ASAP7_75t_L g11564 ( 
.A(n_10220),
.Y(n_11564)
);

BUFx2_ASAP7_75t_L g11565 ( 
.A(n_10249),
.Y(n_11565)
);

NAND2xp5_ASAP7_75t_SL g11566 ( 
.A(n_10229),
.B(n_4949),
.Y(n_11566)
);

AOI22xp5_ASAP7_75t_L g11567 ( 
.A1(n_10276),
.A2(n_588),
.B1(n_586),
.B2(n_587),
.Y(n_11567)
);

NAND2xp5_ASAP7_75t_SL g11568 ( 
.A(n_10229),
.B(n_4951),
.Y(n_11568)
);

AOI21xp5_ASAP7_75t_L g11569 ( 
.A1(n_10324),
.A2(n_4953),
.B(n_4952),
.Y(n_11569)
);

CKINVDCx5p33_ASAP7_75t_R g11570 ( 
.A(n_10350),
.Y(n_11570)
);

NAND2xp5_ASAP7_75t_L g11571 ( 
.A(n_10229),
.B(n_586),
.Y(n_11571)
);

AOI21xp5_ASAP7_75t_L g11572 ( 
.A1(n_10324),
.A2(n_4955),
.B(n_4954),
.Y(n_11572)
);

OAI21xp5_ASAP7_75t_L g11573 ( 
.A1(n_10276),
.A2(n_587),
.B(n_588),
.Y(n_11573)
);

AOI21xp5_ASAP7_75t_L g11574 ( 
.A1(n_10324),
.A2(n_4958),
.B(n_4956),
.Y(n_11574)
);

INVx1_ASAP7_75t_L g11575 ( 
.A(n_10291),
.Y(n_11575)
);

NAND2xp5_ASAP7_75t_L g11576 ( 
.A(n_10229),
.B(n_589),
.Y(n_11576)
);

NAND2xp5_ASAP7_75t_L g11577 ( 
.A(n_10229),
.B(n_589),
.Y(n_11577)
);

AOI21xp5_ASAP7_75t_L g11578 ( 
.A1(n_10324),
.A2(n_4960),
.B(n_4959),
.Y(n_11578)
);

INVx3_ASAP7_75t_L g11579 ( 
.A(n_10227),
.Y(n_11579)
);

NAND2xp5_ASAP7_75t_L g11580 ( 
.A(n_10229),
.B(n_590),
.Y(n_11580)
);

NAND2xp5_ASAP7_75t_L g11581 ( 
.A(n_10229),
.B(n_590),
.Y(n_11581)
);

INVx2_ASAP7_75t_L g11582 ( 
.A(n_10220),
.Y(n_11582)
);

AOI21xp5_ASAP7_75t_L g11583 ( 
.A1(n_10324),
.A2(n_4962),
.B(n_4961),
.Y(n_11583)
);

A2O1A1Ixp33_ASAP7_75t_L g11584 ( 
.A1(n_10276),
.A2(n_593),
.B(n_591),
.C(n_592),
.Y(n_11584)
);

AOI21xp5_ASAP7_75t_L g11585 ( 
.A1(n_10324),
.A2(n_4964),
.B(n_4963),
.Y(n_11585)
);

NAND2xp5_ASAP7_75t_L g11586 ( 
.A(n_10229),
.B(n_591),
.Y(n_11586)
);

AOI21x1_ASAP7_75t_L g11587 ( 
.A1(n_10392),
.A2(n_4967),
.B(n_4966),
.Y(n_11587)
);

AOI21xp5_ASAP7_75t_L g11588 ( 
.A1(n_10324),
.A2(n_4970),
.B(n_4968),
.Y(n_11588)
);

AOI21xp5_ASAP7_75t_L g11589 ( 
.A1(n_10324),
.A2(n_4973),
.B(n_4971),
.Y(n_11589)
);

NAND2x1p5_ASAP7_75t_L g11590 ( 
.A(n_10283),
.B(n_4975),
.Y(n_11590)
);

NAND2xp5_ASAP7_75t_L g11591 ( 
.A(n_10229),
.B(n_592),
.Y(n_11591)
);

AOI21xp5_ASAP7_75t_L g11592 ( 
.A1(n_10324),
.A2(n_4977),
.B(n_4976),
.Y(n_11592)
);

NAND2xp5_ASAP7_75t_L g11593 ( 
.A(n_10229),
.B(n_594),
.Y(n_11593)
);

OAI21xp5_ASAP7_75t_L g11594 ( 
.A1(n_10276),
.A2(n_594),
.B(n_595),
.Y(n_11594)
);

OAI21xp5_ASAP7_75t_L g11595 ( 
.A1(n_10276),
.A2(n_595),
.B(n_596),
.Y(n_11595)
);

AOI21xp5_ASAP7_75t_L g11596 ( 
.A1(n_10324),
.A2(n_4981),
.B(n_4978),
.Y(n_11596)
);

INVx2_ASAP7_75t_L g11597 ( 
.A(n_10220),
.Y(n_11597)
);

NOR3xp33_ASAP7_75t_L g11598 ( 
.A(n_10276),
.B(n_596),
.C(n_597),
.Y(n_11598)
);

AND2x6_ASAP7_75t_L g11599 ( 
.A(n_10598),
.B(n_4982),
.Y(n_11599)
);

INVx3_ASAP7_75t_L g11600 ( 
.A(n_10227),
.Y(n_11600)
);

AOI21x1_ASAP7_75t_L g11601 ( 
.A1(n_10392),
.A2(n_4985),
.B(n_4984),
.Y(n_11601)
);

NAND2xp5_ASAP7_75t_L g11602 ( 
.A(n_10229),
.B(n_597),
.Y(n_11602)
);

AOI21xp5_ASAP7_75t_L g11603 ( 
.A1(n_10324),
.A2(n_4987),
.B(n_4986),
.Y(n_11603)
);

AOI21xp5_ASAP7_75t_L g11604 ( 
.A1(n_10855),
.A2(n_4990),
.B(n_4988),
.Y(n_11604)
);

NAND2xp5_ASAP7_75t_SL g11605 ( 
.A(n_10826),
.B(n_4992),
.Y(n_11605)
);

NAND2xp5_ASAP7_75t_L g11606 ( 
.A(n_11015),
.B(n_598),
.Y(n_11606)
);

INVx1_ASAP7_75t_L g11607 ( 
.A(n_11111),
.Y(n_11607)
);

NOR2xp33_ASAP7_75t_L g11608 ( 
.A(n_10856),
.B(n_598),
.Y(n_11608)
);

AOI22xp5_ASAP7_75t_L g11609 ( 
.A1(n_11440),
.A2(n_601),
.B1(n_599),
.B2(n_600),
.Y(n_11609)
);

AOI21xp5_ASAP7_75t_L g11610 ( 
.A1(n_10839),
.A2(n_4995),
.B(n_4993),
.Y(n_11610)
);

OAI22xp5_ASAP7_75t_L g11611 ( 
.A1(n_11383),
.A2(n_602),
.B1(n_599),
.B2(n_601),
.Y(n_11611)
);

A2O1A1Ixp33_ASAP7_75t_L g11612 ( 
.A1(n_11527),
.A2(n_604),
.B(n_602),
.C(n_603),
.Y(n_11612)
);

NAND2xp5_ASAP7_75t_L g11613 ( 
.A(n_11060),
.B(n_605),
.Y(n_11613)
);

BUFx6f_ASAP7_75t_L g11614 ( 
.A(n_11398),
.Y(n_11614)
);

A2O1A1Ixp33_ASAP7_75t_L g11615 ( 
.A1(n_11534),
.A2(n_11555),
.B(n_11550),
.C(n_11412),
.Y(n_11615)
);

AOI22xp5_ASAP7_75t_L g11616 ( 
.A1(n_11467),
.A2(n_607),
.B1(n_605),
.B2(n_606),
.Y(n_11616)
);

AOI21xp5_ASAP7_75t_L g11617 ( 
.A1(n_10945),
.A2(n_5000),
.B(n_4996),
.Y(n_11617)
);

A2O1A1Ixp33_ASAP7_75t_SL g11618 ( 
.A1(n_11501),
.A2(n_608),
.B(n_606),
.C(n_607),
.Y(n_11618)
);

OR2x6_ASAP7_75t_SL g11619 ( 
.A(n_11451),
.B(n_608),
.Y(n_11619)
);

AOI21xp5_ASAP7_75t_L g11620 ( 
.A1(n_11095),
.A2(n_5002),
.B(n_5001),
.Y(n_11620)
);

A2O1A1Ixp33_ASAP7_75t_L g11621 ( 
.A1(n_11396),
.A2(n_612),
.B(n_609),
.C(n_610),
.Y(n_11621)
);

NOR2xp33_ASAP7_75t_SL g11622 ( 
.A(n_11051),
.B(n_5003),
.Y(n_11622)
);

NAND2xp5_ASAP7_75t_L g11623 ( 
.A(n_10949),
.B(n_609),
.Y(n_11623)
);

OAI21xp33_ASAP7_75t_L g11624 ( 
.A1(n_11598),
.A2(n_610),
.B(n_612),
.Y(n_11624)
);

INVx1_ASAP7_75t_L g11625 ( 
.A(n_11186),
.Y(n_11625)
);

AND2x2_ASAP7_75t_L g11626 ( 
.A(n_10859),
.B(n_613),
.Y(n_11626)
);

INVx1_ASAP7_75t_L g11627 ( 
.A(n_11246),
.Y(n_11627)
);

INVx2_ASAP7_75t_SL g11628 ( 
.A(n_11211),
.Y(n_11628)
);

A2O1A1Ixp33_ASAP7_75t_L g11629 ( 
.A1(n_11418),
.A2(n_615),
.B(n_613),
.C(n_614),
.Y(n_11629)
);

INVx2_ASAP7_75t_L g11630 ( 
.A(n_11266),
.Y(n_11630)
);

AOI21xp5_ASAP7_75t_L g11631 ( 
.A1(n_10828),
.A2(n_5005),
.B(n_5004),
.Y(n_11631)
);

AOI21xp5_ASAP7_75t_L g11632 ( 
.A1(n_11438),
.A2(n_5008),
.B(n_5007),
.Y(n_11632)
);

INVx1_ASAP7_75t_L g11633 ( 
.A(n_11245),
.Y(n_11633)
);

NAND2xp5_ASAP7_75t_L g11634 ( 
.A(n_11439),
.B(n_615),
.Y(n_11634)
);

NAND2xp5_ASAP7_75t_L g11635 ( 
.A(n_11450),
.B(n_616),
.Y(n_11635)
);

NAND2xp5_ASAP7_75t_L g11636 ( 
.A(n_11503),
.B(n_616),
.Y(n_11636)
);

NAND2xp5_ASAP7_75t_L g11637 ( 
.A(n_10907),
.B(n_617),
.Y(n_11637)
);

NOR2xp33_ASAP7_75t_L g11638 ( 
.A(n_11389),
.B(n_617),
.Y(n_11638)
);

NAND2xp5_ASAP7_75t_L g11639 ( 
.A(n_10924),
.B(n_618),
.Y(n_11639)
);

AOI21xp5_ASAP7_75t_L g11640 ( 
.A1(n_11444),
.A2(n_5011),
.B(n_5010),
.Y(n_11640)
);

OAI22xp5_ASAP7_75t_L g11641 ( 
.A1(n_11021),
.A2(n_620),
.B1(n_618),
.B2(n_619),
.Y(n_11641)
);

INVx1_ASAP7_75t_L g11642 ( 
.A(n_10829),
.Y(n_11642)
);

NOR2xp67_ASAP7_75t_L g11643 ( 
.A(n_11076),
.B(n_619),
.Y(n_11643)
);

INVx1_ASAP7_75t_L g11644 ( 
.A(n_10834),
.Y(n_11644)
);

AOI21xp5_ASAP7_75t_L g11645 ( 
.A1(n_11459),
.A2(n_5013),
.B(n_5012),
.Y(n_11645)
);

OAI22xp5_ASAP7_75t_L g11646 ( 
.A1(n_11401),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_11646)
);

OAI21xp5_ASAP7_75t_L g11647 ( 
.A1(n_11385),
.A2(n_5015),
.B(n_5014),
.Y(n_11647)
);

OR2x2_ASAP7_75t_L g11648 ( 
.A(n_11413),
.B(n_622),
.Y(n_11648)
);

AOI21xp5_ASAP7_75t_L g11649 ( 
.A1(n_11463),
.A2(n_5017),
.B(n_5016),
.Y(n_11649)
);

NAND2xp5_ASAP7_75t_SL g11650 ( 
.A(n_11480),
.B(n_5020),
.Y(n_11650)
);

OAI21x1_ASAP7_75t_L g11651 ( 
.A1(n_10911),
.A2(n_5023),
.B(n_5022),
.Y(n_11651)
);

INVx1_ASAP7_75t_L g11652 ( 
.A(n_10866),
.Y(n_11652)
);

INVx1_ASAP7_75t_L g11653 ( 
.A(n_10912),
.Y(n_11653)
);

NOR2xp33_ASAP7_75t_L g11654 ( 
.A(n_11369),
.B(n_623),
.Y(n_11654)
);

OAI21x1_ASAP7_75t_L g11655 ( 
.A1(n_10994),
.A2(n_10982),
.B(n_11218),
.Y(n_11655)
);

OAI22xp5_ASAP7_75t_L g11656 ( 
.A1(n_11469),
.A2(n_11549),
.B1(n_11567),
.B2(n_11537),
.Y(n_11656)
);

AND2x2_ASAP7_75t_L g11657 ( 
.A(n_11363),
.B(n_624),
.Y(n_11657)
);

NAND2xp5_ASAP7_75t_SL g11658 ( 
.A(n_11493),
.B(n_5025),
.Y(n_11658)
);

AOI21xp5_ASAP7_75t_L g11659 ( 
.A1(n_11504),
.A2(n_5028),
.B(n_5026),
.Y(n_11659)
);

INVx1_ASAP7_75t_L g11660 ( 
.A(n_10917),
.Y(n_11660)
);

NAND2xp5_ASAP7_75t_L g11661 ( 
.A(n_10959),
.B(n_11014),
.Y(n_11661)
);

INVx1_ASAP7_75t_L g11662 ( 
.A(n_10948),
.Y(n_11662)
);

NAND2xp5_ASAP7_75t_L g11663 ( 
.A(n_10875),
.B(n_625),
.Y(n_11663)
);

AOI21xp5_ASAP7_75t_L g11664 ( 
.A1(n_11523),
.A2(n_5031),
.B(n_5029),
.Y(n_11664)
);

AOI22xp5_ASAP7_75t_L g11665 ( 
.A1(n_11391),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.Y(n_11665)
);

AND3x2_ASAP7_75t_L g11666 ( 
.A(n_11573),
.B(n_626),
.C(n_627),
.Y(n_11666)
);

NAND2xp5_ASAP7_75t_L g11667 ( 
.A(n_11520),
.B(n_628),
.Y(n_11667)
);

NAND2xp5_ASAP7_75t_L g11668 ( 
.A(n_11565),
.B(n_628),
.Y(n_11668)
);

AOI22xp5_ASAP7_75t_L g11669 ( 
.A1(n_11392),
.A2(n_631),
.B1(n_629),
.B2(n_630),
.Y(n_11669)
);

NAND2xp5_ASAP7_75t_SL g11670 ( 
.A(n_11594),
.B(n_5032),
.Y(n_11670)
);

BUFx2_ASAP7_75t_L g11671 ( 
.A(n_11046),
.Y(n_11671)
);

NAND2xp5_ASAP7_75t_SL g11672 ( 
.A(n_11595),
.B(n_5033),
.Y(n_11672)
);

AOI22xp5_ASAP7_75t_L g11673 ( 
.A1(n_11394),
.A2(n_631),
.B1(n_629),
.B2(n_630),
.Y(n_11673)
);

NAND2xp5_ASAP7_75t_L g11674 ( 
.A(n_10852),
.B(n_632),
.Y(n_11674)
);

OAI22xp5_ASAP7_75t_L g11675 ( 
.A1(n_11525),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.Y(n_11675)
);

NAND3xp33_ASAP7_75t_L g11676 ( 
.A(n_11399),
.B(n_634),
.C(n_635),
.Y(n_11676)
);

INVx3_ASAP7_75t_L g11677 ( 
.A(n_11398),
.Y(n_11677)
);

NOR2xp33_ASAP7_75t_L g11678 ( 
.A(n_10887),
.B(n_635),
.Y(n_11678)
);

NOR2xp33_ASAP7_75t_L g11679 ( 
.A(n_11406),
.B(n_637),
.Y(n_11679)
);

A2O1A1Ixp33_ASAP7_75t_L g11680 ( 
.A1(n_11400),
.A2(n_11485),
.B(n_11502),
.C(n_11484),
.Y(n_11680)
);

AOI22xp5_ASAP7_75t_L g11681 ( 
.A1(n_11166),
.A2(n_641),
.B1(n_638),
.B2(n_640),
.Y(n_11681)
);

AOI21x1_ASAP7_75t_L g11682 ( 
.A1(n_10872),
.A2(n_638),
.B(n_640),
.Y(n_11682)
);

AOI21xp5_ASAP7_75t_L g11683 ( 
.A1(n_11077),
.A2(n_5035),
.B(n_5034),
.Y(n_11683)
);

AOI21xp5_ASAP7_75t_L g11684 ( 
.A1(n_10969),
.A2(n_5037),
.B(n_5036),
.Y(n_11684)
);

NAND2xp5_ASAP7_75t_SL g11685 ( 
.A(n_11048),
.B(n_5038),
.Y(n_11685)
);

AOI21xp5_ASAP7_75t_L g11686 ( 
.A1(n_10980),
.A2(n_642),
.B(n_643),
.Y(n_11686)
);

INVxp67_ASAP7_75t_L g11687 ( 
.A(n_10962),
.Y(n_11687)
);

BUFx8_ASAP7_75t_L g11688 ( 
.A(n_10879),
.Y(n_11688)
);

NAND2xp5_ASAP7_75t_L g11689 ( 
.A(n_10892),
.B(n_11397),
.Y(n_11689)
);

OAI22xp5_ASAP7_75t_L g11690 ( 
.A1(n_10831),
.A2(n_10878),
.B1(n_11424),
.B2(n_11380),
.Y(n_11690)
);

BUFx4f_ASAP7_75t_L g11691 ( 
.A(n_11143),
.Y(n_11691)
);

NAND2xp5_ASAP7_75t_SL g11692 ( 
.A(n_11019),
.B(n_642),
.Y(n_11692)
);

BUFx6f_ASAP7_75t_L g11693 ( 
.A(n_10991),
.Y(n_11693)
);

NAND2xp5_ASAP7_75t_SL g11694 ( 
.A(n_10904),
.B(n_644),
.Y(n_11694)
);

A2O1A1Ixp33_ASAP7_75t_L g11695 ( 
.A1(n_10935),
.A2(n_646),
.B(n_644),
.C(n_645),
.Y(n_11695)
);

O2A1O1Ixp33_ASAP7_75t_L g11696 ( 
.A1(n_11518),
.A2(n_648),
.B(n_645),
.C(n_647),
.Y(n_11696)
);

OAI22xp33_ASAP7_75t_L g11697 ( 
.A1(n_11203),
.A2(n_650),
.B1(n_647),
.B2(n_649),
.Y(n_11697)
);

NAND2xp5_ASAP7_75t_SL g11698 ( 
.A(n_11136),
.B(n_649),
.Y(n_11698)
);

INVx2_ASAP7_75t_L g11699 ( 
.A(n_11237),
.Y(n_11699)
);

AOI21xp5_ASAP7_75t_L g11700 ( 
.A1(n_10842),
.A2(n_650),
.B(n_651),
.Y(n_11700)
);

NOR2xp33_ASAP7_75t_L g11701 ( 
.A(n_11579),
.B(n_652),
.Y(n_11701)
);

NOR3xp33_ASAP7_75t_L g11702 ( 
.A(n_11489),
.B(n_652),
.C(n_653),
.Y(n_11702)
);

INVxp67_ASAP7_75t_SL g11703 ( 
.A(n_11092),
.Y(n_11703)
);

CKINVDCx8_ASAP7_75t_R g11704 ( 
.A(n_11471),
.Y(n_11704)
);

BUFx12f_ASAP7_75t_L g11705 ( 
.A(n_11448),
.Y(n_11705)
);

O2A1O1Ixp5_ASAP7_75t_L g11706 ( 
.A1(n_11539),
.A2(n_656),
.B(n_654),
.C(n_655),
.Y(n_11706)
);

NAND2xp5_ASAP7_75t_L g11707 ( 
.A(n_11306),
.B(n_654),
.Y(n_11707)
);

NAND2xp5_ASAP7_75t_SL g11708 ( 
.A(n_11318),
.B(n_11310),
.Y(n_11708)
);

NOR2xp33_ASAP7_75t_L g11709 ( 
.A(n_11600),
.B(n_655),
.Y(n_11709)
);

OAI22xp5_ASAP7_75t_L g11710 ( 
.A1(n_11554),
.A2(n_658),
.B1(n_656),
.B2(n_657),
.Y(n_11710)
);

INVx1_ASAP7_75t_L g11711 ( 
.A(n_10951),
.Y(n_11711)
);

AOI21xp5_ASAP7_75t_L g11712 ( 
.A1(n_11138),
.A2(n_11160),
.B(n_11159),
.Y(n_11712)
);

NOR2xp33_ASAP7_75t_L g11713 ( 
.A(n_11156),
.B(n_657),
.Y(n_11713)
);

NAND2xp5_ASAP7_75t_SL g11714 ( 
.A(n_11318),
.B(n_658),
.Y(n_11714)
);

AOI21xp5_ASAP7_75t_L g11715 ( 
.A1(n_11172),
.A2(n_659),
.B(n_660),
.Y(n_11715)
);

NAND2xp5_ASAP7_75t_L g11716 ( 
.A(n_10920),
.B(n_659),
.Y(n_11716)
);

AOI21xp5_ASAP7_75t_L g11717 ( 
.A1(n_11105),
.A2(n_660),
.B(n_661),
.Y(n_11717)
);

AOI22xp5_ASAP7_75t_L g11718 ( 
.A1(n_11235),
.A2(n_11037),
.B1(n_11113),
.B2(n_10915),
.Y(n_11718)
);

INVx1_ASAP7_75t_L g11719 ( 
.A(n_10967),
.Y(n_11719)
);

NAND2xp5_ASAP7_75t_L g11720 ( 
.A(n_10979),
.B(n_661),
.Y(n_11720)
);

BUFx6f_ASAP7_75t_L g11721 ( 
.A(n_10991),
.Y(n_11721)
);

O2A1O1Ixp33_ASAP7_75t_L g11722 ( 
.A1(n_11584),
.A2(n_10847),
.B(n_11251),
.C(n_10964),
.Y(n_11722)
);

NAND2xp5_ASAP7_75t_L g11723 ( 
.A(n_11271),
.B(n_662),
.Y(n_11723)
);

NAND2xp5_ASAP7_75t_SL g11724 ( 
.A(n_11318),
.B(n_662),
.Y(n_11724)
);

AO32x1_ASAP7_75t_L g11725 ( 
.A1(n_11365),
.A2(n_665),
.A3(n_663),
.B1(n_664),
.B2(n_666),
.Y(n_11725)
);

AOI21xp5_ASAP7_75t_L g11726 ( 
.A1(n_11096),
.A2(n_663),
.B(n_664),
.Y(n_11726)
);

AND2x4_ASAP7_75t_L g11727 ( 
.A(n_11132),
.B(n_665),
.Y(n_11727)
);

NOR2xp33_ASAP7_75t_L g11728 ( 
.A(n_10884),
.B(n_666),
.Y(n_11728)
);

OAI22xp5_ASAP7_75t_L g11729 ( 
.A1(n_11347),
.A2(n_669),
.B1(n_667),
.B2(n_668),
.Y(n_11729)
);

NOR2xp33_ASAP7_75t_L g11730 ( 
.A(n_10954),
.B(n_10984),
.Y(n_11730)
);

O2A1O1Ixp33_ASAP7_75t_SL g11731 ( 
.A1(n_11372),
.A2(n_669),
.B(n_667),
.C(n_668),
.Y(n_11731)
);

AND2x2_ASAP7_75t_L g11732 ( 
.A(n_11370),
.B(n_670),
.Y(n_11732)
);

O2A1O1Ixp33_ASAP7_75t_L g11733 ( 
.A1(n_11207),
.A2(n_672),
.B(n_670),
.C(n_671),
.Y(n_11733)
);

INVx3_ASAP7_75t_L g11734 ( 
.A(n_10905),
.Y(n_11734)
);

NOR2xp33_ASAP7_75t_L g11735 ( 
.A(n_11087),
.B(n_671),
.Y(n_11735)
);

INVx1_ASAP7_75t_L g11736 ( 
.A(n_11010),
.Y(n_11736)
);

INVx2_ASAP7_75t_SL g11737 ( 
.A(n_11211),
.Y(n_11737)
);

BUFx3_ASAP7_75t_L g11738 ( 
.A(n_10991),
.Y(n_11738)
);

AOI21xp5_ASAP7_75t_L g11739 ( 
.A1(n_11100),
.A2(n_672),
.B(n_673),
.Y(n_11739)
);

INVx4_ASAP7_75t_L g11740 ( 
.A(n_11559),
.Y(n_11740)
);

AOI21xp5_ASAP7_75t_L g11741 ( 
.A1(n_10840),
.A2(n_10835),
.B(n_10843),
.Y(n_11741)
);

BUFx2_ASAP7_75t_L g11742 ( 
.A(n_10981),
.Y(n_11742)
);

BUFx2_ASAP7_75t_L g11743 ( 
.A(n_11017),
.Y(n_11743)
);

NAND2xp5_ASAP7_75t_L g11744 ( 
.A(n_11273),
.B(n_673),
.Y(n_11744)
);

BUFx12f_ASAP7_75t_L g11745 ( 
.A(n_11482),
.Y(n_11745)
);

NAND2xp5_ASAP7_75t_L g11746 ( 
.A(n_10961),
.B(n_674),
.Y(n_11746)
);

INVx1_ASAP7_75t_L g11747 ( 
.A(n_11011),
.Y(n_11747)
);

CKINVDCx20_ASAP7_75t_R g11748 ( 
.A(n_11476),
.Y(n_11748)
);

NAND2xp5_ASAP7_75t_L g11749 ( 
.A(n_10989),
.B(n_674),
.Y(n_11749)
);

INVx2_ASAP7_75t_L g11750 ( 
.A(n_11247),
.Y(n_11750)
);

NAND3xp33_ASAP7_75t_SL g11751 ( 
.A(n_11517),
.B(n_675),
.C(n_676),
.Y(n_11751)
);

OAI21x1_ASAP7_75t_L g11752 ( 
.A1(n_11119),
.A2(n_675),
.B(n_676),
.Y(n_11752)
);

AND2x2_ASAP7_75t_L g11753 ( 
.A(n_11317),
.B(n_677),
.Y(n_11753)
);

NAND2xp5_ASAP7_75t_L g11754 ( 
.A(n_10870),
.B(n_677),
.Y(n_11754)
);

NAND2xp5_ASAP7_75t_SL g11755 ( 
.A(n_11285),
.B(n_678),
.Y(n_11755)
);

INVx1_ASAP7_75t_L g11756 ( 
.A(n_11054),
.Y(n_11756)
);

OAI22xp5_ASAP7_75t_SL g11757 ( 
.A1(n_10928),
.A2(n_680),
.B1(n_678),
.B2(n_679),
.Y(n_11757)
);

AOI21xp5_ASAP7_75t_L g11758 ( 
.A1(n_10851),
.A2(n_679),
.B(n_680),
.Y(n_11758)
);

NOR2xp33_ASAP7_75t_L g11759 ( 
.A(n_11320),
.B(n_681),
.Y(n_11759)
);

NOR2xp33_ASAP7_75t_L g11760 ( 
.A(n_11342),
.B(n_681),
.Y(n_11760)
);

BUFx2_ASAP7_75t_SL g11761 ( 
.A(n_10919),
.Y(n_11761)
);

INVxp67_ASAP7_75t_SL g11762 ( 
.A(n_11003),
.Y(n_11762)
);

AOI21xp5_ASAP7_75t_L g11763 ( 
.A1(n_11085),
.A2(n_682),
.B(n_683),
.Y(n_11763)
);

NOR2xp33_ASAP7_75t_L g11764 ( 
.A(n_11067),
.B(n_683),
.Y(n_11764)
);

O2A1O1Ixp5_ASAP7_75t_L g11765 ( 
.A1(n_11231),
.A2(n_686),
.B(n_684),
.C(n_685),
.Y(n_11765)
);

NAND2xp5_ASAP7_75t_L g11766 ( 
.A(n_10916),
.B(n_684),
.Y(n_11766)
);

INVx1_ASAP7_75t_L g11767 ( 
.A(n_11055),
.Y(n_11767)
);

AOI22x1_ASAP7_75t_L g11768 ( 
.A1(n_11552),
.A2(n_687),
.B1(n_685),
.B2(n_686),
.Y(n_11768)
);

AOI22xp5_ASAP7_75t_L g11769 ( 
.A1(n_11135),
.A2(n_689),
.B1(n_687),
.B2(n_688),
.Y(n_11769)
);

NAND2xp5_ASAP7_75t_L g11770 ( 
.A(n_11334),
.B(n_690),
.Y(n_11770)
);

BUFx3_ASAP7_75t_L g11771 ( 
.A(n_11061),
.Y(n_11771)
);

NAND2xp5_ASAP7_75t_L g11772 ( 
.A(n_11255),
.B(n_690),
.Y(n_11772)
);

NAND2xp5_ASAP7_75t_L g11773 ( 
.A(n_11151),
.B(n_691),
.Y(n_11773)
);

AOI21xp5_ASAP7_75t_L g11774 ( 
.A1(n_11088),
.A2(n_691),
.B(n_692),
.Y(n_11774)
);

AO21x1_ASAP7_75t_L g11775 ( 
.A1(n_11377),
.A2(n_693),
.B(n_694),
.Y(n_11775)
);

CKINVDCx5p33_ASAP7_75t_R g11776 ( 
.A(n_11570),
.Y(n_11776)
);

AOI21xp5_ASAP7_75t_L g11777 ( 
.A1(n_10836),
.A2(n_693),
.B(n_694),
.Y(n_11777)
);

CKINVDCx6p67_ASAP7_75t_R g11778 ( 
.A(n_11214),
.Y(n_11778)
);

OAI22xp5_ASAP7_75t_L g11779 ( 
.A1(n_11281),
.A2(n_697),
.B1(n_695),
.B2(n_696),
.Y(n_11779)
);

BUFx8_ASAP7_75t_L g11780 ( 
.A(n_11206),
.Y(n_11780)
);

AOI22xp5_ASAP7_75t_L g11781 ( 
.A1(n_11009),
.A2(n_697),
.B1(n_695),
.B2(n_696),
.Y(n_11781)
);

O2A1O1Ixp33_ASAP7_75t_L g11782 ( 
.A1(n_11137),
.A2(n_700),
.B(n_698),
.C(n_699),
.Y(n_11782)
);

INVx2_ASAP7_75t_L g11783 ( 
.A(n_11261),
.Y(n_11783)
);

BUFx2_ASAP7_75t_SL g11784 ( 
.A(n_11455),
.Y(n_11784)
);

AOI21xp5_ASAP7_75t_L g11785 ( 
.A1(n_11351),
.A2(n_698),
.B(n_699),
.Y(n_11785)
);

NAND2xp5_ASAP7_75t_L g11786 ( 
.A(n_11053),
.B(n_700),
.Y(n_11786)
);

OAI21x1_ASAP7_75t_L g11787 ( 
.A1(n_11184),
.A2(n_701),
.B(n_702),
.Y(n_11787)
);

NAND2xp5_ASAP7_75t_L g11788 ( 
.A(n_11319),
.B(n_701),
.Y(n_11788)
);

NAND2xp5_ASAP7_75t_L g11789 ( 
.A(n_10833),
.B(n_702),
.Y(n_11789)
);

AOI21xp5_ASAP7_75t_L g11790 ( 
.A1(n_11202),
.A2(n_703),
.B(n_704),
.Y(n_11790)
);

INVx3_ASAP7_75t_L g11791 ( 
.A(n_10905),
.Y(n_11791)
);

AOI21xp5_ASAP7_75t_L g11792 ( 
.A1(n_11202),
.A2(n_704),
.B(n_705),
.Y(n_11792)
);

A2O1A1Ixp33_ASAP7_75t_L g11793 ( 
.A1(n_11213),
.A2(n_708),
.B(n_706),
.C(n_707),
.Y(n_11793)
);

NAND2xp5_ASAP7_75t_L g11794 ( 
.A(n_10891),
.B(n_707),
.Y(n_11794)
);

AOI21xp5_ASAP7_75t_L g11795 ( 
.A1(n_11229),
.A2(n_708),
.B(n_709),
.Y(n_11795)
);

NAND2xp5_ASAP7_75t_L g11796 ( 
.A(n_10903),
.B(n_709),
.Y(n_11796)
);

AND2x4_ASAP7_75t_L g11797 ( 
.A(n_11287),
.B(n_710),
.Y(n_11797)
);

O2A1O1Ixp33_ASAP7_75t_SL g11798 ( 
.A1(n_10968),
.A2(n_712),
.B(n_710),
.C(n_711),
.Y(n_11798)
);

NAND2xp5_ASAP7_75t_L g11799 ( 
.A(n_10926),
.B(n_711),
.Y(n_11799)
);

INVx2_ASAP7_75t_L g11800 ( 
.A(n_11058),
.Y(n_11800)
);

NOR2xp33_ASAP7_75t_L g11801 ( 
.A(n_11050),
.B(n_713),
.Y(n_11801)
);

NAND2xp5_ASAP7_75t_L g11802 ( 
.A(n_11005),
.B(n_713),
.Y(n_11802)
);

NAND2xp5_ASAP7_75t_SL g11803 ( 
.A(n_11099),
.B(n_714),
.Y(n_11803)
);

O2A1O1Ixp33_ASAP7_75t_L g11804 ( 
.A1(n_11179),
.A2(n_716),
.B(n_714),
.C(n_715),
.Y(n_11804)
);

OAI21xp5_ASAP7_75t_L g11805 ( 
.A1(n_11128),
.A2(n_715),
.B(n_716),
.Y(n_11805)
);

INVx1_ASAP7_75t_L g11806 ( 
.A(n_11059),
.Y(n_11806)
);

NOR2xp33_ASAP7_75t_SL g11807 ( 
.A(n_11147),
.B(n_717),
.Y(n_11807)
);

NOR2xp33_ASAP7_75t_L g11808 ( 
.A(n_11112),
.B(n_717),
.Y(n_11808)
);

AOI21xp5_ASAP7_75t_L g11809 ( 
.A1(n_10993),
.A2(n_718),
.B(n_719),
.Y(n_11809)
);

OAI22xp5_ASAP7_75t_L g11810 ( 
.A1(n_11264),
.A2(n_720),
.B1(n_718),
.B2(n_719),
.Y(n_11810)
);

NAND2xp5_ASAP7_75t_L g11811 ( 
.A(n_11006),
.B(n_721),
.Y(n_11811)
);

AOI21xp5_ASAP7_75t_L g11812 ( 
.A1(n_10993),
.A2(n_721),
.B(n_722),
.Y(n_11812)
);

INVx2_ASAP7_75t_L g11813 ( 
.A(n_11068),
.Y(n_11813)
);

O2A1O1Ixp5_ASAP7_75t_SL g11814 ( 
.A1(n_10972),
.A2(n_724),
.B(n_722),
.C(n_723),
.Y(n_11814)
);

OAI22xp5_ASAP7_75t_L g11815 ( 
.A1(n_11016),
.A2(n_726),
.B1(n_724),
.B2(n_725),
.Y(n_11815)
);

O2A1O1Ixp33_ASAP7_75t_L g11816 ( 
.A1(n_11224),
.A2(n_728),
.B(n_725),
.C(n_727),
.Y(n_11816)
);

NOR2xp33_ASAP7_75t_L g11817 ( 
.A(n_11086),
.B(n_727),
.Y(n_11817)
);

A2O1A1Ixp33_ASAP7_75t_L g11818 ( 
.A1(n_11198),
.A2(n_730),
.B(n_728),
.C(n_729),
.Y(n_11818)
);

AND2x4_ASAP7_75t_L g11819 ( 
.A(n_11368),
.B(n_729),
.Y(n_11819)
);

NAND2xp5_ASAP7_75t_L g11820 ( 
.A(n_11018),
.B(n_730),
.Y(n_11820)
);

OAI21xp5_ASAP7_75t_L g11821 ( 
.A1(n_10837),
.A2(n_731),
.B(n_732),
.Y(n_11821)
);

AOI21xp5_ASAP7_75t_L g11822 ( 
.A1(n_10947),
.A2(n_731),
.B(n_733),
.Y(n_11822)
);

INVx2_ASAP7_75t_L g11823 ( 
.A(n_11073),
.Y(n_11823)
);

HB1xp67_ASAP7_75t_L g11824 ( 
.A(n_11104),
.Y(n_11824)
);

OAI21x1_ASAP7_75t_L g11825 ( 
.A1(n_10881),
.A2(n_733),
.B(n_734),
.Y(n_11825)
);

AND2x4_ASAP7_75t_L g11826 ( 
.A(n_11064),
.B(n_735),
.Y(n_11826)
);

AND2x2_ASAP7_75t_L g11827 ( 
.A(n_11108),
.B(n_735),
.Y(n_11827)
);

INVx1_ASAP7_75t_L g11828 ( 
.A(n_11123),
.Y(n_11828)
);

NAND3xp33_ASAP7_75t_L g11829 ( 
.A(n_10965),
.B(n_736),
.C(n_737),
.Y(n_11829)
);

AOI22xp5_ASAP7_75t_L g11830 ( 
.A1(n_11381),
.A2(n_740),
.B1(n_738),
.B2(n_739),
.Y(n_11830)
);

NAND2xp5_ASAP7_75t_SL g11831 ( 
.A(n_11362),
.B(n_739),
.Y(n_11831)
);

NAND3xp33_ASAP7_75t_SL g11832 ( 
.A(n_11041),
.B(n_10930),
.C(n_10925),
.Y(n_11832)
);

BUFx3_ASAP7_75t_L g11833 ( 
.A(n_10853),
.Y(n_11833)
);

OAI22xp5_ASAP7_75t_L g11834 ( 
.A1(n_11102),
.A2(n_11289),
.B1(n_10880),
.B2(n_11190),
.Y(n_11834)
);

AOI22x1_ASAP7_75t_L g11835 ( 
.A1(n_11089),
.A2(n_742),
.B1(n_740),
.B2(n_741),
.Y(n_11835)
);

OAI21xp5_ASAP7_75t_L g11836 ( 
.A1(n_10825),
.A2(n_742),
.B(n_743),
.Y(n_11836)
);

OA22x2_ASAP7_75t_L g11837 ( 
.A1(n_11313),
.A2(n_745),
.B1(n_743),
.B2(n_744),
.Y(n_11837)
);

INVx1_ASAP7_75t_L g11838 ( 
.A(n_11154),
.Y(n_11838)
);

AOI21xp5_ASAP7_75t_L g11839 ( 
.A1(n_11408),
.A2(n_745),
.B(n_746),
.Y(n_11839)
);

NAND2xp5_ASAP7_75t_L g11840 ( 
.A(n_11082),
.B(n_746),
.Y(n_11840)
);

INVx3_ASAP7_75t_L g11841 ( 
.A(n_10905),
.Y(n_11841)
);

INVx2_ASAP7_75t_L g11842 ( 
.A(n_11163),
.Y(n_11842)
);

OAI22xp5_ASAP7_75t_L g11843 ( 
.A1(n_11079),
.A2(n_11241),
.B1(n_11395),
.B2(n_11388),
.Y(n_11843)
);

AO21x2_ASAP7_75t_L g11844 ( 
.A1(n_11097),
.A2(n_747),
.B(n_748),
.Y(n_11844)
);

NAND2xp5_ASAP7_75t_SL g11845 ( 
.A(n_10858),
.B(n_747),
.Y(n_11845)
);

OR2x2_ASAP7_75t_L g11846 ( 
.A(n_11284),
.B(n_750),
.Y(n_11846)
);

AOI21xp5_ASAP7_75t_L g11847 ( 
.A1(n_11415),
.A2(n_750),
.B(n_751),
.Y(n_11847)
);

AOI22x1_ASAP7_75t_L g11848 ( 
.A1(n_11139),
.A2(n_753),
.B1(n_751),
.B2(n_752),
.Y(n_11848)
);

INVx1_ASAP7_75t_L g11849 ( 
.A(n_11168),
.Y(n_11849)
);

INVx3_ASAP7_75t_L g11850 ( 
.A(n_10944),
.Y(n_11850)
);

NOR2xp33_ASAP7_75t_L g11851 ( 
.A(n_11115),
.B(n_752),
.Y(n_11851)
);

AOI21xp5_ASAP7_75t_L g11852 ( 
.A1(n_11428),
.A2(n_753),
.B(n_754),
.Y(n_11852)
);

AOI21xp5_ASAP7_75t_L g11853 ( 
.A1(n_11434),
.A2(n_754),
.B(n_755),
.Y(n_11853)
);

INVx1_ASAP7_75t_L g11854 ( 
.A(n_11189),
.Y(n_11854)
);

OR2x6_ASAP7_75t_SL g11855 ( 
.A(n_11341),
.B(n_755),
.Y(n_11855)
);

AOI21xp5_ASAP7_75t_L g11856 ( 
.A1(n_11457),
.A2(n_756),
.B(n_757),
.Y(n_11856)
);

AOI21xp5_ASAP7_75t_L g11857 ( 
.A1(n_11462),
.A2(n_756),
.B(n_758),
.Y(n_11857)
);

OA22x2_ASAP7_75t_L g11858 ( 
.A1(n_11042),
.A2(n_760),
.B1(n_758),
.B2(n_759),
.Y(n_11858)
);

NOR2xp33_ASAP7_75t_L g11859 ( 
.A(n_11336),
.B(n_11348),
.Y(n_11859)
);

A2O1A1Ixp33_ASAP7_75t_L g11860 ( 
.A1(n_10854),
.A2(n_762),
.B(n_760),
.C(n_761),
.Y(n_11860)
);

NAND2xp5_ASAP7_75t_SL g11861 ( 
.A(n_11386),
.B(n_762),
.Y(n_11861)
);

NAND2xp5_ASAP7_75t_SL g11862 ( 
.A(n_11464),
.B(n_763),
.Y(n_11862)
);

O2A1O1Ixp33_ASAP7_75t_SL g11863 ( 
.A1(n_11353),
.A2(n_10983),
.B(n_10977),
.C(n_10995),
.Y(n_11863)
);

O2A1O1Ixp33_ASAP7_75t_SL g11864 ( 
.A1(n_11002),
.A2(n_765),
.B(n_763),
.C(n_764),
.Y(n_11864)
);

AOI21xp5_ASAP7_75t_L g11865 ( 
.A1(n_11468),
.A2(n_765),
.B(n_766),
.Y(n_11865)
);

AOI21xp5_ASAP7_75t_L g11866 ( 
.A1(n_11481),
.A2(n_766),
.B(n_767),
.Y(n_11866)
);

A2O1A1Ixp33_ASAP7_75t_L g11867 ( 
.A1(n_11355),
.A2(n_770),
.B(n_768),
.C(n_769),
.Y(n_11867)
);

AOI21xp5_ASAP7_75t_L g11868 ( 
.A1(n_11533),
.A2(n_770),
.B(n_771),
.Y(n_11868)
);

AND2x4_ASAP7_75t_L g11869 ( 
.A(n_11107),
.B(n_772),
.Y(n_11869)
);

NAND2xp5_ASAP7_75t_L g11870 ( 
.A(n_11114),
.B(n_772),
.Y(n_11870)
);

AOI21xp5_ASAP7_75t_L g11871 ( 
.A1(n_11547),
.A2(n_773),
.B(n_774),
.Y(n_11871)
);

OR2x6_ASAP7_75t_L g11872 ( 
.A(n_11079),
.B(n_774),
.Y(n_11872)
);

O2A1O1Ixp33_ASAP7_75t_L g11873 ( 
.A1(n_11433),
.A2(n_777),
.B(n_775),
.C(n_776),
.Y(n_11873)
);

AOI21xp33_ASAP7_75t_L g11874 ( 
.A1(n_11442),
.A2(n_775),
.B(n_776),
.Y(n_11874)
);

BUFx6f_ASAP7_75t_L g11875 ( 
.A(n_10944),
.Y(n_11875)
);

NAND2x1p5_ASAP7_75t_L g11876 ( 
.A(n_11447),
.B(n_11149),
.Y(n_11876)
);

NOR2xp33_ASAP7_75t_L g11877 ( 
.A(n_11336),
.B(n_777),
.Y(n_11877)
);

NAND2xp5_ASAP7_75t_SL g11878 ( 
.A(n_11423),
.B(n_778),
.Y(n_11878)
);

INVx1_ASAP7_75t_L g11879 ( 
.A(n_11230),
.Y(n_11879)
);

INVxp33_ASAP7_75t_L g11880 ( 
.A(n_11127),
.Y(n_11880)
);

OAI22xp5_ASAP7_75t_SL g11881 ( 
.A1(n_11314),
.A2(n_780),
.B1(n_778),
.B2(n_779),
.Y(n_11881)
);

INVx1_ASAP7_75t_L g11882 ( 
.A(n_11252),
.Y(n_11882)
);

OAI22xp5_ASAP7_75t_L g11883 ( 
.A1(n_11241),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_11883)
);

OAI22x1_ASAP7_75t_L g11884 ( 
.A1(n_11356),
.A2(n_784),
.B1(n_782),
.B2(n_783),
.Y(n_11884)
);

OAI22xp5_ASAP7_75t_L g11885 ( 
.A1(n_11491),
.A2(n_785),
.B1(n_782),
.B2(n_784),
.Y(n_11885)
);

AOI21xp5_ASAP7_75t_L g11886 ( 
.A1(n_11551),
.A2(n_786),
.B(n_787),
.Y(n_11886)
);

BUFx3_ASAP7_75t_L g11887 ( 
.A(n_11513),
.Y(n_11887)
);

AOI21xp5_ASAP7_75t_L g11888 ( 
.A1(n_11563),
.A2(n_786),
.B(n_787),
.Y(n_11888)
);

O2A1O1Ixp5_ASAP7_75t_L g11889 ( 
.A1(n_11167),
.A2(n_791),
.B(n_788),
.C(n_789),
.Y(n_11889)
);

OAI21xp5_ASAP7_75t_L g11890 ( 
.A1(n_10824),
.A2(n_788),
.B(n_789),
.Y(n_11890)
);

NAND2xp5_ASAP7_75t_L g11891 ( 
.A(n_11425),
.B(n_791),
.Y(n_11891)
);

NOR2xp33_ASAP7_75t_L g11892 ( 
.A(n_11336),
.B(n_792),
.Y(n_11892)
);

AOI21xp5_ASAP7_75t_L g11893 ( 
.A1(n_11566),
.A2(n_792),
.B(n_793),
.Y(n_11893)
);

AOI33xp33_ASAP7_75t_L g11894 ( 
.A1(n_10877),
.A2(n_11191),
.A3(n_11328),
.B1(n_10893),
.B2(n_11238),
.B3(n_11316),
.Y(n_11894)
);

OAI22xp5_ASAP7_75t_L g11895 ( 
.A1(n_11505),
.A2(n_795),
.B1(n_793),
.B2(n_794),
.Y(n_11895)
);

BUFx8_ASAP7_75t_L g11896 ( 
.A(n_11499),
.Y(n_11896)
);

INVx2_ASAP7_75t_L g11897 ( 
.A(n_11256),
.Y(n_11897)
);

NAND2xp5_ASAP7_75t_L g11898 ( 
.A(n_11443),
.B(n_794),
.Y(n_11898)
);

NOR2xp33_ASAP7_75t_L g11899 ( 
.A(n_11348),
.B(n_795),
.Y(n_11899)
);

INVx4_ASAP7_75t_L g11900 ( 
.A(n_10944),
.Y(n_11900)
);

OR2x6_ASAP7_75t_L g11901 ( 
.A(n_11315),
.B(n_797),
.Y(n_11901)
);

NOR2xp33_ASAP7_75t_L g11902 ( 
.A(n_11348),
.B(n_797),
.Y(n_11902)
);

A2O1A1Ixp33_ASAP7_75t_L g11903 ( 
.A1(n_11359),
.A2(n_800),
.B(n_798),
.C(n_799),
.Y(n_11903)
);

NAND3xp33_ASAP7_75t_L g11904 ( 
.A(n_11173),
.B(n_798),
.C(n_799),
.Y(n_11904)
);

AOI22xp33_ASAP7_75t_L g11905 ( 
.A1(n_11535),
.A2(n_803),
.B1(n_801),
.B2(n_802),
.Y(n_11905)
);

OR2x6_ASAP7_75t_L g11906 ( 
.A(n_11321),
.B(n_801),
.Y(n_11906)
);

NAND2xp5_ASAP7_75t_SL g11907 ( 
.A(n_11431),
.B(n_802),
.Y(n_11907)
);

NAND2x1p5_ASAP7_75t_L g11908 ( 
.A(n_11196),
.B(n_803),
.Y(n_11908)
);

A2O1A1Ixp33_ASAP7_75t_L g11909 ( 
.A1(n_11371),
.A2(n_806),
.B(n_804),
.C(n_805),
.Y(n_11909)
);

AOI21xp5_ASAP7_75t_L g11910 ( 
.A1(n_11568),
.A2(n_804),
.B(n_805),
.Y(n_11910)
);

OAI22xp5_ASAP7_75t_SL g11911 ( 
.A1(n_11292),
.A2(n_808),
.B1(n_806),
.B2(n_807),
.Y(n_11911)
);

INVx3_ASAP7_75t_L g11912 ( 
.A(n_11460),
.Y(n_11912)
);

NAND2xp5_ASAP7_75t_L g11913 ( 
.A(n_11452),
.B(n_807),
.Y(n_11913)
);

AOI22xp33_ASAP7_75t_L g11914 ( 
.A1(n_11548),
.A2(n_10940),
.B1(n_11109),
.B2(n_11283),
.Y(n_11914)
);

BUFx6f_ASAP7_75t_L g11915 ( 
.A(n_11460),
.Y(n_11915)
);

INVx3_ASAP7_75t_SL g11916 ( 
.A(n_11127),
.Y(n_11916)
);

CKINVDCx10_ASAP7_75t_R g11917 ( 
.A(n_11526),
.Y(n_11917)
);

AOI21xp5_ASAP7_75t_L g11918 ( 
.A1(n_11103),
.A2(n_808),
.B(n_809),
.Y(n_11918)
);

NAND2xp5_ASAP7_75t_L g11919 ( 
.A(n_11454),
.B(n_809),
.Y(n_11919)
);

INVx1_ASAP7_75t_L g11920 ( 
.A(n_11410),
.Y(n_11920)
);

AOI21xp5_ASAP7_75t_L g11921 ( 
.A1(n_11382),
.A2(n_810),
.B(n_811),
.Y(n_11921)
);

A2O1A1Ixp33_ASAP7_75t_SL g11922 ( 
.A1(n_11174),
.A2(n_812),
.B(n_810),
.C(n_811),
.Y(n_11922)
);

AO21x1_ASAP7_75t_L g11923 ( 
.A1(n_11374),
.A2(n_813),
.B(n_814),
.Y(n_11923)
);

INVxp33_ASAP7_75t_SL g11924 ( 
.A(n_11199),
.Y(n_11924)
);

AOI21xp5_ASAP7_75t_L g11925 ( 
.A1(n_11393),
.A2(n_813),
.B(n_814),
.Y(n_11925)
);

AOI21xp5_ASAP7_75t_L g11926 ( 
.A1(n_11402),
.A2(n_815),
.B(n_816),
.Y(n_11926)
);

O2A1O1Ixp33_ASAP7_75t_L g11927 ( 
.A1(n_11038),
.A2(n_817),
.B(n_815),
.C(n_816),
.Y(n_11927)
);

O2A1O1Ixp33_ASAP7_75t_L g11928 ( 
.A1(n_11169),
.A2(n_819),
.B(n_817),
.C(n_818),
.Y(n_11928)
);

NOR2xp33_ASAP7_75t_L g11929 ( 
.A(n_11346),
.B(n_818),
.Y(n_11929)
);

INVx1_ASAP7_75t_L g11930 ( 
.A(n_11414),
.Y(n_11930)
);

NAND2xp5_ASAP7_75t_SL g11931 ( 
.A(n_11127),
.B(n_819),
.Y(n_11931)
);

AOI21xp5_ASAP7_75t_L g11932 ( 
.A1(n_11403),
.A2(n_820),
.B(n_821),
.Y(n_11932)
);

NAND2xp5_ASAP7_75t_L g11933 ( 
.A(n_11474),
.B(n_820),
.Y(n_11933)
);

NAND2xp5_ASAP7_75t_L g11934 ( 
.A(n_11510),
.B(n_821),
.Y(n_11934)
);

AOI21xp5_ASAP7_75t_L g11935 ( 
.A1(n_11404),
.A2(n_822),
.B(n_823),
.Y(n_11935)
);

INVx1_ASAP7_75t_L g11936 ( 
.A(n_11420),
.Y(n_11936)
);

HB1xp67_ASAP7_75t_L g11937 ( 
.A(n_11441),
.Y(n_11937)
);

AOI22xp5_ASAP7_75t_L g11938 ( 
.A1(n_11056),
.A2(n_11081),
.B1(n_11141),
.B2(n_11093),
.Y(n_11938)
);

NAND2xp5_ASAP7_75t_SL g11939 ( 
.A(n_11049),
.B(n_822),
.Y(n_11939)
);

INVx1_ASAP7_75t_L g11940 ( 
.A(n_11445),
.Y(n_11940)
);

NAND2xp5_ASAP7_75t_L g11941 ( 
.A(n_11532),
.B(n_823),
.Y(n_11941)
);

AOI22xp5_ASAP7_75t_L g11942 ( 
.A1(n_10902),
.A2(n_826),
.B1(n_824),
.B2(n_825),
.Y(n_11942)
);

NOR2x1_ASAP7_75t_L g11943 ( 
.A(n_11270),
.B(n_824),
.Y(n_11943)
);

NAND2xp5_ASAP7_75t_L g11944 ( 
.A(n_11542),
.B(n_827),
.Y(n_11944)
);

INVx2_ASAP7_75t_L g11945 ( 
.A(n_11458),
.Y(n_11945)
);

CKINVDCx5p33_ASAP7_75t_R g11946 ( 
.A(n_10963),
.Y(n_11946)
);

AND2x4_ASAP7_75t_L g11947 ( 
.A(n_11544),
.B(n_827),
.Y(n_11947)
);

INVx1_ASAP7_75t_L g11948 ( 
.A(n_11472),
.Y(n_11948)
);

A2O1A1Ixp33_ASAP7_75t_SL g11949 ( 
.A1(n_11193),
.A2(n_830),
.B(n_828),
.C(n_829),
.Y(n_11949)
);

AOI21x1_ASAP7_75t_L g11950 ( 
.A1(n_11262),
.A2(n_828),
.B(n_829),
.Y(n_11950)
);

INVx1_ASAP7_75t_L g11951 ( 
.A(n_11495),
.Y(n_11951)
);

AOI22xp5_ASAP7_75t_L g11952 ( 
.A1(n_10886),
.A2(n_833),
.B1(n_831),
.B2(n_832),
.Y(n_11952)
);

NOR3xp33_ASAP7_75t_L g11953 ( 
.A(n_11209),
.B(n_831),
.C(n_832),
.Y(n_11953)
);

A2O1A1Ixp33_ASAP7_75t_L g11954 ( 
.A1(n_11290),
.A2(n_835),
.B(n_833),
.C(n_834),
.Y(n_11954)
);

OAI21xp33_ASAP7_75t_L g11955 ( 
.A1(n_10992),
.A2(n_834),
.B(n_835),
.Y(n_11955)
);

NAND2xp5_ASAP7_75t_L g11956 ( 
.A(n_11546),
.B(n_836),
.Y(n_11956)
);

NOR2xp33_ASAP7_75t_L g11957 ( 
.A(n_10871),
.B(n_10896),
.Y(n_11957)
);

O2A1O1Ixp33_ASAP7_75t_L g11958 ( 
.A1(n_11177),
.A2(n_11274),
.B(n_11344),
.C(n_11332),
.Y(n_11958)
);

AOI21xp5_ASAP7_75t_L g11959 ( 
.A1(n_11409),
.A2(n_836),
.B(n_837),
.Y(n_11959)
);

NOR2xp33_ASAP7_75t_L g11960 ( 
.A(n_11031),
.B(n_837),
.Y(n_11960)
);

BUFx8_ASAP7_75t_L g11961 ( 
.A(n_11301),
.Y(n_11961)
);

AOI21xp5_ASAP7_75t_L g11962 ( 
.A1(n_11416),
.A2(n_838),
.B(n_839),
.Y(n_11962)
);

NAND2xp5_ASAP7_75t_L g11963 ( 
.A(n_11560),
.B(n_840),
.Y(n_11963)
);

NOR2xp33_ASAP7_75t_L g11964 ( 
.A(n_11023),
.B(n_841),
.Y(n_11964)
);

OAI21xp5_ASAP7_75t_L g11965 ( 
.A1(n_11421),
.A2(n_841),
.B(n_842),
.Y(n_11965)
);

NAND2xp5_ASAP7_75t_L g11966 ( 
.A(n_11564),
.B(n_842),
.Y(n_11966)
);

AOI21xp5_ASAP7_75t_L g11967 ( 
.A1(n_11422),
.A2(n_843),
.B(n_844),
.Y(n_11967)
);

A2O1A1Ixp33_ASAP7_75t_L g11968 ( 
.A1(n_11045),
.A2(n_11075),
.B(n_11094),
.C(n_11217),
.Y(n_11968)
);

AOI21xp5_ASAP7_75t_L g11969 ( 
.A1(n_11429),
.A2(n_843),
.B(n_844),
.Y(n_11969)
);

NAND2xp5_ASAP7_75t_SL g11970 ( 
.A(n_11309),
.B(n_845),
.Y(n_11970)
);

NAND2xp5_ASAP7_75t_L g11971 ( 
.A(n_11582),
.B(n_846),
.Y(n_11971)
);

NOR2xp33_ASAP7_75t_L g11972 ( 
.A(n_11242),
.B(n_846),
.Y(n_11972)
);

NOR2xp33_ASAP7_75t_L g11973 ( 
.A(n_11352),
.B(n_847),
.Y(n_11973)
);

O2A1O1Ixp33_ASAP7_75t_L g11974 ( 
.A1(n_11152),
.A2(n_849),
.B(n_847),
.C(n_848),
.Y(n_11974)
);

BUFx6f_ASAP7_75t_L g11975 ( 
.A(n_11460),
.Y(n_11975)
);

AOI21xp5_ASAP7_75t_L g11976 ( 
.A1(n_11432),
.A2(n_849),
.B(n_850),
.Y(n_11976)
);

BUFx6f_ASAP7_75t_L g11977 ( 
.A(n_11492),
.Y(n_11977)
);

NOR2xp33_ASAP7_75t_L g11978 ( 
.A(n_11326),
.B(n_850),
.Y(n_11978)
);

AOI21xp5_ASAP7_75t_L g11979 ( 
.A1(n_11436),
.A2(n_851),
.B(n_852),
.Y(n_11979)
);

AOI21x1_ASAP7_75t_L g11980 ( 
.A1(n_11322),
.A2(n_851),
.B(n_853),
.Y(n_11980)
);

AND2x4_ASAP7_75t_L g11981 ( 
.A(n_11597),
.B(n_853),
.Y(n_11981)
);

AOI21xp5_ASAP7_75t_L g11982 ( 
.A1(n_11437),
.A2(n_854),
.B(n_855),
.Y(n_11982)
);

NAND2xp5_ASAP7_75t_SL g11983 ( 
.A(n_11027),
.B(n_854),
.Y(n_11983)
);

OAI21x1_ASAP7_75t_L g11984 ( 
.A1(n_11522),
.A2(n_856),
.B(n_857),
.Y(n_11984)
);

NAND2xp5_ASAP7_75t_SL g11985 ( 
.A(n_11084),
.B(n_856),
.Y(n_11985)
);

INVx1_ASAP7_75t_L g11986 ( 
.A(n_11511),
.Y(n_11986)
);

AOI22xp33_ASAP7_75t_L g11987 ( 
.A1(n_11373),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.Y(n_11987)
);

NAND2xp5_ASAP7_75t_SL g11988 ( 
.A(n_11243),
.B(n_858),
.Y(n_11988)
);

INVx4_ASAP7_75t_L g11989 ( 
.A(n_11492),
.Y(n_11989)
);

AO21x1_ASAP7_75t_L g11990 ( 
.A1(n_11034),
.A2(n_11057),
.B(n_11305),
.Y(n_11990)
);

AOI21xp5_ASAP7_75t_L g11991 ( 
.A1(n_11470),
.A2(n_859),
.B(n_860),
.Y(n_11991)
);

NOR2xp67_ASAP7_75t_SL g11992 ( 
.A(n_11343),
.B(n_860),
.Y(n_11992)
);

NAND2xp5_ASAP7_75t_L g11993 ( 
.A(n_11126),
.B(n_861),
.Y(n_11993)
);

AOI21xp5_ASAP7_75t_L g11994 ( 
.A1(n_11473),
.A2(n_861),
.B(n_862),
.Y(n_11994)
);

AND2x2_ASAP7_75t_L g11995 ( 
.A(n_11514),
.B(n_11553),
.Y(n_11995)
);

OAI21x1_ASAP7_75t_L g11996 ( 
.A1(n_11142),
.A2(n_862),
.B(n_863),
.Y(n_11996)
);

O2A1O1Ixp33_ASAP7_75t_L g11997 ( 
.A1(n_11308),
.A2(n_865),
.B(n_863),
.C(n_864),
.Y(n_11997)
);

NAND2xp5_ASAP7_75t_SL g11998 ( 
.A(n_11181),
.B(n_865),
.Y(n_11998)
);

NOR2xp33_ASAP7_75t_L g11999 ( 
.A(n_11208),
.B(n_866),
.Y(n_11999)
);

NAND2xp5_ASAP7_75t_L g12000 ( 
.A(n_11133),
.B(n_866),
.Y(n_12000)
);

OA21x2_ASAP7_75t_L g12001 ( 
.A1(n_11222),
.A2(n_867),
.B(n_868),
.Y(n_12001)
);

INVx2_ASAP7_75t_L g12002 ( 
.A(n_11575),
.Y(n_12002)
);

INVx2_ASAP7_75t_L g12003 ( 
.A(n_11221),
.Y(n_12003)
);

INVx1_ASAP7_75t_L g12004 ( 
.A(n_11153),
.Y(n_12004)
);

NAND2xp5_ASAP7_75t_L g12005 ( 
.A(n_11146),
.B(n_867),
.Y(n_12005)
);

AND2x2_ASAP7_75t_L g12006 ( 
.A(n_11106),
.B(n_868),
.Y(n_12006)
);

A2O1A1Ixp33_ASAP7_75t_L g12007 ( 
.A1(n_10996),
.A2(n_871),
.B(n_869),
.C(n_870),
.Y(n_12007)
);

NAND2xp5_ASAP7_75t_L g12008 ( 
.A(n_11155),
.B(n_870),
.Y(n_12008)
);

AOI21xp5_ASAP7_75t_L g12009 ( 
.A1(n_11475),
.A2(n_871),
.B(n_873),
.Y(n_12009)
);

INVx3_ASAP7_75t_L g12010 ( 
.A(n_11492),
.Y(n_12010)
);

AOI21xp5_ASAP7_75t_L g12011 ( 
.A1(n_11477),
.A2(n_873),
.B(n_874),
.Y(n_12011)
);

NAND2xp5_ASAP7_75t_L g12012 ( 
.A(n_11161),
.B(n_875),
.Y(n_12012)
);

NAND2xp5_ASAP7_75t_SL g12013 ( 
.A(n_11022),
.B(n_875),
.Y(n_12013)
);

NAND2xp5_ASAP7_75t_L g12014 ( 
.A(n_11201),
.B(n_11216),
.Y(n_12014)
);

INVx3_ASAP7_75t_L g12015 ( 
.A(n_11531),
.Y(n_12015)
);

AOI21xp5_ASAP7_75t_L g12016 ( 
.A1(n_11487),
.A2(n_876),
.B(n_877),
.Y(n_12016)
);

NAND2xp5_ASAP7_75t_L g12017 ( 
.A(n_11259),
.B(n_876),
.Y(n_12017)
);

AOI21xp5_ASAP7_75t_L g12018 ( 
.A1(n_11494),
.A2(n_878),
.B(n_879),
.Y(n_12018)
);

INVx11_ASAP7_75t_L g12019 ( 
.A(n_11323),
.Y(n_12019)
);

OAI22xp5_ASAP7_75t_L g12020 ( 
.A1(n_11157),
.A2(n_881),
.B1(n_878),
.B2(n_880),
.Y(n_12020)
);

NOR3xp33_ASAP7_75t_L g12021 ( 
.A(n_11197),
.B(n_880),
.C(n_881),
.Y(n_12021)
);

NAND2xp5_ASAP7_75t_L g12022 ( 
.A(n_11384),
.B(n_882),
.Y(n_12022)
);

CKINVDCx10_ASAP7_75t_R g12023 ( 
.A(n_11376),
.Y(n_12023)
);

AOI21xp5_ASAP7_75t_L g12024 ( 
.A1(n_11507),
.A2(n_11515),
.B(n_11512),
.Y(n_12024)
);

NAND2xp5_ASAP7_75t_L g12025 ( 
.A(n_11405),
.B(n_882),
.Y(n_12025)
);

A2O1A1Ixp33_ASAP7_75t_L g12026 ( 
.A1(n_11294),
.A2(n_886),
.B(n_884),
.C(n_885),
.Y(n_12026)
);

HB1xp67_ASAP7_75t_L g12027 ( 
.A(n_11263),
.Y(n_12027)
);

NAND2xp5_ASAP7_75t_L g12028 ( 
.A(n_11407),
.B(n_884),
.Y(n_12028)
);

A2O1A1Ixp33_ASAP7_75t_SL g12029 ( 
.A1(n_11117),
.A2(n_887),
.B(n_885),
.C(n_886),
.Y(n_12029)
);

NAND2xp5_ASAP7_75t_L g12030 ( 
.A(n_11411),
.B(n_888),
.Y(n_12030)
);

AOI21xp5_ASAP7_75t_L g12031 ( 
.A1(n_11516),
.A2(n_888),
.B(n_889),
.Y(n_12031)
);

AOI21xp5_ASAP7_75t_L g12032 ( 
.A1(n_11519),
.A2(n_889),
.B(n_890),
.Y(n_12032)
);

NAND2xp5_ASAP7_75t_L g12033 ( 
.A(n_11417),
.B(n_11435),
.Y(n_12033)
);

OAI22xp5_ASAP7_75t_L g12034 ( 
.A1(n_11331),
.A2(n_892),
.B1(n_890),
.B2(n_891),
.Y(n_12034)
);

AOI21xp5_ASAP7_75t_L g12035 ( 
.A1(n_11521),
.A2(n_891),
.B(n_892),
.Y(n_12035)
);

BUFx2_ASAP7_75t_L g12036 ( 
.A(n_11240),
.Y(n_12036)
);

A2O1A1Ixp33_ASAP7_75t_L g12037 ( 
.A1(n_11300),
.A2(n_895),
.B(n_893),
.C(n_894),
.Y(n_12037)
);

NAND2xp5_ASAP7_75t_L g12038 ( 
.A(n_11453),
.B(n_893),
.Y(n_12038)
);

OAI21xp5_ASAP7_75t_L g12039 ( 
.A1(n_11524),
.A2(n_895),
.B(n_896),
.Y(n_12039)
);

NOR2xp33_ASAP7_75t_L g12040 ( 
.A(n_10997),
.B(n_896),
.Y(n_12040)
);

AND2x2_ASAP7_75t_L g12041 ( 
.A(n_11226),
.B(n_897),
.Y(n_12041)
);

AOI222xp33_ASAP7_75t_L g12042 ( 
.A1(n_11299),
.A2(n_900),
.B1(n_902),
.B2(n_898),
.C1(n_899),
.C2(n_901),
.Y(n_12042)
);

AND2x4_ASAP7_75t_L g12043 ( 
.A(n_11008),
.B(n_898),
.Y(n_12043)
);

OAI22xp5_ASAP7_75t_L g12044 ( 
.A1(n_11354),
.A2(n_901),
.B1(n_899),
.B2(n_900),
.Y(n_12044)
);

A2O1A1Ixp33_ASAP7_75t_L g12045 ( 
.A1(n_11040),
.A2(n_904),
.B(n_902),
.C(n_903),
.Y(n_12045)
);

AOI22xp5_ASAP7_75t_L g12046 ( 
.A1(n_10895),
.A2(n_906),
.B1(n_903),
.B2(n_905),
.Y(n_12046)
);

NAND2xp5_ASAP7_75t_L g12047 ( 
.A(n_11461),
.B(n_905),
.Y(n_12047)
);

O2A1O1Ixp5_ASAP7_75t_L g12048 ( 
.A1(n_11364),
.A2(n_909),
.B(n_907),
.C(n_908),
.Y(n_12048)
);

OAI21xp5_ASAP7_75t_L g12049 ( 
.A1(n_11536),
.A2(n_908),
.B(n_909),
.Y(n_12049)
);

NAND2xp5_ASAP7_75t_L g12050 ( 
.A(n_11465),
.B(n_910),
.Y(n_12050)
);

AOI21x1_ASAP7_75t_L g12051 ( 
.A1(n_10929),
.A2(n_911),
.B(n_912),
.Y(n_12051)
);

INVx3_ASAP7_75t_L g12052 ( 
.A(n_11531),
.Y(n_12052)
);

INVx1_ASAP7_75t_L g12053 ( 
.A(n_11258),
.Y(n_12053)
);

AOI21xp5_ASAP7_75t_L g12054 ( 
.A1(n_11538),
.A2(n_911),
.B(n_912),
.Y(n_12054)
);

BUFx3_ASAP7_75t_L g12055 ( 
.A(n_11531),
.Y(n_12055)
);

INVx1_ASAP7_75t_L g12056 ( 
.A(n_11236),
.Y(n_12056)
);

O2A1O1Ixp33_ASAP7_75t_L g12057 ( 
.A1(n_11185),
.A2(n_915),
.B(n_913),
.C(n_914),
.Y(n_12057)
);

INVx2_ASAP7_75t_L g12058 ( 
.A(n_11116),
.Y(n_12058)
);

AOI21x1_ASAP7_75t_L g12059 ( 
.A1(n_11361),
.A2(n_914),
.B(n_915),
.Y(n_12059)
);

AOI21xp5_ASAP7_75t_L g12060 ( 
.A1(n_11543),
.A2(n_917),
.B(n_918),
.Y(n_12060)
);

INVx1_ASAP7_75t_L g12061 ( 
.A(n_11239),
.Y(n_12061)
);

NAND2xp33_ASAP7_75t_L g12062 ( 
.A(n_10846),
.B(n_917),
.Y(n_12062)
);

INVx2_ASAP7_75t_L g12063 ( 
.A(n_11121),
.Y(n_12063)
);

INVx2_ASAP7_75t_L g12064 ( 
.A(n_11125),
.Y(n_12064)
);

NOR2xp33_ASAP7_75t_L g12065 ( 
.A(n_11248),
.B(n_919),
.Y(n_12065)
);

AOI21xp5_ASAP7_75t_L g12066 ( 
.A1(n_11557),
.A2(n_919),
.B(n_920),
.Y(n_12066)
);

NAND2xp5_ASAP7_75t_SL g12067 ( 
.A(n_11304),
.B(n_920),
.Y(n_12067)
);

AOI22xp5_ASAP7_75t_L g12068 ( 
.A1(n_11175),
.A2(n_923),
.B1(n_921),
.B2(n_922),
.Y(n_12068)
);

AOI21xp5_ASAP7_75t_L g12069 ( 
.A1(n_11558),
.A2(n_922),
.B(n_924),
.Y(n_12069)
);

NAND2xp33_ASAP7_75t_L g12070 ( 
.A(n_10846),
.B(n_924),
.Y(n_12070)
);

AOI21xp5_ASAP7_75t_L g12071 ( 
.A1(n_11561),
.A2(n_925),
.B(n_926),
.Y(n_12071)
);

OAI22xp5_ASAP7_75t_L g12072 ( 
.A1(n_11345),
.A2(n_927),
.B1(n_925),
.B2(n_926),
.Y(n_12072)
);

A2O1A1Ixp33_ASAP7_75t_L g12073 ( 
.A1(n_11047),
.A2(n_929),
.B(n_927),
.C(n_928),
.Y(n_12073)
);

OAI22xp5_ASAP7_75t_L g12074 ( 
.A1(n_11349),
.A2(n_930),
.B1(n_928),
.B2(n_929),
.Y(n_12074)
);

BUFx6f_ASAP7_75t_L g12075 ( 
.A(n_11110),
.Y(n_12075)
);

NAND2xp5_ASAP7_75t_L g12076 ( 
.A(n_11466),
.B(n_930),
.Y(n_12076)
);

NAND2xp5_ASAP7_75t_SL g12077 ( 
.A(n_11311),
.B(n_931),
.Y(n_12077)
);

AOI21xp5_ASAP7_75t_L g12078 ( 
.A1(n_11569),
.A2(n_931),
.B(n_932),
.Y(n_12078)
);

NOR2xp33_ASAP7_75t_L g12079 ( 
.A(n_11278),
.B(n_932),
.Y(n_12079)
);

INVx2_ASAP7_75t_L g12080 ( 
.A(n_11131),
.Y(n_12080)
);

CKINVDCx8_ASAP7_75t_R g12081 ( 
.A(n_11134),
.Y(n_12081)
);

INVx2_ASAP7_75t_L g12082 ( 
.A(n_11140),
.Y(n_12082)
);

AOI21xp5_ASAP7_75t_L g12083 ( 
.A1(n_11572),
.A2(n_933),
.B(n_934),
.Y(n_12083)
);

O2A1O1Ixp33_ASAP7_75t_L g12084 ( 
.A1(n_10966),
.A2(n_936),
.B(n_934),
.C(n_935),
.Y(n_12084)
);

AND2x2_ASAP7_75t_L g12085 ( 
.A(n_11205),
.B(n_935),
.Y(n_12085)
);

AOI21xp5_ASAP7_75t_L g12086 ( 
.A1(n_11574),
.A2(n_936),
.B(n_937),
.Y(n_12086)
);

A2O1A1Ixp33_ASAP7_75t_L g12087 ( 
.A1(n_11052),
.A2(n_939),
.B(n_937),
.C(n_938),
.Y(n_12087)
);

INVx1_ASAP7_75t_L g12088 ( 
.A(n_11250),
.Y(n_12088)
);

NAND3xp33_ASAP7_75t_L g12089 ( 
.A(n_11366),
.B(n_938),
.C(n_939),
.Y(n_12089)
);

NAND2xp5_ASAP7_75t_L g12090 ( 
.A(n_11478),
.B(n_940),
.Y(n_12090)
);

A2O1A1Ixp33_ASAP7_75t_L g12091 ( 
.A1(n_11063),
.A2(n_11065),
.B(n_11066),
.C(n_11120),
.Y(n_12091)
);

NAND2xp5_ASAP7_75t_L g12092 ( 
.A(n_11483),
.B(n_940),
.Y(n_12092)
);

NAND2xp5_ASAP7_75t_L g12093 ( 
.A(n_11488),
.B(n_941),
.Y(n_12093)
);

NAND2xp5_ASAP7_75t_SL g12094 ( 
.A(n_11277),
.B(n_941),
.Y(n_12094)
);

INVx2_ASAP7_75t_L g12095 ( 
.A(n_11162),
.Y(n_12095)
);

OAI22xp5_ASAP7_75t_L g12096 ( 
.A1(n_11360),
.A2(n_11367),
.B1(n_11333),
.B2(n_11335),
.Y(n_12096)
);

NAND2xp5_ASAP7_75t_SL g12097 ( 
.A(n_11327),
.B(n_942),
.Y(n_12097)
);

INVx2_ASAP7_75t_L g12098 ( 
.A(n_11165),
.Y(n_12098)
);

O2A1O1Ixp33_ASAP7_75t_L g12099 ( 
.A1(n_11312),
.A2(n_944),
.B(n_942),
.C(n_943),
.Y(n_12099)
);

O2A1O1Ixp33_ASAP7_75t_L g12100 ( 
.A1(n_11426),
.A2(n_10941),
.B(n_11043),
.C(n_11375),
.Y(n_12100)
);

NOR2xp33_ASAP7_75t_L g12101 ( 
.A(n_11298),
.B(n_943),
.Y(n_12101)
);

BUFx6f_ASAP7_75t_L g12102 ( 
.A(n_11134),
.Y(n_12102)
);

NAND2xp5_ASAP7_75t_SL g12103 ( 
.A(n_11329),
.B(n_944),
.Y(n_12103)
);

CKINVDCx10_ASAP7_75t_R g12104 ( 
.A(n_11357),
.Y(n_12104)
);

OAI22xp5_ASAP7_75t_L g12105 ( 
.A1(n_11020),
.A2(n_11496),
.B1(n_11506),
.B2(n_11490),
.Y(n_12105)
);

INVx1_ASAP7_75t_L g12106 ( 
.A(n_11253),
.Y(n_12106)
);

BUFx2_ASAP7_75t_L g12107 ( 
.A(n_11240),
.Y(n_12107)
);

AND2x2_ASAP7_75t_L g12108 ( 
.A(n_11387),
.B(n_945),
.Y(n_12108)
);

NOR2xp33_ASAP7_75t_SL g12109 ( 
.A(n_11269),
.B(n_945),
.Y(n_12109)
);

NAND2xp5_ASAP7_75t_SL g12110 ( 
.A(n_11033),
.B(n_946),
.Y(n_12110)
);

AOI21xp5_ASAP7_75t_L g12111 ( 
.A1(n_11578),
.A2(n_946),
.B(n_947),
.Y(n_12111)
);

INVx2_ASAP7_75t_L g12112 ( 
.A(n_11170),
.Y(n_12112)
);

AND2x2_ASAP7_75t_L g12113 ( 
.A(n_11419),
.B(n_947),
.Y(n_12113)
);

AOI21xp5_ASAP7_75t_L g12114 ( 
.A1(n_11583),
.A2(n_948),
.B(n_949),
.Y(n_12114)
);

NOR2xp67_ASAP7_75t_L g12115 ( 
.A(n_11004),
.B(n_948),
.Y(n_12115)
);

AOI21xp5_ASAP7_75t_L g12116 ( 
.A1(n_11585),
.A2(n_949),
.B(n_950),
.Y(n_12116)
);

INVx1_ASAP7_75t_L g12117 ( 
.A(n_11254),
.Y(n_12117)
);

NAND2xp5_ASAP7_75t_L g12118 ( 
.A(n_11509),
.B(n_950),
.Y(n_12118)
);

OAI21xp5_ASAP7_75t_L g12119 ( 
.A1(n_11588),
.A2(n_951),
.B(n_952),
.Y(n_12119)
);

OAI22xp5_ASAP7_75t_SL g12120 ( 
.A1(n_11036),
.A2(n_954),
.B1(n_952),
.B2(n_953),
.Y(n_12120)
);

AND2x2_ASAP7_75t_L g12121 ( 
.A(n_11446),
.B(n_953),
.Y(n_12121)
);

INVx1_ASAP7_75t_L g12122 ( 
.A(n_11171),
.Y(n_12122)
);

AOI21xp5_ASAP7_75t_L g12123 ( 
.A1(n_11589),
.A2(n_954),
.B(n_955),
.Y(n_12123)
);

AOI22xp33_ASAP7_75t_L g12124 ( 
.A1(n_11244),
.A2(n_11339),
.B1(n_11599),
.B2(n_10846),
.Y(n_12124)
);

OAI21xp33_ASAP7_75t_SL g12125 ( 
.A1(n_11188),
.A2(n_955),
.B(n_956),
.Y(n_12125)
);

AND2x6_ASAP7_75t_L g12126 ( 
.A(n_11240),
.B(n_956),
.Y(n_12126)
);

NAND2xp5_ASAP7_75t_L g12127 ( 
.A(n_11528),
.B(n_957),
.Y(n_12127)
);

NAND3xp33_ASAP7_75t_L g12128 ( 
.A(n_11122),
.B(n_957),
.C(n_958),
.Y(n_12128)
);

NOR2xp33_ASAP7_75t_L g12129 ( 
.A(n_11307),
.B(n_958),
.Y(n_12129)
);

AO21x1_ASAP7_75t_L g12130 ( 
.A1(n_11330),
.A2(n_959),
.B(n_960),
.Y(n_12130)
);

AOI21xp5_ASAP7_75t_L g12131 ( 
.A1(n_11592),
.A2(n_959),
.B(n_960),
.Y(n_12131)
);

INVx2_ASAP7_75t_L g12132 ( 
.A(n_11176),
.Y(n_12132)
);

INVxp67_ASAP7_75t_L g12133 ( 
.A(n_11144),
.Y(n_12133)
);

NAND2xp5_ASAP7_75t_L g12134 ( 
.A(n_11530),
.B(n_961),
.Y(n_12134)
);

NOR2xp33_ASAP7_75t_L g12135 ( 
.A(n_11545),
.B(n_962),
.Y(n_12135)
);

OAI321xp33_ASAP7_75t_L g12136 ( 
.A1(n_10873),
.A2(n_10885),
.A3(n_10849),
.B1(n_10838),
.B2(n_10933),
.C(n_11013),
.Y(n_12136)
);

INVx1_ASAP7_75t_SL g12137 ( 
.A(n_11265),
.Y(n_12137)
);

NAND2xp5_ASAP7_75t_L g12138 ( 
.A(n_11556),
.B(n_962),
.Y(n_12138)
);

NOR2xp33_ASAP7_75t_L g12139 ( 
.A(n_11562),
.B(n_11571),
.Y(n_12139)
);

NOR2xp33_ASAP7_75t_L g12140 ( 
.A(n_11576),
.B(n_963),
.Y(n_12140)
);

OAI21xp33_ASAP7_75t_L g12141 ( 
.A1(n_11039),
.A2(n_963),
.B(n_964),
.Y(n_12141)
);

NOR2xp33_ASAP7_75t_L g12142 ( 
.A(n_11577),
.B(n_965),
.Y(n_12142)
);

NAND2xp5_ASAP7_75t_SL g12143 ( 
.A(n_11158),
.B(n_965),
.Y(n_12143)
);

INVx1_ASAP7_75t_L g12144 ( 
.A(n_11178),
.Y(n_12144)
);

NAND2xp5_ASAP7_75t_SL g12145 ( 
.A(n_11291),
.B(n_966),
.Y(n_12145)
);

OAI22xp5_ASAP7_75t_L g12146 ( 
.A1(n_11580),
.A2(n_968),
.B1(n_966),
.B2(n_967),
.Y(n_12146)
);

NAND2xp5_ASAP7_75t_L g12147 ( 
.A(n_11581),
.B(n_967),
.Y(n_12147)
);

NAND2xp5_ASAP7_75t_SL g12148 ( 
.A(n_11586),
.B(n_968),
.Y(n_12148)
);

CKINVDCx10_ASAP7_75t_R g12149 ( 
.A(n_11379),
.Y(n_12149)
);

NAND2xp5_ASAP7_75t_L g12150 ( 
.A(n_11591),
.B(n_969),
.Y(n_12150)
);

NAND2xp5_ASAP7_75t_L g12151 ( 
.A(n_11593),
.B(n_970),
.Y(n_12151)
);

NAND2xp5_ASAP7_75t_L g12152 ( 
.A(n_11602),
.B(n_970),
.Y(n_12152)
);

NAND2xp5_ASAP7_75t_L g12153 ( 
.A(n_10923),
.B(n_10927),
.Y(n_12153)
);

INVx1_ASAP7_75t_L g12154 ( 
.A(n_11180),
.Y(n_12154)
);

NAND2xp5_ASAP7_75t_L g12155 ( 
.A(n_10936),
.B(n_971),
.Y(n_12155)
);

NAND2xp5_ASAP7_75t_L g12156 ( 
.A(n_10937),
.B(n_971),
.Y(n_12156)
);

INVx2_ASAP7_75t_L g12157 ( 
.A(n_11182),
.Y(n_12157)
);

NAND2xp5_ASAP7_75t_L g12158 ( 
.A(n_10943),
.B(n_972),
.Y(n_12158)
);

NOR2xp33_ASAP7_75t_SL g12159 ( 
.A(n_11124),
.B(n_972),
.Y(n_12159)
);

AND2x4_ASAP7_75t_L g12160 ( 
.A(n_10848),
.B(n_973),
.Y(n_12160)
);

BUFx2_ASAP7_75t_L g12161 ( 
.A(n_11134),
.Y(n_12161)
);

AOI21xp5_ASAP7_75t_L g12162 ( 
.A1(n_11596),
.A2(n_973),
.B(n_974),
.Y(n_12162)
);

NOR2xp33_ASAP7_75t_L g12163 ( 
.A(n_11338),
.B(n_974),
.Y(n_12163)
);

NAND2xp5_ASAP7_75t_L g12164 ( 
.A(n_10974),
.B(n_975),
.Y(n_12164)
);

INVx1_ASAP7_75t_L g12165 ( 
.A(n_11183),
.Y(n_12165)
);

AOI21xp5_ASAP7_75t_L g12166 ( 
.A1(n_11603),
.A2(n_975),
.B(n_976),
.Y(n_12166)
);

O2A1O1Ixp5_ASAP7_75t_L g12167 ( 
.A1(n_11118),
.A2(n_978),
.B(n_976),
.C(n_977),
.Y(n_12167)
);

AOI22xp33_ASAP7_75t_L g12168 ( 
.A1(n_10846),
.A2(n_980),
.B1(n_978),
.B2(n_979),
.Y(n_12168)
);

OR2x6_ASAP7_75t_L g12169 ( 
.A(n_10909),
.B(n_980),
.Y(n_12169)
);

NAND2xp5_ASAP7_75t_L g12170 ( 
.A(n_10985),
.B(n_981),
.Y(n_12170)
);

AOI22xp33_ASAP7_75t_L g12171 ( 
.A1(n_11599),
.A2(n_983),
.B1(n_981),
.B2(n_982),
.Y(n_12171)
);

INVxp67_ASAP7_75t_L g12172 ( 
.A(n_11130),
.Y(n_12172)
);

AO21x1_ASAP7_75t_L g12173 ( 
.A1(n_10894),
.A2(n_982),
.B(n_983),
.Y(n_12173)
);

NOR2xp33_ASAP7_75t_L g12174 ( 
.A(n_11378),
.B(n_984),
.Y(n_12174)
);

AOI22xp5_ASAP7_75t_L g12175 ( 
.A1(n_11599),
.A2(n_986),
.B1(n_984),
.B2(n_985),
.Y(n_12175)
);

NOR2xp33_ASAP7_75t_L g12176 ( 
.A(n_11449),
.B(n_985),
.Y(n_12176)
);

INVx2_ASAP7_75t_L g12177 ( 
.A(n_11219),
.Y(n_12177)
);

OR2x6_ASAP7_75t_L g12178 ( 
.A(n_11590),
.B(n_987),
.Y(n_12178)
);

OAI22xp5_ASAP7_75t_L g12179 ( 
.A1(n_11062),
.A2(n_989),
.B1(n_987),
.B2(n_988),
.Y(n_12179)
);

NOR3xp33_ASAP7_75t_L g12180 ( 
.A(n_11286),
.B(n_988),
.C(n_989),
.Y(n_12180)
);

NAND2xp5_ASAP7_75t_SL g12181 ( 
.A(n_11215),
.B(n_990),
.Y(n_12181)
);

A2O1A1Ixp33_ASAP7_75t_L g12182 ( 
.A1(n_11101),
.A2(n_993),
.B(n_991),
.C(n_992),
.Y(n_12182)
);

AND2x4_ASAP7_75t_L g12183 ( 
.A(n_11390),
.B(n_991),
.Y(n_12183)
);

AOI21xp5_ASAP7_75t_L g12184 ( 
.A1(n_11150),
.A2(n_11232),
.B(n_11001),
.Y(n_12184)
);

AOI21xp5_ASAP7_75t_L g12185 ( 
.A1(n_10999),
.A2(n_992),
.B(n_993),
.Y(n_12185)
);

BUFx12f_ASAP7_75t_L g12186 ( 
.A(n_11025),
.Y(n_12186)
);

AND2x2_ASAP7_75t_L g12187 ( 
.A(n_11456),
.B(n_994),
.Y(n_12187)
);

INVx2_ASAP7_75t_L g12188 ( 
.A(n_11223),
.Y(n_12188)
);

NAND2xp5_ASAP7_75t_SL g12189 ( 
.A(n_11295),
.B(n_994),
.Y(n_12189)
);

AO32x2_ASAP7_75t_L g12190 ( 
.A1(n_11228),
.A2(n_997),
.A3(n_995),
.B1(n_996),
.B2(n_998),
.Y(n_12190)
);

NAND2x1p5_ASAP7_75t_L g12191 ( 
.A(n_11145),
.B(n_11044),
.Y(n_12191)
);

NAND2xp5_ASAP7_75t_L g12192 ( 
.A(n_11000),
.B(n_995),
.Y(n_12192)
);

AOI21xp5_ASAP7_75t_L g12193 ( 
.A1(n_10860),
.A2(n_996),
.B(n_998),
.Y(n_12193)
);

BUFx8_ASAP7_75t_L g12194 ( 
.A(n_10901),
.Y(n_12194)
);

NAND2xp5_ASAP7_75t_L g12195 ( 
.A(n_10958),
.B(n_999),
.Y(n_12195)
);

NAND2xp5_ASAP7_75t_L g12196 ( 
.A(n_10971),
.B(n_999),
.Y(n_12196)
);

NOR2xp33_ASAP7_75t_L g12197 ( 
.A(n_11486),
.B(n_1000),
.Y(n_12197)
);

AOI21xp5_ASAP7_75t_L g12198 ( 
.A1(n_10861),
.A2(n_10868),
.B(n_10862),
.Y(n_12198)
);

NAND2xp5_ASAP7_75t_SL g12199 ( 
.A(n_11288),
.B(n_1000),
.Y(n_12199)
);

AOI22xp5_ASAP7_75t_L g12200 ( 
.A1(n_11599),
.A2(n_10864),
.B1(n_10900),
.B2(n_10850),
.Y(n_12200)
);

NAND2xp5_ASAP7_75t_SL g12201 ( 
.A(n_11337),
.B(n_1001),
.Y(n_12201)
);

NAND2xp5_ASAP7_75t_L g12202 ( 
.A(n_10973),
.B(n_1001),
.Y(n_12202)
);

AOI21xp5_ASAP7_75t_L g12203 ( 
.A1(n_10869),
.A2(n_10876),
.B(n_10874),
.Y(n_12203)
);

O2A1O1Ixp33_ASAP7_75t_SL g12204 ( 
.A1(n_11069),
.A2(n_1004),
.B(n_1002),
.C(n_1003),
.Y(n_12204)
);

AND2x2_ASAP7_75t_L g12205 ( 
.A(n_11541),
.B(n_1002),
.Y(n_12205)
);

NAND2xp5_ASAP7_75t_L g12206 ( 
.A(n_10827),
.B(n_1003),
.Y(n_12206)
);

INVx2_ASAP7_75t_L g12207 ( 
.A(n_11164),
.Y(n_12207)
);

BUFx2_ASAP7_75t_L g12208 ( 
.A(n_11029),
.Y(n_12208)
);

NOR2xp33_ASAP7_75t_L g12209 ( 
.A(n_11035),
.B(n_1005),
.Y(n_12209)
);

OAI22x1_ASAP7_75t_L g12210 ( 
.A1(n_11540),
.A2(n_1007),
.B1(n_1005),
.B2(n_1006),
.Y(n_12210)
);

AOI21xp5_ASAP7_75t_L g12211 ( 
.A1(n_10883),
.A2(n_1006),
.B(n_1007),
.Y(n_12211)
);

NAND2xp5_ASAP7_75t_L g12212 ( 
.A(n_10830),
.B(n_1008),
.Y(n_12212)
);

NAND2xp5_ASAP7_75t_SL g12213 ( 
.A(n_11340),
.B(n_1009),
.Y(n_12213)
);

AOI21xp5_ASAP7_75t_L g12214 ( 
.A1(n_10888),
.A2(n_1009),
.B(n_1010),
.Y(n_12214)
);

NAND2xp5_ASAP7_75t_L g12215 ( 
.A(n_10841),
.B(n_1010),
.Y(n_12215)
);

AOI21xp5_ASAP7_75t_L g12216 ( 
.A1(n_10889),
.A2(n_10897),
.B(n_10890),
.Y(n_12216)
);

AOI21xp5_ASAP7_75t_L g12217 ( 
.A1(n_10906),
.A2(n_1011),
.B(n_1012),
.Y(n_12217)
);

AO21x1_ASAP7_75t_L g12218 ( 
.A1(n_11071),
.A2(n_11074),
.B(n_11072),
.Y(n_12218)
);

NOR2xp33_ASAP7_75t_L g12219 ( 
.A(n_11080),
.B(n_1013),
.Y(n_12219)
);

NAND2xp5_ASAP7_75t_L g12220 ( 
.A(n_10844),
.B(n_1013),
.Y(n_12220)
);

OAI22xp5_ASAP7_75t_L g12221 ( 
.A1(n_11083),
.A2(n_1016),
.B1(n_1014),
.B2(n_1015),
.Y(n_12221)
);

HB1xp67_ASAP7_75t_L g12222 ( 
.A(n_11227),
.Y(n_12222)
);

AOI21xp5_ASAP7_75t_L g12223 ( 
.A1(n_10910),
.A2(n_1014),
.B(n_1015),
.Y(n_12223)
);

INVx2_ASAP7_75t_L g12224 ( 
.A(n_11234),
.Y(n_12224)
);

AO32x2_ASAP7_75t_L g12225 ( 
.A1(n_11296),
.A2(n_1018),
.A3(n_1016),
.B1(n_1017),
.B2(n_1019),
.Y(n_12225)
);

NAND2xp5_ASAP7_75t_SL g12226 ( 
.A(n_11350),
.B(n_1017),
.Y(n_12226)
);

NAND2xp5_ASAP7_75t_SL g12227 ( 
.A(n_10987),
.B(n_1019),
.Y(n_12227)
);

INVx2_ASAP7_75t_SL g12228 ( 
.A(n_11508),
.Y(n_12228)
);

O2A1O1Ixp33_ASAP7_75t_L g12229 ( 
.A1(n_11098),
.A2(n_11267),
.B(n_11268),
.C(n_11324),
.Y(n_12229)
);

NAND2xp5_ASAP7_75t_L g12230 ( 
.A(n_10845),
.B(n_10863),
.Y(n_12230)
);

NOR2xp67_ASAP7_75t_SL g12231 ( 
.A(n_11129),
.B(n_1020),
.Y(n_12231)
);

AO21x1_ASAP7_75t_L g12232 ( 
.A1(n_10865),
.A2(n_10882),
.B(n_10867),
.Y(n_12232)
);

AOI21xp5_ASAP7_75t_L g12233 ( 
.A1(n_10913),
.A2(n_1020),
.B(n_1021),
.Y(n_12233)
);

AOI21xp5_ASAP7_75t_L g12234 ( 
.A1(n_10918),
.A2(n_1021),
.B(n_1022),
.Y(n_12234)
);

HB1xp67_ASAP7_75t_L g12235 ( 
.A(n_11282),
.Y(n_12235)
);

NAND2xp5_ASAP7_75t_SL g12236 ( 
.A(n_11032),
.B(n_1022),
.Y(n_12236)
);

BUFx8_ASAP7_75t_L g12237 ( 
.A(n_11210),
.Y(n_12237)
);

NAND2xp5_ASAP7_75t_L g12238 ( 
.A(n_10898),
.B(n_1023),
.Y(n_12238)
);

NAND2xp5_ASAP7_75t_L g12239 ( 
.A(n_10899),
.B(n_1023),
.Y(n_12239)
);

NOR2xp33_ASAP7_75t_L g12240 ( 
.A(n_11293),
.B(n_1024),
.Y(n_12240)
);

OAI22xp5_ASAP7_75t_L g12241 ( 
.A1(n_10914),
.A2(n_1026),
.B1(n_1024),
.B2(n_1025),
.Y(n_12241)
);

NOR2xp33_ASAP7_75t_L g12242 ( 
.A(n_11297),
.B(n_1025),
.Y(n_12242)
);

NAND2xp5_ASAP7_75t_L g12243 ( 
.A(n_10921),
.B(n_1027),
.Y(n_12243)
);

INVx3_ASAP7_75t_L g12244 ( 
.A(n_11529),
.Y(n_12244)
);

NAND2xp5_ASAP7_75t_L g12245 ( 
.A(n_11026),
.B(n_1028),
.Y(n_12245)
);

O2A1O1Ixp33_ASAP7_75t_L g12246 ( 
.A1(n_11090),
.A2(n_1030),
.B(n_1028),
.C(n_1029),
.Y(n_12246)
);

NOR2xp33_ASAP7_75t_SL g12247 ( 
.A(n_10857),
.B(n_1029),
.Y(n_12247)
);

NOR2xp33_ASAP7_75t_L g12248 ( 
.A(n_10908),
.B(n_1030),
.Y(n_12248)
);

OAI21xp5_ASAP7_75t_L g12249 ( 
.A1(n_10998),
.A2(n_1031),
.B(n_1032),
.Y(n_12249)
);

AND2x2_ASAP7_75t_L g12250 ( 
.A(n_11028),
.B(n_11030),
.Y(n_12250)
);

INVx1_ASAP7_75t_L g12251 ( 
.A(n_11427),
.Y(n_12251)
);

INVx2_ASAP7_75t_L g12252 ( 
.A(n_11276),
.Y(n_12252)
);

NOR2xp33_ASAP7_75t_L g12253 ( 
.A(n_11280),
.B(n_1031),
.Y(n_12253)
);

AOI21xp5_ASAP7_75t_L g12254 ( 
.A1(n_10922),
.A2(n_1032),
.B(n_1033),
.Y(n_12254)
);

NOR3xp33_ASAP7_75t_L g12255 ( 
.A(n_10976),
.B(n_1033),
.C(n_1034),
.Y(n_12255)
);

BUFx3_ASAP7_75t_L g12256 ( 
.A(n_11358),
.Y(n_12256)
);

AOI21xp5_ASAP7_75t_L g12257 ( 
.A1(n_10931),
.A2(n_1034),
.B(n_1035),
.Y(n_12257)
);

INVx1_ASAP7_75t_L g12258 ( 
.A(n_11427),
.Y(n_12258)
);

NOR2xp33_ASAP7_75t_R g12259 ( 
.A(n_10832),
.B(n_1035),
.Y(n_12259)
);

CKINVDCx16_ASAP7_75t_R g12260 ( 
.A(n_11325),
.Y(n_12260)
);

AOI21xp5_ASAP7_75t_L g12261 ( 
.A1(n_10932),
.A2(n_1036),
.B(n_1037),
.Y(n_12261)
);

AOI21xp5_ASAP7_75t_L g12262 ( 
.A1(n_10934),
.A2(n_1037),
.B(n_1038),
.Y(n_12262)
);

INVx2_ASAP7_75t_L g12263 ( 
.A(n_11430),
.Y(n_12263)
);

OAI21xp5_ASAP7_75t_L g12264 ( 
.A1(n_10956),
.A2(n_1038),
.B(n_1039),
.Y(n_12264)
);

NOR2xp33_ASAP7_75t_L g12265 ( 
.A(n_11249),
.B(n_1039),
.Y(n_12265)
);

BUFx6f_ASAP7_75t_L g12266 ( 
.A(n_10988),
.Y(n_12266)
);

INVx2_ASAP7_75t_L g12267 ( 
.A(n_11479),
.Y(n_12267)
);

NAND2xp5_ASAP7_75t_L g12268 ( 
.A(n_11279),
.B(n_1040),
.Y(n_12268)
);

NOR2xp33_ASAP7_75t_L g12269 ( 
.A(n_11091),
.B(n_1040),
.Y(n_12269)
);

NOR2xp33_ASAP7_75t_L g12270 ( 
.A(n_11070),
.B(n_1041),
.Y(n_12270)
);

NAND2xp5_ASAP7_75t_L g12271 ( 
.A(n_11233),
.B(n_1041),
.Y(n_12271)
);

OAI22xp5_ASAP7_75t_L g12272 ( 
.A1(n_11497),
.A2(n_1045),
.B1(n_1042),
.B2(n_1044),
.Y(n_12272)
);

O2A1O1Ixp5_ASAP7_75t_L g12273 ( 
.A1(n_10938),
.A2(n_1046),
.B(n_1042),
.C(n_1044),
.Y(n_12273)
);

AOI21xp5_ASAP7_75t_L g12274 ( 
.A1(n_10939),
.A2(n_1047),
.B(n_1048),
.Y(n_12274)
);

NAND2xp5_ASAP7_75t_SL g12275 ( 
.A(n_11078),
.B(n_1047),
.Y(n_12275)
);

NAND2xp5_ASAP7_75t_L g12276 ( 
.A(n_10957),
.B(n_10960),
.Y(n_12276)
);

INVx3_ASAP7_75t_SL g12277 ( 
.A(n_11302),
.Y(n_12277)
);

INVx1_ASAP7_75t_L g12278 ( 
.A(n_11427),
.Y(n_12278)
);

INVx2_ASAP7_75t_L g12279 ( 
.A(n_11498),
.Y(n_12279)
);

AO22x1_ASAP7_75t_L g12280 ( 
.A1(n_11500),
.A2(n_11601),
.B1(n_11587),
.B2(n_10975),
.Y(n_12280)
);

NOR3xp33_ASAP7_75t_L g12281 ( 
.A(n_11148),
.B(n_1049),
.C(n_1050),
.Y(n_12281)
);

INVx2_ASAP7_75t_L g12282 ( 
.A(n_11187),
.Y(n_12282)
);

AOI21xp5_ASAP7_75t_L g12283 ( 
.A1(n_10942),
.A2(n_1049),
.B(n_1050),
.Y(n_12283)
);

O2A1O1Ixp33_ASAP7_75t_L g12284 ( 
.A1(n_10970),
.A2(n_1053),
.B(n_1051),
.C(n_1052),
.Y(n_12284)
);

AO21x1_ASAP7_75t_L g12285 ( 
.A1(n_10978),
.A2(n_10990),
.B(n_10986),
.Y(n_12285)
);

INVx1_ASAP7_75t_L g12286 ( 
.A(n_11192),
.Y(n_12286)
);

OR2x6_ASAP7_75t_L g12287 ( 
.A(n_11257),
.B(n_1051),
.Y(n_12287)
);

BUFx6f_ASAP7_75t_L g12288 ( 
.A(n_11303),
.Y(n_12288)
);

INVx2_ASAP7_75t_L g12289 ( 
.A(n_11194),
.Y(n_12289)
);

BUFx2_ASAP7_75t_L g12290 ( 
.A(n_11260),
.Y(n_12290)
);

NAND2xp5_ASAP7_75t_L g12291 ( 
.A(n_10946),
.B(n_11195),
.Y(n_12291)
);

NAND2xp5_ASAP7_75t_L g12292 ( 
.A(n_11200),
.B(n_1052),
.Y(n_12292)
);

INVx1_ASAP7_75t_L g12293 ( 
.A(n_11204),
.Y(n_12293)
);

NAND2xp5_ASAP7_75t_L g12294 ( 
.A(n_11212),
.B(n_1053),
.Y(n_12294)
);

AOI21xp5_ASAP7_75t_L g12295 ( 
.A1(n_11272),
.A2(n_1054),
.B(n_1055),
.Y(n_12295)
);

NOR2xp33_ASAP7_75t_L g12296 ( 
.A(n_11275),
.B(n_1054),
.Y(n_12296)
);

NAND2xp5_ASAP7_75t_SL g12297 ( 
.A(n_11220),
.B(n_11225),
.Y(n_12297)
);

NAND2xp5_ASAP7_75t_L g12298 ( 
.A(n_10952),
.B(n_1056),
.Y(n_12298)
);

NAND2xp5_ASAP7_75t_SL g12299 ( 
.A(n_10950),
.B(n_1056),
.Y(n_12299)
);

OAI21xp33_ASAP7_75t_L g12300 ( 
.A1(n_10953),
.A2(n_1057),
.B(n_1058),
.Y(n_12300)
);

A2O1A1Ixp33_ASAP7_75t_L g12301 ( 
.A1(n_11007),
.A2(n_1060),
.B(n_1057),
.C(n_1059),
.Y(n_12301)
);

BUFx12f_ASAP7_75t_L g12302 ( 
.A(n_11012),
.Y(n_12302)
);

BUFx8_ASAP7_75t_L g12303 ( 
.A(n_11024),
.Y(n_12303)
);

OAI22xp5_ASAP7_75t_L g12304 ( 
.A1(n_10955),
.A2(n_1062),
.B1(n_1059),
.B2(n_1061),
.Y(n_12304)
);

O2A1O1Ixp33_ASAP7_75t_L g12305 ( 
.A1(n_11380),
.A2(n_1063),
.B(n_1061),
.C(n_1062),
.Y(n_12305)
);

AOI21xp5_ASAP7_75t_L g12306 ( 
.A1(n_10855),
.A2(n_1063),
.B(n_1064),
.Y(n_12306)
);

INVxp33_ASAP7_75t_SL g12307 ( 
.A(n_11451),
.Y(n_12307)
);

OAI22xp5_ASAP7_75t_L g12308 ( 
.A1(n_11383),
.A2(n_1067),
.B1(n_1065),
.B2(n_1066),
.Y(n_12308)
);

INVx1_ASAP7_75t_L g12309 ( 
.A(n_11111),
.Y(n_12309)
);

AOI21x1_ASAP7_75t_L g12310 ( 
.A1(n_10855),
.A2(n_1065),
.B(n_1066),
.Y(n_12310)
);

AOI21xp5_ASAP7_75t_L g12311 ( 
.A1(n_10855),
.A2(n_1067),
.B(n_1068),
.Y(n_12311)
);

INVx3_ASAP7_75t_L g12312 ( 
.A(n_11398),
.Y(n_12312)
);

NOR2xp33_ASAP7_75t_R g12313 ( 
.A(n_11451),
.B(n_1068),
.Y(n_12313)
);

HB1xp67_ASAP7_75t_L g12314 ( 
.A(n_11015),
.Y(n_12314)
);

O2A1O1Ixp33_ASAP7_75t_L g12315 ( 
.A1(n_11380),
.A2(n_1071),
.B(n_1069),
.C(n_1070),
.Y(n_12315)
);

AOI21xp5_ASAP7_75t_L g12316 ( 
.A1(n_10855),
.A2(n_1069),
.B(n_1070),
.Y(n_12316)
);

NAND2xp5_ASAP7_75t_SL g12317 ( 
.A(n_10855),
.B(n_1072),
.Y(n_12317)
);

AOI21xp5_ASAP7_75t_L g12318 ( 
.A1(n_10855),
.A2(n_1072),
.B(n_1073),
.Y(n_12318)
);

AOI21xp5_ASAP7_75t_L g12319 ( 
.A1(n_10855),
.A2(n_1074),
.B(n_1076),
.Y(n_12319)
);

O2A1O1Ixp5_ASAP7_75t_L g12320 ( 
.A1(n_11396),
.A2(n_1078),
.B(n_1074),
.C(n_1077),
.Y(n_12320)
);

AOI21xp5_ASAP7_75t_L g12321 ( 
.A1(n_10855),
.A2(n_1077),
.B(n_1079),
.Y(n_12321)
);

BUFx6f_ASAP7_75t_L g12322 ( 
.A(n_11398),
.Y(n_12322)
);

INVx4_ASAP7_75t_L g12323 ( 
.A(n_11559),
.Y(n_12323)
);

INVx1_ASAP7_75t_L g12324 ( 
.A(n_11111),
.Y(n_12324)
);

OAI21xp5_ASAP7_75t_L g12325 ( 
.A1(n_10855),
.A2(n_1080),
.B(n_1081),
.Y(n_12325)
);

NAND2xp5_ASAP7_75t_L g12326 ( 
.A(n_11015),
.B(n_1081),
.Y(n_12326)
);

BUFx6f_ASAP7_75t_L g12327 ( 
.A(n_11398),
.Y(n_12327)
);

AOI21x1_ASAP7_75t_L g12328 ( 
.A1(n_10855),
.A2(n_1082),
.B(n_1083),
.Y(n_12328)
);

NOR2xp33_ASAP7_75t_R g12329 ( 
.A(n_11451),
.B(n_1082),
.Y(n_12329)
);

NOR2xp33_ASAP7_75t_L g12330 ( 
.A(n_10856),
.B(n_1083),
.Y(n_12330)
);

NOR2x1p5_ASAP7_75t_L g12331 ( 
.A(n_11376),
.B(n_1084),
.Y(n_12331)
);

OAI21xp33_ASAP7_75t_L g12332 ( 
.A1(n_10826),
.A2(n_1084),
.B(n_1085),
.Y(n_12332)
);

O2A1O1Ixp33_ASAP7_75t_SL g12333 ( 
.A1(n_11251),
.A2(n_1087),
.B(n_1085),
.C(n_1086),
.Y(n_12333)
);

AND2x2_ASAP7_75t_L g12334 ( 
.A(n_10859),
.B(n_1088),
.Y(n_12334)
);

BUFx6f_ASAP7_75t_L g12335 ( 
.A(n_11398),
.Y(n_12335)
);

BUFx8_ASAP7_75t_L g12336 ( 
.A(n_10879),
.Y(n_12336)
);

NAND2xp5_ASAP7_75t_L g12337 ( 
.A(n_11015),
.B(n_1089),
.Y(n_12337)
);

NAND2xp5_ASAP7_75t_L g12338 ( 
.A(n_11015),
.B(n_1089),
.Y(n_12338)
);

OAI22xp5_ASAP7_75t_L g12339 ( 
.A1(n_11383),
.A2(n_1092),
.B1(n_1090),
.B2(n_1091),
.Y(n_12339)
);

NOR2xp33_ASAP7_75t_L g12340 ( 
.A(n_10856),
.B(n_1090),
.Y(n_12340)
);

NAND2xp5_ASAP7_75t_SL g12341 ( 
.A(n_10855),
.B(n_1091),
.Y(n_12341)
);

OAI21x1_ASAP7_75t_L g12342 ( 
.A1(n_10911),
.A2(n_1092),
.B(n_1093),
.Y(n_12342)
);

OAI22xp5_ASAP7_75t_L g12343 ( 
.A1(n_11383),
.A2(n_1095),
.B1(n_1093),
.B2(n_1094),
.Y(n_12343)
);

AOI21xp5_ASAP7_75t_L g12344 ( 
.A1(n_10855),
.A2(n_1094),
.B(n_1096),
.Y(n_12344)
);

NAND2xp5_ASAP7_75t_L g12345 ( 
.A(n_11015),
.B(n_1096),
.Y(n_12345)
);

NAND2xp5_ASAP7_75t_L g12346 ( 
.A(n_11015),
.B(n_1097),
.Y(n_12346)
);

BUFx3_ASAP7_75t_L g12347 ( 
.A(n_10991),
.Y(n_12347)
);

AOI21xp5_ASAP7_75t_L g12348 ( 
.A1(n_10855),
.A2(n_1097),
.B(n_1098),
.Y(n_12348)
);

NOR2xp33_ASAP7_75t_L g12349 ( 
.A(n_10856),
.B(n_1099),
.Y(n_12349)
);

AOI21xp5_ASAP7_75t_L g12350 ( 
.A1(n_10855),
.A2(n_1100),
.B(n_1101),
.Y(n_12350)
);

OAI22xp5_ASAP7_75t_L g12351 ( 
.A1(n_11383),
.A2(n_1102),
.B1(n_1100),
.B2(n_1101),
.Y(n_12351)
);

AND2x2_ASAP7_75t_L g12352 ( 
.A(n_10859),
.B(n_1102),
.Y(n_12352)
);

OA22x2_ASAP7_75t_L g12353 ( 
.A1(n_10928),
.A2(n_1105),
.B1(n_1103),
.B2(n_1104),
.Y(n_12353)
);

AOI21xp5_ASAP7_75t_L g12354 ( 
.A1(n_10855),
.A2(n_1103),
.B(n_1104),
.Y(n_12354)
);

AOI22xp5_ASAP7_75t_L g12355 ( 
.A1(n_10826),
.A2(n_1108),
.B1(n_1106),
.B2(n_1107),
.Y(n_12355)
);

AOI21xp5_ASAP7_75t_L g12356 ( 
.A1(n_10855),
.A2(n_1107),
.B(n_1109),
.Y(n_12356)
);

INVx2_ASAP7_75t_L g12357 ( 
.A(n_11266),
.Y(n_12357)
);

AOI21xp5_ASAP7_75t_L g12358 ( 
.A1(n_10855),
.A2(n_1110),
.B(n_1111),
.Y(n_12358)
);

CKINVDCx5p33_ASAP7_75t_R g12359 ( 
.A(n_11087),
.Y(n_12359)
);

AO21x1_ASAP7_75t_L g12360 ( 
.A1(n_11377),
.A2(n_1111),
.B(n_1112),
.Y(n_12360)
);

NAND2xp5_ASAP7_75t_SL g12361 ( 
.A(n_10855),
.B(n_1112),
.Y(n_12361)
);

BUFx6f_ASAP7_75t_L g12362 ( 
.A(n_11398),
.Y(n_12362)
);

AOI21xp5_ASAP7_75t_L g12363 ( 
.A1(n_10855),
.A2(n_1113),
.B(n_1114),
.Y(n_12363)
);

O2A1O1Ixp33_ASAP7_75t_L g12364 ( 
.A1(n_11380),
.A2(n_1115),
.B(n_1113),
.C(n_1114),
.Y(n_12364)
);

AOI21xp5_ASAP7_75t_L g12365 ( 
.A1(n_10855),
.A2(n_1115),
.B(n_1116),
.Y(n_12365)
);

INVx1_ASAP7_75t_L g12366 ( 
.A(n_11111),
.Y(n_12366)
);

O2A1O1Ixp33_ASAP7_75t_SL g12367 ( 
.A1(n_11251),
.A2(n_1118),
.B(n_1116),
.C(n_1117),
.Y(n_12367)
);

AOI22xp33_ASAP7_75t_L g12368 ( 
.A1(n_10826),
.A2(n_1120),
.B1(n_1117),
.B2(n_1119),
.Y(n_12368)
);

NAND2xp5_ASAP7_75t_SL g12369 ( 
.A(n_10855),
.B(n_1119),
.Y(n_12369)
);

HB1xp67_ASAP7_75t_L g12370 ( 
.A(n_11015),
.Y(n_12370)
);

AOI21xp5_ASAP7_75t_L g12371 ( 
.A1(n_10855),
.A2(n_1120),
.B(n_1121),
.Y(n_12371)
);

NAND2xp5_ASAP7_75t_SL g12372 ( 
.A(n_10855),
.B(n_1121),
.Y(n_12372)
);

AND2x4_ASAP7_75t_L g12373 ( 
.A(n_10907),
.B(n_1124),
.Y(n_12373)
);

INVxp67_ASAP7_75t_L g12374 ( 
.A(n_10949),
.Y(n_12374)
);

INVx3_ASAP7_75t_L g12375 ( 
.A(n_11398),
.Y(n_12375)
);

AND2x4_ASAP7_75t_L g12376 ( 
.A(n_10907),
.B(n_1124),
.Y(n_12376)
);

NAND2xp5_ASAP7_75t_L g12377 ( 
.A(n_11015),
.B(n_1125),
.Y(n_12377)
);

OA22x2_ASAP7_75t_L g12378 ( 
.A1(n_10928),
.A2(n_1127),
.B1(n_1125),
.B2(n_1126),
.Y(n_12378)
);

NAND2xp5_ASAP7_75t_SL g12379 ( 
.A(n_10855),
.B(n_1127),
.Y(n_12379)
);

INVx1_ASAP7_75t_SL g12380 ( 
.A(n_11067),
.Y(n_12380)
);

OA22x2_ASAP7_75t_L g12381 ( 
.A1(n_10928),
.A2(n_1130),
.B1(n_1128),
.B2(n_1129),
.Y(n_12381)
);

O2A1O1Ixp5_ASAP7_75t_L g12382 ( 
.A1(n_11396),
.A2(n_1130),
.B(n_1128),
.C(n_1129),
.Y(n_12382)
);

A2O1A1Ixp33_ASAP7_75t_L g12383 ( 
.A1(n_10826),
.A2(n_1133),
.B(n_1131),
.C(n_1132),
.Y(n_12383)
);

BUFx6f_ASAP7_75t_L g12384 ( 
.A(n_11398),
.Y(n_12384)
);

OAI22xp5_ASAP7_75t_L g12385 ( 
.A1(n_11383),
.A2(n_1136),
.B1(n_1134),
.B2(n_1135),
.Y(n_12385)
);

O2A1O1Ixp33_ASAP7_75t_L g12386 ( 
.A1(n_11380),
.A2(n_1139),
.B(n_1137),
.C(n_1138),
.Y(n_12386)
);

NOR2xp33_ASAP7_75t_L g12387 ( 
.A(n_10856),
.B(n_1137),
.Y(n_12387)
);

BUFx12f_ASAP7_75t_L g12388 ( 
.A(n_10879),
.Y(n_12388)
);

NAND2xp5_ASAP7_75t_L g12389 ( 
.A(n_11015),
.B(n_1138),
.Y(n_12389)
);

BUFx6f_ASAP7_75t_L g12390 ( 
.A(n_11398),
.Y(n_12390)
);

AOI21xp5_ASAP7_75t_L g12391 ( 
.A1(n_10855),
.A2(n_1139),
.B(n_1140),
.Y(n_12391)
);

NAND2xp5_ASAP7_75t_SL g12392 ( 
.A(n_10855),
.B(n_1141),
.Y(n_12392)
);

AOI21xp5_ASAP7_75t_L g12393 ( 
.A1(n_10855),
.A2(n_1141),
.B(n_1142),
.Y(n_12393)
);

AOI22xp5_ASAP7_75t_L g12394 ( 
.A1(n_10826),
.A2(n_1145),
.B1(n_1142),
.B2(n_1143),
.Y(n_12394)
);

INVx2_ASAP7_75t_L g12395 ( 
.A(n_11266),
.Y(n_12395)
);

INVx1_ASAP7_75t_L g12396 ( 
.A(n_11111),
.Y(n_12396)
);

INVx1_ASAP7_75t_L g12397 ( 
.A(n_11111),
.Y(n_12397)
);

NAND2xp5_ASAP7_75t_L g12398 ( 
.A(n_11015),
.B(n_1143),
.Y(n_12398)
);

AOI21xp5_ASAP7_75t_L g12399 ( 
.A1(n_10855),
.A2(n_1145),
.B(n_1146),
.Y(n_12399)
);

NAND2xp5_ASAP7_75t_L g12400 ( 
.A(n_11015),
.B(n_1147),
.Y(n_12400)
);

INVxp67_ASAP7_75t_L g12401 ( 
.A(n_10949),
.Y(n_12401)
);

CKINVDCx14_ASAP7_75t_R g12402 ( 
.A(n_11087),
.Y(n_12402)
);

OR2x6_ASAP7_75t_SL g12403 ( 
.A(n_11451),
.B(n_1147),
.Y(n_12403)
);

NAND2xp5_ASAP7_75t_L g12404 ( 
.A(n_11015),
.B(n_1148),
.Y(n_12404)
);

OAI21xp5_ASAP7_75t_L g12405 ( 
.A1(n_10855),
.A2(n_1148),
.B(n_1149),
.Y(n_12405)
);

O2A1O1Ixp33_ASAP7_75t_L g12406 ( 
.A1(n_11380),
.A2(n_1152),
.B(n_1150),
.C(n_1151),
.Y(n_12406)
);

AND2x4_ASAP7_75t_L g12407 ( 
.A(n_10907),
.B(n_1150),
.Y(n_12407)
);

OR2x2_ASAP7_75t_L g12408 ( 
.A(n_11015),
.B(n_1151),
.Y(n_12408)
);

NAND2xp5_ASAP7_75t_L g12409 ( 
.A(n_11015),
.B(n_1152),
.Y(n_12409)
);

NOR2x1_ASAP7_75t_SL g12410 ( 
.A(n_10911),
.B(n_1153),
.Y(n_12410)
);

AOI21xp5_ASAP7_75t_L g12411 ( 
.A1(n_10855),
.A2(n_1153),
.B(n_1154),
.Y(n_12411)
);

AOI21xp5_ASAP7_75t_L g12412 ( 
.A1(n_10855),
.A2(n_1155),
.B(n_1156),
.Y(n_12412)
);

OAI21xp5_ASAP7_75t_L g12413 ( 
.A1(n_10855),
.A2(n_1155),
.B(n_1156),
.Y(n_12413)
);

NAND2xp5_ASAP7_75t_L g12414 ( 
.A(n_11015),
.B(n_1157),
.Y(n_12414)
);

CKINVDCx8_ASAP7_75t_R g12415 ( 
.A(n_11471),
.Y(n_12415)
);

AOI21xp5_ASAP7_75t_L g12416 ( 
.A1(n_10855),
.A2(n_1157),
.B(n_1158),
.Y(n_12416)
);

INVx2_ASAP7_75t_L g12417 ( 
.A(n_11266),
.Y(n_12417)
);

INVx1_ASAP7_75t_L g12418 ( 
.A(n_11111),
.Y(n_12418)
);

NOR2xp33_ASAP7_75t_L g12419 ( 
.A(n_10856),
.B(n_1158),
.Y(n_12419)
);

OAI22xp5_ASAP7_75t_L g12420 ( 
.A1(n_11383),
.A2(n_1162),
.B1(n_1160),
.B2(n_1161),
.Y(n_12420)
);

NAND2xp5_ASAP7_75t_L g12421 ( 
.A(n_11015),
.B(n_1160),
.Y(n_12421)
);

INVx4_ASAP7_75t_L g12422 ( 
.A(n_11559),
.Y(n_12422)
);

NAND2xp5_ASAP7_75t_L g12423 ( 
.A(n_11015),
.B(n_1161),
.Y(n_12423)
);

NAND2xp5_ASAP7_75t_L g12424 ( 
.A(n_11015),
.B(n_1163),
.Y(n_12424)
);

AOI21xp5_ASAP7_75t_L g12425 ( 
.A1(n_10855),
.A2(n_1164),
.B(n_1165),
.Y(n_12425)
);

NOR2xp67_ASAP7_75t_L g12426 ( 
.A(n_11076),
.B(n_1164),
.Y(n_12426)
);

INVx2_ASAP7_75t_L g12427 ( 
.A(n_11266),
.Y(n_12427)
);

AOI22xp5_ASAP7_75t_L g12428 ( 
.A1(n_10826),
.A2(n_1169),
.B1(n_1166),
.B2(n_1168),
.Y(n_12428)
);

AOI21xp5_ASAP7_75t_L g12429 ( 
.A1(n_10855),
.A2(n_1166),
.B(n_1168),
.Y(n_12429)
);

AOI21xp5_ASAP7_75t_L g12430 ( 
.A1(n_10855),
.A2(n_1170),
.B(n_1171),
.Y(n_12430)
);

NAND2xp5_ASAP7_75t_L g12431 ( 
.A(n_11015),
.B(n_1170),
.Y(n_12431)
);

INVx1_ASAP7_75t_SL g12432 ( 
.A(n_11067),
.Y(n_12432)
);

INVx3_ASAP7_75t_SL g12433 ( 
.A(n_11451),
.Y(n_12433)
);

INVx3_ASAP7_75t_SL g12434 ( 
.A(n_11451),
.Y(n_12434)
);

OAI22xp5_ASAP7_75t_L g12435 ( 
.A1(n_11383),
.A2(n_1176),
.B1(n_1174),
.B2(n_1175),
.Y(n_12435)
);

NOR2xp33_ASAP7_75t_L g12436 ( 
.A(n_10856),
.B(n_1174),
.Y(n_12436)
);

O2A1O1Ixp33_ASAP7_75t_SL g12437 ( 
.A1(n_11251),
.A2(n_1177),
.B(n_1175),
.C(n_1176),
.Y(n_12437)
);

BUFx3_ASAP7_75t_L g12438 ( 
.A(n_10991),
.Y(n_12438)
);

OAI22xp5_ASAP7_75t_L g12439 ( 
.A1(n_11383),
.A2(n_1179),
.B1(n_1177),
.B2(n_1178),
.Y(n_12439)
);

NAND2xp5_ASAP7_75t_L g12440 ( 
.A(n_11015),
.B(n_1178),
.Y(n_12440)
);

NAND2xp5_ASAP7_75t_L g12441 ( 
.A(n_11015),
.B(n_1179),
.Y(n_12441)
);

OR2x2_ASAP7_75t_L g12442 ( 
.A(n_11015),
.B(n_1180),
.Y(n_12442)
);

HB1xp67_ASAP7_75t_L g12443 ( 
.A(n_11015),
.Y(n_12443)
);

A2O1A1Ixp33_ASAP7_75t_L g12444 ( 
.A1(n_10826),
.A2(n_1182),
.B(n_1180),
.C(n_1181),
.Y(n_12444)
);

INVx2_ASAP7_75t_L g12445 ( 
.A(n_11266),
.Y(n_12445)
);

AOI22xp5_ASAP7_75t_L g12446 ( 
.A1(n_10826),
.A2(n_1183),
.B1(n_1181),
.B2(n_1182),
.Y(n_12446)
);

NAND2xp5_ASAP7_75t_SL g12447 ( 
.A(n_10855),
.B(n_1183),
.Y(n_12447)
);

AOI21xp5_ASAP7_75t_L g12448 ( 
.A1(n_10855),
.A2(n_1184),
.B(n_1185),
.Y(n_12448)
);

O2A1O1Ixp33_ASAP7_75t_L g12449 ( 
.A1(n_11380),
.A2(n_1186),
.B(n_1184),
.C(n_1185),
.Y(n_12449)
);

AOI21xp5_ASAP7_75t_L g12450 ( 
.A1(n_10855),
.A2(n_1187),
.B(n_1188),
.Y(n_12450)
);

BUFx8_ASAP7_75t_L g12451 ( 
.A(n_10879),
.Y(n_12451)
);

AOI221xp5_ASAP7_75t_L g12452 ( 
.A1(n_10826),
.A2(n_1190),
.B1(n_1187),
.B2(n_1189),
.C(n_1191),
.Y(n_12452)
);

AND2x4_ASAP7_75t_L g12453 ( 
.A(n_10907),
.B(n_1189),
.Y(n_12453)
);

NOR2xp33_ASAP7_75t_L g12454 ( 
.A(n_10856),
.B(n_1191),
.Y(n_12454)
);

NOR2xp33_ASAP7_75t_SL g12455 ( 
.A(n_11051),
.B(n_1192),
.Y(n_12455)
);

AO32x1_ASAP7_75t_L g12456 ( 
.A1(n_11365),
.A2(n_1194),
.A3(n_1192),
.B1(n_1193),
.B2(n_1195),
.Y(n_12456)
);

O2A1O1Ixp33_ASAP7_75t_L g12457 ( 
.A1(n_11380),
.A2(n_1195),
.B(n_1193),
.C(n_1194),
.Y(n_12457)
);

OR2x6_ASAP7_75t_SL g12458 ( 
.A(n_11451),
.B(n_1196),
.Y(n_12458)
);

INVx1_ASAP7_75t_L g12459 ( 
.A(n_11111),
.Y(n_12459)
);

BUFx8_ASAP7_75t_SL g12460 ( 
.A(n_10879),
.Y(n_12460)
);

OAI22xp5_ASAP7_75t_L g12461 ( 
.A1(n_11383),
.A2(n_1199),
.B1(n_1197),
.B2(n_1198),
.Y(n_12461)
);

BUFx6f_ASAP7_75t_L g12462 ( 
.A(n_11398),
.Y(n_12462)
);

AOI21xp5_ASAP7_75t_L g12463 ( 
.A1(n_10855),
.A2(n_1197),
.B(n_1199),
.Y(n_12463)
);

INVx1_ASAP7_75t_L g12464 ( 
.A(n_11111),
.Y(n_12464)
);

INVx3_ASAP7_75t_L g12465 ( 
.A(n_11398),
.Y(n_12465)
);

INVx1_ASAP7_75t_L g12466 ( 
.A(n_11111),
.Y(n_12466)
);

NAND2xp5_ASAP7_75t_L g12467 ( 
.A(n_11015),
.B(n_1200),
.Y(n_12467)
);

OAI22xp5_ASAP7_75t_L g12468 ( 
.A1(n_11383),
.A2(n_1202),
.B1(n_1200),
.B2(n_1201),
.Y(n_12468)
);

O2A1O1Ixp5_ASAP7_75t_L g12469 ( 
.A1(n_11396),
.A2(n_1203),
.B(n_1201),
.C(n_1202),
.Y(n_12469)
);

NOR2xp33_ASAP7_75t_L g12470 ( 
.A(n_10856),
.B(n_1203),
.Y(n_12470)
);

NAND2xp5_ASAP7_75t_L g12471 ( 
.A(n_11015),
.B(n_1204),
.Y(n_12471)
);

OAI21xp5_ASAP7_75t_L g12472 ( 
.A1(n_10855),
.A2(n_1204),
.B(n_1205),
.Y(n_12472)
);

AOI22xp33_ASAP7_75t_L g12473 ( 
.A1(n_10826),
.A2(n_1208),
.B1(n_1206),
.B2(n_1207),
.Y(n_12473)
);

NAND2xp5_ASAP7_75t_L g12474 ( 
.A(n_11015),
.B(n_1206),
.Y(n_12474)
);

INVx2_ASAP7_75t_L g12475 ( 
.A(n_11266),
.Y(n_12475)
);

INVx1_ASAP7_75t_L g12476 ( 
.A(n_11111),
.Y(n_12476)
);

NAND2xp5_ASAP7_75t_SL g12477 ( 
.A(n_10855),
.B(n_1207),
.Y(n_12477)
);

AOI21xp5_ASAP7_75t_L g12478 ( 
.A1(n_10855),
.A2(n_1208),
.B(n_1209),
.Y(n_12478)
);

NAND2xp5_ASAP7_75t_L g12479 ( 
.A(n_11015),
.B(n_1209),
.Y(n_12479)
);

INVx2_ASAP7_75t_L g12480 ( 
.A(n_11266),
.Y(n_12480)
);

INVx2_ASAP7_75t_L g12481 ( 
.A(n_11266),
.Y(n_12481)
);

AOI21xp5_ASAP7_75t_L g12482 ( 
.A1(n_10855),
.A2(n_1210),
.B(n_1211),
.Y(n_12482)
);

NAND2xp5_ASAP7_75t_L g12483 ( 
.A(n_11015),
.B(n_1211),
.Y(n_12483)
);

NOR3xp33_ASAP7_75t_L g12484 ( 
.A(n_10826),
.B(n_1212),
.C(n_1213),
.Y(n_12484)
);

AOI21xp5_ASAP7_75t_L g12485 ( 
.A1(n_10855),
.A2(n_1212),
.B(n_1213),
.Y(n_12485)
);

AOI21xp5_ASAP7_75t_L g12486 ( 
.A1(n_10855),
.A2(n_1214),
.B(n_1215),
.Y(n_12486)
);

AOI21xp5_ASAP7_75t_L g12487 ( 
.A1(n_10855),
.A2(n_1215),
.B(n_1216),
.Y(n_12487)
);

AOI22xp5_ASAP7_75t_L g12488 ( 
.A1(n_10826),
.A2(n_1218),
.B1(n_1216),
.B2(n_1217),
.Y(n_12488)
);

AND2x2_ASAP7_75t_L g12489 ( 
.A(n_10859),
.B(n_1217),
.Y(n_12489)
);

NAND2xp5_ASAP7_75t_SL g12490 ( 
.A(n_10855),
.B(n_1218),
.Y(n_12490)
);

NOR2xp33_ASAP7_75t_SL g12491 ( 
.A(n_11051),
.B(n_1219),
.Y(n_12491)
);

AOI21xp5_ASAP7_75t_L g12492 ( 
.A1(n_10855),
.A2(n_1219),
.B(n_1220),
.Y(n_12492)
);

INVx2_ASAP7_75t_L g12493 ( 
.A(n_11266),
.Y(n_12493)
);

AOI21xp5_ASAP7_75t_L g12494 ( 
.A1(n_10855),
.A2(n_1220),
.B(n_1221),
.Y(n_12494)
);

OAI22xp5_ASAP7_75t_L g12495 ( 
.A1(n_11383),
.A2(n_1225),
.B1(n_1222),
.B2(n_1224),
.Y(n_12495)
);

NAND2xp5_ASAP7_75t_L g12496 ( 
.A(n_11015),
.B(n_1224),
.Y(n_12496)
);

NOR2xp33_ASAP7_75t_L g12497 ( 
.A(n_10856),
.B(n_1225),
.Y(n_12497)
);

NOR2xp33_ASAP7_75t_R g12498 ( 
.A(n_11451),
.B(n_1226),
.Y(n_12498)
);

NAND2xp5_ASAP7_75t_SL g12499 ( 
.A(n_10855),
.B(n_1226),
.Y(n_12499)
);

AND2x2_ASAP7_75t_L g12500 ( 
.A(n_10859),
.B(n_1227),
.Y(n_12500)
);

NOR2xp33_ASAP7_75t_L g12501 ( 
.A(n_10856),
.B(n_1227),
.Y(n_12501)
);

NOR2xp33_ASAP7_75t_L g12502 ( 
.A(n_10856),
.B(n_1228),
.Y(n_12502)
);

AOI21xp5_ASAP7_75t_L g12503 ( 
.A1(n_10855),
.A2(n_1228),
.B(n_1229),
.Y(n_12503)
);

NAND2xp5_ASAP7_75t_L g12504 ( 
.A(n_11015),
.B(n_1230),
.Y(n_12504)
);

NAND2xp5_ASAP7_75t_SL g12505 ( 
.A(n_10855),
.B(n_1230),
.Y(n_12505)
);

AOI22x1_ASAP7_75t_L g12506 ( 
.A1(n_11517),
.A2(n_1233),
.B1(n_1231),
.B2(n_1232),
.Y(n_12506)
);

AOI21xp5_ASAP7_75t_L g12507 ( 
.A1(n_10855),
.A2(n_1231),
.B(n_1232),
.Y(n_12507)
);

BUFx6f_ASAP7_75t_L g12508 ( 
.A(n_11398),
.Y(n_12508)
);

NOR2xp33_ASAP7_75t_L g12509 ( 
.A(n_10856),
.B(n_1234),
.Y(n_12509)
);

AOI21xp5_ASAP7_75t_L g12510 ( 
.A1(n_10855),
.A2(n_1234),
.B(n_1235),
.Y(n_12510)
);

INVx1_ASAP7_75t_L g12511 ( 
.A(n_11111),
.Y(n_12511)
);

AOI21xp5_ASAP7_75t_L g12512 ( 
.A1(n_10855),
.A2(n_1235),
.B(n_1236),
.Y(n_12512)
);

O2A1O1Ixp33_ASAP7_75t_L g12513 ( 
.A1(n_11380),
.A2(n_1238),
.B(n_1236),
.C(n_1237),
.Y(n_12513)
);

NAND2xp5_ASAP7_75t_L g12514 ( 
.A(n_11015),
.B(n_1237),
.Y(n_12514)
);

AOI21xp5_ASAP7_75t_L g12515 ( 
.A1(n_10855),
.A2(n_1238),
.B(n_1239),
.Y(n_12515)
);

NAND2xp5_ASAP7_75t_SL g12516 ( 
.A(n_10855),
.B(n_1239),
.Y(n_12516)
);

AND2x4_ASAP7_75t_L g12517 ( 
.A(n_10907),
.B(n_1240),
.Y(n_12517)
);

NAND2xp5_ASAP7_75t_L g12518 ( 
.A(n_11015),
.B(n_1241),
.Y(n_12518)
);

NOR2xp33_ASAP7_75t_L g12519 ( 
.A(n_10856),
.B(n_1241),
.Y(n_12519)
);

AOI22xp5_ASAP7_75t_L g12520 ( 
.A1(n_11832),
.A2(n_1244),
.B1(n_1242),
.B2(n_1243),
.Y(n_12520)
);

INVx3_ASAP7_75t_L g12521 ( 
.A(n_12102),
.Y(n_12521)
);

A2O1A1Ixp33_ASAP7_75t_L g12522 ( 
.A1(n_11722),
.A2(n_1244),
.B(n_1242),
.C(n_1243),
.Y(n_12522)
);

CKINVDCx20_ASAP7_75t_R g12523 ( 
.A(n_11748),
.Y(n_12523)
);

AOI22xp5_ASAP7_75t_L g12524 ( 
.A1(n_11656),
.A2(n_1247),
.B1(n_1245),
.B2(n_1246),
.Y(n_12524)
);

BUFx2_ASAP7_75t_L g12525 ( 
.A(n_11671),
.Y(n_12525)
);

NOR2xp33_ASAP7_75t_L g12526 ( 
.A(n_11924),
.B(n_1245),
.Y(n_12526)
);

INVx2_ASAP7_75t_L g12527 ( 
.A(n_11783),
.Y(n_12527)
);

NAND2xp5_ASAP7_75t_SL g12528 ( 
.A(n_12260),
.B(n_12232),
.Y(n_12528)
);

AND2x2_ASAP7_75t_L g12529 ( 
.A(n_11742),
.B(n_1246),
.Y(n_12529)
);

NAND2xp5_ASAP7_75t_L g12530 ( 
.A(n_12314),
.B(n_1247),
.Y(n_12530)
);

NOR2xp33_ASAP7_75t_L g12531 ( 
.A(n_11957),
.B(n_1248),
.Y(n_12531)
);

NAND2xp5_ASAP7_75t_L g12532 ( 
.A(n_12370),
.B(n_1248),
.Y(n_12532)
);

NAND2xp5_ASAP7_75t_L g12533 ( 
.A(n_12443),
.B(n_1249),
.Y(n_12533)
);

NAND2xp5_ASAP7_75t_L g12534 ( 
.A(n_11661),
.B(n_1249),
.Y(n_12534)
);

NAND2xp5_ASAP7_75t_L g12535 ( 
.A(n_12374),
.B(n_1250),
.Y(n_12535)
);

OR2x2_ASAP7_75t_L g12536 ( 
.A(n_11607),
.B(n_1250),
.Y(n_12536)
);

BUFx3_ASAP7_75t_L g12537 ( 
.A(n_11896),
.Y(n_12537)
);

NAND2xp5_ASAP7_75t_L g12538 ( 
.A(n_12401),
.B(n_1251),
.Y(n_12538)
);

HB1xp67_ASAP7_75t_L g12539 ( 
.A(n_11824),
.Y(n_12539)
);

INVx2_ASAP7_75t_L g12540 ( 
.A(n_11800),
.Y(n_12540)
);

AND2x2_ASAP7_75t_L g12541 ( 
.A(n_11743),
.B(n_11687),
.Y(n_12541)
);

CKINVDCx5p33_ASAP7_75t_R g12542 ( 
.A(n_11917),
.Y(n_12542)
);

BUFx6f_ASAP7_75t_L g12543 ( 
.A(n_11614),
.Y(n_12543)
);

CKINVDCx5p33_ASAP7_75t_R g12544 ( 
.A(n_12460),
.Y(n_12544)
);

AND3x1_ASAP7_75t_SL g12545 ( 
.A(n_12331),
.B(n_1251),
.C(n_1252),
.Y(n_12545)
);

NAND2xp5_ASAP7_75t_SL g12546 ( 
.A(n_12218),
.B(n_1252),
.Y(n_12546)
);

OAI21xp5_ASAP7_75t_L g12547 ( 
.A1(n_11680),
.A2(n_1253),
.B(n_1254),
.Y(n_12547)
);

INVx1_ASAP7_75t_L g12548 ( 
.A(n_11937),
.Y(n_12548)
);

OAI22xp5_ASAP7_75t_L g12549 ( 
.A1(n_11718),
.A2(n_1255),
.B1(n_1253),
.B2(n_1254),
.Y(n_12549)
);

INVx3_ASAP7_75t_L g12550 ( 
.A(n_12102),
.Y(n_12550)
);

NAND2xp5_ASAP7_75t_L g12551 ( 
.A(n_12004),
.B(n_1255),
.Y(n_12551)
);

BUFx6f_ASAP7_75t_L g12552 ( 
.A(n_11614),
.Y(n_12552)
);

CKINVDCx5p33_ASAP7_75t_R g12553 ( 
.A(n_12359),
.Y(n_12553)
);

NAND2xp5_ASAP7_75t_L g12554 ( 
.A(n_12003),
.B(n_1256),
.Y(n_12554)
);

INVx2_ASAP7_75t_SL g12555 ( 
.A(n_11961),
.Y(n_12555)
);

NAND2xp5_ASAP7_75t_L g12556 ( 
.A(n_11703),
.B(n_1256),
.Y(n_12556)
);

INVx2_ASAP7_75t_L g12557 ( 
.A(n_11813),
.Y(n_12557)
);

HB1xp67_ASAP7_75t_L g12558 ( 
.A(n_11625),
.Y(n_12558)
);

AOI22xp5_ASAP7_75t_L g12559 ( 
.A1(n_11751),
.A2(n_11953),
.B1(n_11690),
.B2(n_12484),
.Y(n_12559)
);

NAND2xp5_ASAP7_75t_L g12560 ( 
.A(n_12222),
.B(n_1257),
.Y(n_12560)
);

INVx2_ASAP7_75t_L g12561 ( 
.A(n_11823),
.Y(n_12561)
);

INVxp33_ASAP7_75t_SL g12562 ( 
.A(n_11776),
.Y(n_12562)
);

INVx1_ASAP7_75t_L g12563 ( 
.A(n_11642),
.Y(n_12563)
);

BUFx3_ASAP7_75t_L g12564 ( 
.A(n_11771),
.Y(n_12564)
);

AND3x1_ASAP7_75t_SL g12565 ( 
.A(n_12452),
.B(n_1257),
.C(n_1258),
.Y(n_12565)
);

NAND3xp33_ASAP7_75t_SL g12566 ( 
.A(n_12325),
.B(n_1258),
.C(n_1259),
.Y(n_12566)
);

INVxp67_ASAP7_75t_SL g12567 ( 
.A(n_11762),
.Y(n_12567)
);

INVx1_ASAP7_75t_L g12568 ( 
.A(n_11644),
.Y(n_12568)
);

AND2x2_ASAP7_75t_L g12569 ( 
.A(n_11627),
.B(n_1259),
.Y(n_12569)
);

CKINVDCx5p33_ASAP7_75t_R g12570 ( 
.A(n_12402),
.Y(n_12570)
);

INVxp67_ASAP7_75t_L g12571 ( 
.A(n_12027),
.Y(n_12571)
);

AND3x1_ASAP7_75t_SL g12572 ( 
.A(n_12251),
.B(n_1260),
.C(n_1261),
.Y(n_12572)
);

OAI22xp5_ASAP7_75t_SL g12573 ( 
.A1(n_11757),
.A2(n_1262),
.B1(n_1260),
.B2(n_1261),
.Y(n_12573)
);

CKINVDCx5p33_ASAP7_75t_R g12574 ( 
.A(n_12023),
.Y(n_12574)
);

AND2x6_ASAP7_75t_L g12575 ( 
.A(n_11943),
.B(n_1262),
.Y(n_12575)
);

CKINVDCx5p33_ASAP7_75t_R g12576 ( 
.A(n_11704),
.Y(n_12576)
);

INVx1_ASAP7_75t_L g12577 ( 
.A(n_11652),
.Y(n_12577)
);

AND2x2_ASAP7_75t_L g12578 ( 
.A(n_12309),
.B(n_1263),
.Y(n_12578)
);

OAI22xp5_ASAP7_75t_L g12579 ( 
.A1(n_11615),
.A2(n_1265),
.B1(n_1263),
.B2(n_1264),
.Y(n_12579)
);

HB1xp67_ASAP7_75t_L g12580 ( 
.A(n_12324),
.Y(n_12580)
);

INVx2_ASAP7_75t_L g12581 ( 
.A(n_11842),
.Y(n_12581)
);

INVxp67_ASAP7_75t_L g12582 ( 
.A(n_12235),
.Y(n_12582)
);

INVx1_ASAP7_75t_L g12583 ( 
.A(n_11653),
.Y(n_12583)
);

NAND2xp5_ASAP7_75t_L g12584 ( 
.A(n_12366),
.B(n_1264),
.Y(n_12584)
);

BUFx6f_ASAP7_75t_L g12585 ( 
.A(n_12322),
.Y(n_12585)
);

INVxp67_ASAP7_75t_L g12586 ( 
.A(n_11730),
.Y(n_12586)
);

AND2x2_ASAP7_75t_L g12587 ( 
.A(n_12511),
.B(n_1265),
.Y(n_12587)
);

NAND2xp5_ASAP7_75t_L g12588 ( 
.A(n_12396),
.B(n_1266),
.Y(n_12588)
);

AND2x2_ASAP7_75t_L g12589 ( 
.A(n_12397),
.B(n_1266),
.Y(n_12589)
);

INVx2_ASAP7_75t_L g12590 ( 
.A(n_11897),
.Y(n_12590)
);

CKINVDCx11_ASAP7_75t_R g12591 ( 
.A(n_12415),
.Y(n_12591)
);

INVx1_ASAP7_75t_L g12592 ( 
.A(n_11660),
.Y(n_12592)
);

NOR2xp33_ASAP7_75t_L g12593 ( 
.A(n_12139),
.B(n_1267),
.Y(n_12593)
);

INVx2_ASAP7_75t_L g12594 ( 
.A(n_11945),
.Y(n_12594)
);

INVx2_ASAP7_75t_L g12595 ( 
.A(n_12002),
.Y(n_12595)
);

AND3x1_ASAP7_75t_SL g12596 ( 
.A(n_12258),
.B(n_12278),
.C(n_11855),
.Y(n_12596)
);

INVx1_ASAP7_75t_L g12597 ( 
.A(n_11662),
.Y(n_12597)
);

NAND2xp5_ASAP7_75t_L g12598 ( 
.A(n_12418),
.B(n_1267),
.Y(n_12598)
);

NAND2xp5_ASAP7_75t_L g12599 ( 
.A(n_12459),
.B(n_1268),
.Y(n_12599)
);

INVx2_ASAP7_75t_L g12600 ( 
.A(n_11995),
.Y(n_12600)
);

NAND2xp5_ASAP7_75t_L g12601 ( 
.A(n_12464),
.B(n_1268),
.Y(n_12601)
);

NAND2xp5_ASAP7_75t_SL g12602 ( 
.A(n_12124),
.B(n_12290),
.Y(n_12602)
);

CKINVDCx5p33_ASAP7_75t_R g12603 ( 
.A(n_12307),
.Y(n_12603)
);

INVx2_ASAP7_75t_L g12604 ( 
.A(n_11630),
.Y(n_12604)
);

INVx1_ASAP7_75t_L g12605 ( 
.A(n_11711),
.Y(n_12605)
);

INVxp67_ASAP7_75t_L g12606 ( 
.A(n_12252),
.Y(n_12606)
);

NAND2xp5_ASAP7_75t_L g12607 ( 
.A(n_12466),
.B(n_1269),
.Y(n_12607)
);

INVx1_ASAP7_75t_L g12608 ( 
.A(n_11719),
.Y(n_12608)
);

OAI21xp5_ASAP7_75t_L g12609 ( 
.A1(n_12306),
.A2(n_1269),
.B(n_1270),
.Y(n_12609)
);

NAND2xp5_ASAP7_75t_SL g12610 ( 
.A(n_12256),
.B(n_11876),
.Y(n_12610)
);

AND2x2_ASAP7_75t_L g12611 ( 
.A(n_12476),
.B(n_1270),
.Y(n_12611)
);

AND2x2_ASAP7_75t_L g12612 ( 
.A(n_12380),
.B(n_1271),
.Y(n_12612)
);

INVx1_ASAP7_75t_L g12613 ( 
.A(n_11736),
.Y(n_12613)
);

NAND2xp5_ASAP7_75t_L g12614 ( 
.A(n_12096),
.B(n_11633),
.Y(n_12614)
);

CKINVDCx16_ASAP7_75t_R g12615 ( 
.A(n_12313),
.Y(n_12615)
);

INVx1_ASAP7_75t_SL g12616 ( 
.A(n_11916),
.Y(n_12616)
);

OAI22xp5_ASAP7_75t_L g12617 ( 
.A1(n_11609),
.A2(n_11616),
.B1(n_11681),
.B2(n_11629),
.Y(n_12617)
);

NAND2xp5_ASAP7_75t_L g12618 ( 
.A(n_11699),
.B(n_1271),
.Y(n_12618)
);

INVx3_ASAP7_75t_L g12619 ( 
.A(n_12081),
.Y(n_12619)
);

NAND2xp5_ASAP7_75t_L g12620 ( 
.A(n_11750),
.B(n_12357),
.Y(n_12620)
);

NAND2xp5_ASAP7_75t_L g12621 ( 
.A(n_12395),
.B(n_1272),
.Y(n_12621)
);

NAND2xp5_ASAP7_75t_SL g12622 ( 
.A(n_12266),
.B(n_1272),
.Y(n_12622)
);

INVx2_ASAP7_75t_L g12623 ( 
.A(n_12417),
.Y(n_12623)
);

INVx2_ASAP7_75t_L g12624 ( 
.A(n_12427),
.Y(n_12624)
);

INVx2_ASAP7_75t_L g12625 ( 
.A(n_12445),
.Y(n_12625)
);

NAND2xp5_ASAP7_75t_L g12626 ( 
.A(n_12475),
.B(n_1273),
.Y(n_12626)
);

INVx2_ASAP7_75t_L g12627 ( 
.A(n_12480),
.Y(n_12627)
);

INVx2_ASAP7_75t_L g12628 ( 
.A(n_12481),
.Y(n_12628)
);

INVx1_ASAP7_75t_L g12629 ( 
.A(n_11747),
.Y(n_12629)
);

INVx1_ASAP7_75t_L g12630 ( 
.A(n_11756),
.Y(n_12630)
);

INVx2_ASAP7_75t_L g12631 ( 
.A(n_12493),
.Y(n_12631)
);

BUFx2_ASAP7_75t_L g12632 ( 
.A(n_12036),
.Y(n_12632)
);

CKINVDCx20_ASAP7_75t_R g12633 ( 
.A(n_11688),
.Y(n_12633)
);

CKINVDCx8_ASAP7_75t_R g12634 ( 
.A(n_11761),
.Y(n_12634)
);

AOI22xp33_ASAP7_75t_SL g12635 ( 
.A1(n_12506),
.A2(n_1275),
.B1(n_1273),
.B2(n_1274),
.Y(n_12635)
);

INVx1_ASAP7_75t_L g12636 ( 
.A(n_11767),
.Y(n_12636)
);

AND2x2_ASAP7_75t_L g12637 ( 
.A(n_12432),
.B(n_1275),
.Y(n_12637)
);

NAND2xp33_ASAP7_75t_R g12638 ( 
.A(n_12329),
.B(n_1277),
.Y(n_12638)
);

NAND2xp5_ASAP7_75t_L g12639 ( 
.A(n_11689),
.B(n_1277),
.Y(n_12639)
);

AND2x2_ASAP7_75t_L g12640 ( 
.A(n_12107),
.B(n_1278),
.Y(n_12640)
);

INVx1_ASAP7_75t_L g12641 ( 
.A(n_11806),
.Y(n_12641)
);

AND2x2_ASAP7_75t_L g12642 ( 
.A(n_12161),
.B(n_1278),
.Y(n_12642)
);

NAND2xp5_ASAP7_75t_L g12643 ( 
.A(n_12207),
.B(n_1279),
.Y(n_12643)
);

OAI22xp5_ASAP7_75t_L g12644 ( 
.A1(n_11621),
.A2(n_1281),
.B1(n_1279),
.B2(n_1280),
.Y(n_12644)
);

NOR2xp33_ASAP7_75t_L g12645 ( 
.A(n_12033),
.B(n_1280),
.Y(n_12645)
);

INVx1_ASAP7_75t_L g12646 ( 
.A(n_11828),
.Y(n_12646)
);

INVx2_ASAP7_75t_L g12647 ( 
.A(n_11838),
.Y(n_12647)
);

AND2x4_ASAP7_75t_L g12648 ( 
.A(n_11738),
.B(n_1281),
.Y(n_12648)
);

INVx2_ASAP7_75t_L g12649 ( 
.A(n_11849),
.Y(n_12649)
);

AND2x2_ASAP7_75t_L g12650 ( 
.A(n_11880),
.B(n_1282),
.Y(n_12650)
);

INVx2_ASAP7_75t_SL g12651 ( 
.A(n_12075),
.Y(n_12651)
);

BUFx2_ASAP7_75t_L g12652 ( 
.A(n_12347),
.Y(n_12652)
);

INVx2_ASAP7_75t_L g12653 ( 
.A(n_11854),
.Y(n_12653)
);

INVx1_ASAP7_75t_L g12654 ( 
.A(n_11879),
.Y(n_12654)
);

NAND2xp5_ASAP7_75t_L g12655 ( 
.A(n_12224),
.B(n_12058),
.Y(n_12655)
);

AND2x2_ASAP7_75t_L g12656 ( 
.A(n_12208),
.B(n_1282),
.Y(n_12656)
);

CKINVDCx5p33_ASAP7_75t_R g12657 ( 
.A(n_11705),
.Y(n_12657)
);

NOR2xp33_ASAP7_75t_L g12658 ( 
.A(n_12153),
.B(n_1283),
.Y(n_12658)
);

INVx1_ASAP7_75t_L g12659 ( 
.A(n_11882),
.Y(n_12659)
);

AND2x2_ASAP7_75t_L g12660 ( 
.A(n_11920),
.B(n_11930),
.Y(n_12660)
);

HB1xp67_ASAP7_75t_L g12661 ( 
.A(n_11936),
.Y(n_12661)
);

INVx2_ASAP7_75t_L g12662 ( 
.A(n_11940),
.Y(n_12662)
);

BUFx2_ASAP7_75t_L g12663 ( 
.A(n_12438),
.Y(n_12663)
);

NAND2xp5_ASAP7_75t_L g12664 ( 
.A(n_12063),
.B(n_1284),
.Y(n_12664)
);

AOI22xp5_ASAP7_75t_L g12665 ( 
.A1(n_11624),
.A2(n_1287),
.B1(n_1285),
.B2(n_1286),
.Y(n_12665)
);

NAND2xp5_ASAP7_75t_L g12666 ( 
.A(n_12064),
.B(n_1285),
.Y(n_12666)
);

INVx2_ASAP7_75t_L g12667 ( 
.A(n_11948),
.Y(n_12667)
);

INVx1_ASAP7_75t_L g12668 ( 
.A(n_11951),
.Y(n_12668)
);

INVx1_ASAP7_75t_L g12669 ( 
.A(n_11986),
.Y(n_12669)
);

AND2x2_ASAP7_75t_L g12670 ( 
.A(n_12250),
.B(n_1286),
.Y(n_12670)
);

CKINVDCx5p33_ASAP7_75t_R g12671 ( 
.A(n_11745),
.Y(n_12671)
);

AO22x1_ASAP7_75t_L g12672 ( 
.A1(n_11654),
.A2(n_1289),
.B1(n_1287),
.B2(n_1288),
.Y(n_12672)
);

NAND2xp5_ASAP7_75t_L g12673 ( 
.A(n_12080),
.B(n_1288),
.Y(n_12673)
);

NAND2xp5_ASAP7_75t_L g12674 ( 
.A(n_12082),
.B(n_1289),
.Y(n_12674)
);

AND2x2_ASAP7_75t_L g12675 ( 
.A(n_11859),
.B(n_1290),
.Y(n_12675)
);

CKINVDCx20_ASAP7_75t_R g12676 ( 
.A(n_12336),
.Y(n_12676)
);

NAND2xp5_ASAP7_75t_L g12677 ( 
.A(n_12095),
.B(n_1291),
.Y(n_12677)
);

AOI22xp5_ASAP7_75t_L g12678 ( 
.A1(n_12062),
.A2(n_1293),
.B1(n_1291),
.B2(n_1292),
.Y(n_12678)
);

OAI22xp5_ASAP7_75t_L g12679 ( 
.A1(n_11793),
.A2(n_1294),
.B1(n_1292),
.B2(n_1293),
.Y(n_12679)
);

BUFx8_ASAP7_75t_SL g12680 ( 
.A(n_12388),
.Y(n_12680)
);

NAND2xp5_ASAP7_75t_L g12681 ( 
.A(n_12098),
.B(n_12112),
.Y(n_12681)
);

INVx3_ASAP7_75t_L g12682 ( 
.A(n_12055),
.Y(n_12682)
);

AND2x2_ASAP7_75t_L g12683 ( 
.A(n_12053),
.B(n_12056),
.Y(n_12683)
);

INVx2_ASAP7_75t_L g12684 ( 
.A(n_12014),
.Y(n_12684)
);

OAI21xp5_ASAP7_75t_L g12685 ( 
.A1(n_12311),
.A2(n_1294),
.B(n_1295),
.Y(n_12685)
);

AND3x1_ASAP7_75t_SL g12686 ( 
.A(n_12061),
.B(n_1295),
.C(n_1296),
.Y(n_12686)
);

NAND2x1_ASAP7_75t_L g12687 ( 
.A(n_12263),
.B(n_1296),
.Y(n_12687)
);

NAND2xp5_ASAP7_75t_L g12688 ( 
.A(n_12132),
.B(n_1297),
.Y(n_12688)
);

NAND2xp5_ASAP7_75t_L g12689 ( 
.A(n_12157),
.B(n_1297),
.Y(n_12689)
);

AND2x2_ASAP7_75t_L g12690 ( 
.A(n_12088),
.B(n_1298),
.Y(n_12690)
);

INVx1_ASAP7_75t_L g12691 ( 
.A(n_11990),
.Y(n_12691)
);

NAND2xp5_ASAP7_75t_L g12692 ( 
.A(n_12177),
.B(n_1298),
.Y(n_12692)
);

AND2x2_ASAP7_75t_SL g12693 ( 
.A(n_12070),
.B(n_12247),
.Y(n_12693)
);

INVx2_ASAP7_75t_L g12694 ( 
.A(n_12188),
.Y(n_12694)
);

INVx2_ASAP7_75t_L g12695 ( 
.A(n_12122),
.Y(n_12695)
);

INVx2_ASAP7_75t_L g12696 ( 
.A(n_12144),
.Y(n_12696)
);

INVx1_ASAP7_75t_L g12697 ( 
.A(n_12408),
.Y(n_12697)
);

BUFx8_ASAP7_75t_L g12698 ( 
.A(n_11833),
.Y(n_12698)
);

OAI21xp5_ASAP7_75t_L g12699 ( 
.A1(n_12316),
.A2(n_1299),
.B(n_1300),
.Y(n_12699)
);

INVx1_ASAP7_75t_L g12700 ( 
.A(n_12442),
.Y(n_12700)
);

BUFx2_ASAP7_75t_L g12701 ( 
.A(n_11693),
.Y(n_12701)
);

INVx2_ASAP7_75t_L g12702 ( 
.A(n_12154),
.Y(n_12702)
);

INVx1_ASAP7_75t_L g12703 ( 
.A(n_12165),
.Y(n_12703)
);

AND2x2_ASAP7_75t_L g12704 ( 
.A(n_12106),
.B(n_1299),
.Y(n_12704)
);

INVx1_ASAP7_75t_L g12705 ( 
.A(n_12117),
.Y(n_12705)
);

NAND2xp5_ASAP7_75t_L g12706 ( 
.A(n_12105),
.B(n_1300),
.Y(n_12706)
);

INVx1_ASAP7_75t_L g12707 ( 
.A(n_11606),
.Y(n_12707)
);

NOR2xp33_ASAP7_75t_L g12708 ( 
.A(n_12230),
.B(n_1301),
.Y(n_12708)
);

NAND2xp5_ASAP7_75t_L g12709 ( 
.A(n_11846),
.B(n_1301),
.Y(n_12709)
);

INVx6_ASAP7_75t_L g12710 ( 
.A(n_11780),
.Y(n_12710)
);

OAI21xp5_ASAP7_75t_L g12711 ( 
.A1(n_12318),
.A2(n_1302),
.B(n_1303),
.Y(n_12711)
);

NAND2xp5_ASAP7_75t_L g12712 ( 
.A(n_12514),
.B(n_1302),
.Y(n_12712)
);

OAI21x1_ASAP7_75t_L g12713 ( 
.A1(n_11655),
.A2(n_12203),
.B(n_12198),
.Y(n_12713)
);

INVx2_ASAP7_75t_L g12714 ( 
.A(n_11613),
.Y(n_12714)
);

INVx1_ASAP7_75t_L g12715 ( 
.A(n_12338),
.Y(n_12715)
);

BUFx6f_ASAP7_75t_L g12716 ( 
.A(n_12322),
.Y(n_12716)
);

INVx2_ASAP7_75t_L g12717 ( 
.A(n_12326),
.Y(n_12717)
);

NAND2xp5_ASAP7_75t_L g12718 ( 
.A(n_12504),
.B(n_1303),
.Y(n_12718)
);

OAI22xp5_ASAP7_75t_L g12719 ( 
.A1(n_11938),
.A2(n_1306),
.B1(n_1304),
.B2(n_1305),
.Y(n_12719)
);

NOR2xp33_ASAP7_75t_R g12720 ( 
.A(n_11946),
.B(n_1305),
.Y(n_12720)
);

AND3x1_ASAP7_75t_SL g12721 ( 
.A(n_11619),
.B(n_1307),
.C(n_1308),
.Y(n_12721)
);

INVx6_ASAP7_75t_L g12722 ( 
.A(n_12451),
.Y(n_12722)
);

INVx1_ASAP7_75t_L g12723 ( 
.A(n_12337),
.Y(n_12723)
);

BUFx3_ASAP7_75t_L g12724 ( 
.A(n_12075),
.Y(n_12724)
);

INVx2_ASAP7_75t_L g12725 ( 
.A(n_12345),
.Y(n_12725)
);

NAND2xp5_ASAP7_75t_L g12726 ( 
.A(n_12518),
.B(n_1307),
.Y(n_12726)
);

AND2x2_ASAP7_75t_SL g12727 ( 
.A(n_12159),
.B(n_1308),
.Y(n_12727)
);

NOR2xp33_ASAP7_75t_R g12728 ( 
.A(n_12149),
.B(n_1309),
.Y(n_12728)
);

CKINVDCx8_ASAP7_75t_R g12729 ( 
.A(n_11784),
.Y(n_12729)
);

BUFx6f_ASAP7_75t_L g12730 ( 
.A(n_12327),
.Y(n_12730)
);

OAI22xp5_ASAP7_75t_SL g12731 ( 
.A1(n_12120),
.A2(n_1312),
.B1(n_1310),
.B2(n_1311),
.Y(n_12731)
);

AND2x2_ASAP7_75t_L g12732 ( 
.A(n_12137),
.B(n_1310),
.Y(n_12732)
);

AND2x2_ASAP7_75t_L g12733 ( 
.A(n_12133),
.B(n_1311),
.Y(n_12733)
);

AND3x1_ASAP7_75t_SL g12734 ( 
.A(n_12403),
.B(n_1313),
.C(n_1314),
.Y(n_12734)
);

CKINVDCx5p33_ASAP7_75t_R g12735 ( 
.A(n_11778),
.Y(n_12735)
);

AND2x4_ASAP7_75t_L g12736 ( 
.A(n_11708),
.B(n_1313),
.Y(n_12736)
);

CKINVDCx8_ASAP7_75t_R g12737 ( 
.A(n_12104),
.Y(n_12737)
);

NAND2xp5_ASAP7_75t_L g12738 ( 
.A(n_12346),
.B(n_1315),
.Y(n_12738)
);

OAI22xp5_ASAP7_75t_SL g12739 ( 
.A1(n_11881),
.A2(n_1317),
.B1(n_1315),
.B2(n_1316),
.Y(n_12739)
);

BUFx2_ASAP7_75t_L g12740 ( 
.A(n_11693),
.Y(n_12740)
);

NOR2x1_ASAP7_75t_L g12741 ( 
.A(n_12377),
.B(n_1316),
.Y(n_12741)
);

NAND2xp5_ASAP7_75t_SL g12742 ( 
.A(n_12266),
.B(n_1317),
.Y(n_12742)
);

INVx2_ASAP7_75t_SL g12743 ( 
.A(n_11875),
.Y(n_12743)
);

INVx2_ASAP7_75t_L g12744 ( 
.A(n_12389),
.Y(n_12744)
);

INVxp67_ASAP7_75t_L g12745 ( 
.A(n_11707),
.Y(n_12745)
);

CKINVDCx11_ASAP7_75t_R g12746 ( 
.A(n_12458),
.Y(n_12746)
);

HB1xp67_ASAP7_75t_L g12747 ( 
.A(n_12398),
.Y(n_12747)
);

HB1xp67_ASAP7_75t_L g12748 ( 
.A(n_12400),
.Y(n_12748)
);

AND2x2_ASAP7_75t_L g12749 ( 
.A(n_12172),
.B(n_1318),
.Y(n_12749)
);

NAND2xp5_ASAP7_75t_L g12750 ( 
.A(n_12404),
.B(n_1318),
.Y(n_12750)
);

BUFx3_ASAP7_75t_L g12751 ( 
.A(n_12186),
.Y(n_12751)
);

INVx4_ASAP7_75t_L g12752 ( 
.A(n_12433),
.Y(n_12752)
);

NOR2x1_ASAP7_75t_L g12753 ( 
.A(n_12409),
.B(n_1319),
.Y(n_12753)
);

NAND3xp33_ASAP7_75t_SL g12754 ( 
.A(n_12405),
.B(n_1319),
.C(n_1321),
.Y(n_12754)
);

BUFx4f_ASAP7_75t_L g12755 ( 
.A(n_12434),
.Y(n_12755)
);

BUFx3_ASAP7_75t_L g12756 ( 
.A(n_11691),
.Y(n_12756)
);

CKINVDCx5p33_ASAP7_75t_R g12757 ( 
.A(n_12019),
.Y(n_12757)
);

INVx1_ASAP7_75t_L g12758 ( 
.A(n_12414),
.Y(n_12758)
);

AND2x4_ASAP7_75t_L g12759 ( 
.A(n_11721),
.B(n_1321),
.Y(n_12759)
);

NAND2xp5_ASAP7_75t_L g12760 ( 
.A(n_12421),
.B(n_1322),
.Y(n_12760)
);

NAND2xp5_ASAP7_75t_L g12761 ( 
.A(n_12423),
.B(n_1322),
.Y(n_12761)
);

INVx2_ASAP7_75t_L g12762 ( 
.A(n_12424),
.Y(n_12762)
);

AND2x2_ASAP7_75t_L g12763 ( 
.A(n_11657),
.B(n_1323),
.Y(n_12763)
);

AND2x2_ASAP7_75t_L g12764 ( 
.A(n_11732),
.B(n_1323),
.Y(n_12764)
);

AND2x2_ASAP7_75t_L g12765 ( 
.A(n_11753),
.B(n_1324),
.Y(n_12765)
);

INVxp67_ASAP7_75t_L g12766 ( 
.A(n_11720),
.Y(n_12766)
);

BUFx3_ASAP7_75t_L g12767 ( 
.A(n_11887),
.Y(n_12767)
);

NOR3xp33_ASAP7_75t_L g12768 ( 
.A(n_11676),
.B(n_1324),
.C(n_1325),
.Y(n_12768)
);

OAI22xp5_ASAP7_75t_SL g12769 ( 
.A1(n_11872),
.A2(n_1327),
.B1(n_1325),
.B2(n_1326),
.Y(n_12769)
);

INVx1_ASAP7_75t_L g12770 ( 
.A(n_12431),
.Y(n_12770)
);

INVx1_ASAP7_75t_L g12771 ( 
.A(n_12440),
.Y(n_12771)
);

NOR2xp33_ASAP7_75t_SL g12772 ( 
.A(n_11740),
.B(n_1326),
.Y(n_12772)
);

OAI221xp5_ASAP7_75t_L g12773 ( 
.A1(n_12413),
.A2(n_12472),
.B1(n_12332),
.B2(n_12394),
.C(n_12428),
.Y(n_12773)
);

INVx2_ASAP7_75t_L g12774 ( 
.A(n_12441),
.Y(n_12774)
);

NAND2xp5_ASAP7_75t_L g12775 ( 
.A(n_12467),
.B(n_1327),
.Y(n_12775)
);

AND2x2_ASAP7_75t_L g12776 ( 
.A(n_11626),
.B(n_1328),
.Y(n_12776)
);

CKINVDCx14_ASAP7_75t_R g12777 ( 
.A(n_12498),
.Y(n_12777)
);

AOI22xp5_ASAP7_75t_L g12778 ( 
.A1(n_11834),
.A2(n_1330),
.B1(n_1328),
.B2(n_1329),
.Y(n_12778)
);

OAI22xp5_ASAP7_75t_L g12779 ( 
.A1(n_11612),
.A2(n_11669),
.B1(n_11673),
.B2(n_11665),
.Y(n_12779)
);

INVxp67_ASAP7_75t_L g12780 ( 
.A(n_11786),
.Y(n_12780)
);

AND2x2_ASAP7_75t_L g12781 ( 
.A(n_12334),
.B(n_1331),
.Y(n_12781)
);

NAND2xp5_ASAP7_75t_L g12782 ( 
.A(n_12471),
.B(n_12474),
.Y(n_12782)
);

NAND2xp5_ASAP7_75t_SL g12783 ( 
.A(n_12288),
.B(n_12200),
.Y(n_12783)
);

NAND2xp5_ASAP7_75t_L g12784 ( 
.A(n_12479),
.B(n_1331),
.Y(n_12784)
);

AND2x2_ASAP7_75t_L g12785 ( 
.A(n_12352),
.B(n_12489),
.Y(n_12785)
);

OR2x2_ASAP7_75t_L g12786 ( 
.A(n_12483),
.B(n_1332),
.Y(n_12786)
);

CKINVDCx5p33_ASAP7_75t_R g12787 ( 
.A(n_12327),
.Y(n_12787)
);

INVx2_ASAP7_75t_L g12788 ( 
.A(n_12496),
.Y(n_12788)
);

OAI22xp5_ASAP7_75t_SL g12789 ( 
.A1(n_11872),
.A2(n_1334),
.B1(n_1332),
.B2(n_1333),
.Y(n_12789)
);

AOI22xp33_ASAP7_75t_L g12790 ( 
.A1(n_12021),
.A2(n_1335),
.B1(n_1333),
.B2(n_1334),
.Y(n_12790)
);

CKINVDCx5p33_ASAP7_75t_R g12791 ( 
.A(n_12335),
.Y(n_12791)
);

AND3x1_ASAP7_75t_SL g12792 ( 
.A(n_12353),
.B(n_1335),
.C(n_1336),
.Y(n_12792)
);

INVx4_ASAP7_75t_L g12793 ( 
.A(n_11875),
.Y(n_12793)
);

INVx2_ASAP7_75t_L g12794 ( 
.A(n_12267),
.Y(n_12794)
);

AND2x2_ASAP7_75t_L g12795 ( 
.A(n_12500),
.B(n_1336),
.Y(n_12795)
);

BUFx6f_ASAP7_75t_L g12796 ( 
.A(n_12335),
.Y(n_12796)
);

AND2x2_ASAP7_75t_L g12797 ( 
.A(n_11721),
.B(n_12373),
.Y(n_12797)
);

INVx1_ASAP7_75t_L g12798 ( 
.A(n_11827),
.Y(n_12798)
);

AND2x2_ASAP7_75t_L g12799 ( 
.A(n_12376),
.B(n_1337),
.Y(n_12799)
);

NAND2xp5_ASAP7_75t_L g12800 ( 
.A(n_12229),
.B(n_1337),
.Y(n_12800)
);

NAND2xp5_ASAP7_75t_L g12801 ( 
.A(n_12135),
.B(n_1338),
.Y(n_12801)
);

NAND2xp5_ASAP7_75t_L g12802 ( 
.A(n_12140),
.B(n_1338),
.Y(n_12802)
);

AOI22xp33_ASAP7_75t_L g12803 ( 
.A1(n_11702),
.A2(n_1341),
.B1(n_1339),
.B2(n_1340),
.Y(n_12803)
);

BUFx3_ASAP7_75t_L g12804 ( 
.A(n_12362),
.Y(n_12804)
);

NAND2xp5_ASAP7_75t_L g12805 ( 
.A(n_12142),
.B(n_1339),
.Y(n_12805)
);

AOI22xp33_ASAP7_75t_L g12806 ( 
.A1(n_11650),
.A2(n_11670),
.B1(n_11672),
.B2(n_11658),
.Y(n_12806)
);

NAND2xp5_ASAP7_75t_L g12807 ( 
.A(n_11746),
.B(n_1341),
.Y(n_12807)
);

INVx2_ASAP7_75t_L g12808 ( 
.A(n_12279),
.Y(n_12808)
);

NAND2xp5_ASAP7_75t_L g12809 ( 
.A(n_11749),
.B(n_1342),
.Y(n_12809)
);

CKINVDCx20_ASAP7_75t_R g12810 ( 
.A(n_12194),
.Y(n_12810)
);

INVx3_ASAP7_75t_L g12811 ( 
.A(n_11900),
.Y(n_12811)
);

INVx2_ASAP7_75t_L g12812 ( 
.A(n_11734),
.Y(n_12812)
);

NAND2xp5_ASAP7_75t_L g12813 ( 
.A(n_11754),
.B(n_1343),
.Y(n_12813)
);

INVx1_ASAP7_75t_L g12814 ( 
.A(n_11788),
.Y(n_12814)
);

AND2x2_ASAP7_75t_L g12815 ( 
.A(n_12407),
.B(n_1343),
.Y(n_12815)
);

NAND2xp33_ASAP7_75t_L g12816 ( 
.A(n_12255),
.B(n_1344),
.Y(n_12816)
);

NAND2xp5_ASAP7_75t_L g12817 ( 
.A(n_11766),
.B(n_1344),
.Y(n_12817)
);

CKINVDCx6p67_ASAP7_75t_R g12818 ( 
.A(n_12323),
.Y(n_12818)
);

INVx2_ASAP7_75t_L g12819 ( 
.A(n_11791),
.Y(n_12819)
);

INVx1_ASAP7_75t_L g12820 ( 
.A(n_11789),
.Y(n_12820)
);

INVx1_ASAP7_75t_L g12821 ( 
.A(n_11794),
.Y(n_12821)
);

NAND2xp5_ASAP7_75t_L g12822 ( 
.A(n_11772),
.B(n_1345),
.Y(n_12822)
);

OR2x2_ASAP7_75t_L g12823 ( 
.A(n_11623),
.B(n_1345),
.Y(n_12823)
);

NAND2xp5_ASAP7_75t_L g12824 ( 
.A(n_11634),
.B(n_1346),
.Y(n_12824)
);

NAND2xp5_ASAP7_75t_L g12825 ( 
.A(n_11635),
.B(n_11636),
.Y(n_12825)
);

NAND2xp5_ASAP7_75t_SL g12826 ( 
.A(n_12288),
.B(n_11698),
.Y(n_12826)
);

AND2x4_ASAP7_75t_L g12827 ( 
.A(n_11989),
.B(n_1346),
.Y(n_12827)
);

OR2x2_ASAP7_75t_L g12828 ( 
.A(n_11637),
.B(n_1347),
.Y(n_12828)
);

NAND2xp5_ASAP7_75t_L g12829 ( 
.A(n_11773),
.B(n_1347),
.Y(n_12829)
);

INVx1_ASAP7_75t_L g12830 ( 
.A(n_11796),
.Y(n_12830)
);

AOI22xp5_ASAP7_75t_L g12831 ( 
.A1(n_11955),
.A2(n_1350),
.B1(n_1348),
.B2(n_1349),
.Y(n_12831)
);

INVx1_ASAP7_75t_L g12832 ( 
.A(n_11799),
.Y(n_12832)
);

NAND2xp5_ASAP7_75t_SL g12833 ( 
.A(n_11643),
.B(n_1348),
.Y(n_12833)
);

A2O1A1Ixp33_ASAP7_75t_L g12834 ( 
.A1(n_11958),
.A2(n_1352),
.B(n_1349),
.C(n_1351),
.Y(n_12834)
);

OAI21xp5_ASAP7_75t_L g12835 ( 
.A1(n_12319),
.A2(n_1351),
.B(n_1352),
.Y(n_12835)
);

NAND2xp5_ASAP7_75t_L g12836 ( 
.A(n_11608),
.B(n_1353),
.Y(n_12836)
);

NAND2x1p5_ASAP7_75t_L g12837 ( 
.A(n_11845),
.B(n_1353),
.Y(n_12837)
);

INVx1_ASAP7_75t_L g12838 ( 
.A(n_11802),
.Y(n_12838)
);

NAND2x1p5_ASAP7_75t_L g12839 ( 
.A(n_11861),
.B(n_1354),
.Y(n_12839)
);

OR2x2_ASAP7_75t_L g12840 ( 
.A(n_11639),
.B(n_1354),
.Y(n_12840)
);

NAND2xp5_ASAP7_75t_L g12841 ( 
.A(n_11638),
.B(n_1355),
.Y(n_12841)
);

A2O1A1Ixp33_ASAP7_75t_L g12842 ( 
.A1(n_11894),
.A2(n_1357),
.B(n_1355),
.C(n_1356),
.Y(n_12842)
);

INVxp67_ASAP7_75t_L g12843 ( 
.A(n_11674),
.Y(n_12843)
);

NAND2xp5_ASAP7_75t_L g12844 ( 
.A(n_12330),
.B(n_1356),
.Y(n_12844)
);

NAND2x1p5_ASAP7_75t_L g12845 ( 
.A(n_11862),
.B(n_1357),
.Y(n_12845)
);

NAND2xp5_ASAP7_75t_L g12846 ( 
.A(n_12340),
.B(n_12349),
.Y(n_12846)
);

AND2x4_ASAP7_75t_L g12847 ( 
.A(n_11628),
.B(n_1358),
.Y(n_12847)
);

INVx1_ASAP7_75t_L g12848 ( 
.A(n_11811),
.Y(n_12848)
);

INVx2_ASAP7_75t_L g12849 ( 
.A(n_11841),
.Y(n_12849)
);

CKINVDCx5p33_ASAP7_75t_R g12850 ( 
.A(n_12362),
.Y(n_12850)
);

OAI221xp5_ASAP7_75t_L g12851 ( 
.A1(n_12355),
.A2(n_1360),
.B1(n_1358),
.B2(n_1359),
.C(n_1361),
.Y(n_12851)
);

BUFx3_ASAP7_75t_L g12852 ( 
.A(n_12384),
.Y(n_12852)
);

BUFx2_ASAP7_75t_L g12853 ( 
.A(n_11850),
.Y(n_12853)
);

INVx2_ASAP7_75t_L g12854 ( 
.A(n_11912),
.Y(n_12854)
);

AND3x1_ASAP7_75t_SL g12855 ( 
.A(n_12378),
.B(n_1359),
.C(n_1360),
.Y(n_12855)
);

NAND2x1p5_ASAP7_75t_L g12856 ( 
.A(n_11988),
.B(n_1361),
.Y(n_12856)
);

NAND2xp5_ASAP7_75t_SL g12857 ( 
.A(n_12426),
.B(n_1362),
.Y(n_12857)
);

NAND2xp5_ASAP7_75t_L g12858 ( 
.A(n_12387),
.B(n_12419),
.Y(n_12858)
);

INVx1_ASAP7_75t_L g12859 ( 
.A(n_11820),
.Y(n_12859)
);

INVx2_ASAP7_75t_L g12860 ( 
.A(n_12010),
.Y(n_12860)
);

AOI22xp5_ASAP7_75t_L g12861 ( 
.A1(n_11710),
.A2(n_1364),
.B1(n_1362),
.B2(n_1363),
.Y(n_12861)
);

INVx2_ASAP7_75t_L g12862 ( 
.A(n_12015),
.Y(n_12862)
);

AND2x2_ASAP7_75t_L g12863 ( 
.A(n_12453),
.B(n_1363),
.Y(n_12863)
);

BUFx4f_ASAP7_75t_L g12864 ( 
.A(n_12384),
.Y(n_12864)
);

OAI22xp5_ASAP7_75t_L g12865 ( 
.A1(n_11829),
.A2(n_11769),
.B1(n_11695),
.B2(n_11904),
.Y(n_12865)
);

INVx2_ASAP7_75t_L g12866 ( 
.A(n_12052),
.Y(n_12866)
);

BUFx4f_ASAP7_75t_L g12867 ( 
.A(n_12390),
.Y(n_12867)
);

AND2x2_ASAP7_75t_L g12868 ( 
.A(n_12517),
.B(n_1364),
.Y(n_12868)
);

NAND2xp5_ASAP7_75t_L g12869 ( 
.A(n_12436),
.B(n_1365),
.Y(n_12869)
);

NAND2xp5_ASAP7_75t_L g12870 ( 
.A(n_12454),
.B(n_1365),
.Y(n_12870)
);

INVx3_ASAP7_75t_L g12871 ( 
.A(n_11915),
.Y(n_12871)
);

NOR3xp33_ASAP7_75t_L g12872 ( 
.A(n_11821),
.B(n_1366),
.C(n_1367),
.Y(n_12872)
);

OAI22xp5_ASAP7_75t_SL g12873 ( 
.A1(n_11911),
.A2(n_1368),
.B1(n_1366),
.B2(n_1367),
.Y(n_12873)
);

INVx1_ASAP7_75t_L g12874 ( 
.A(n_11840),
.Y(n_12874)
);

BUFx4f_ASAP7_75t_L g12875 ( 
.A(n_12390),
.Y(n_12875)
);

INVxp67_ASAP7_75t_L g12876 ( 
.A(n_11663),
.Y(n_12876)
);

NAND2xp5_ASAP7_75t_L g12877 ( 
.A(n_12470),
.B(n_1368),
.Y(n_12877)
);

NAND2xp5_ASAP7_75t_L g12878 ( 
.A(n_12497),
.B(n_1369),
.Y(n_12878)
);

INVx1_ASAP7_75t_L g12879 ( 
.A(n_11870),
.Y(n_12879)
);

OAI22xp5_ASAP7_75t_L g12880 ( 
.A1(n_11952),
.A2(n_1371),
.B1(n_1369),
.B2(n_1370),
.Y(n_12880)
);

INVx2_ASAP7_75t_L g12881 ( 
.A(n_11915),
.Y(n_12881)
);

NAND2xp5_ASAP7_75t_L g12882 ( 
.A(n_12501),
.B(n_12502),
.Y(n_12882)
);

A2O1A1Ixp33_ASAP7_75t_L g12883 ( 
.A1(n_11785),
.A2(n_1373),
.B(n_1370),
.C(n_1372),
.Y(n_12883)
);

AND2x2_ASAP7_75t_L g12884 ( 
.A(n_11727),
.B(n_1374),
.Y(n_12884)
);

INVx1_ASAP7_75t_L g12885 ( 
.A(n_11891),
.Y(n_12885)
);

INVx1_ASAP7_75t_L g12886 ( 
.A(n_11898),
.Y(n_12886)
);

NAND2xp5_ASAP7_75t_SL g12887 ( 
.A(n_12277),
.B(n_1375),
.Y(n_12887)
);

AND2x2_ASAP7_75t_L g12888 ( 
.A(n_12041),
.B(n_1376),
.Y(n_12888)
);

AND2x2_ASAP7_75t_L g12889 ( 
.A(n_11677),
.B(n_1376),
.Y(n_12889)
);

HB1xp67_ASAP7_75t_L g12890 ( 
.A(n_11913),
.Y(n_12890)
);

NAND2xp5_ASAP7_75t_L g12891 ( 
.A(n_12509),
.B(n_1377),
.Y(n_12891)
);

INVx1_ASAP7_75t_L g12892 ( 
.A(n_11919),
.Y(n_12892)
);

INVx1_ASAP7_75t_L g12893 ( 
.A(n_11933),
.Y(n_12893)
);

OR2x2_ASAP7_75t_L g12894 ( 
.A(n_11667),
.B(n_1377),
.Y(n_12894)
);

NAND2xp5_ASAP7_75t_L g12895 ( 
.A(n_12519),
.B(n_1378),
.Y(n_12895)
);

AND3x1_ASAP7_75t_SL g12896 ( 
.A(n_12381),
.B(n_1378),
.C(n_1379),
.Y(n_12896)
);

BUFx2_ASAP7_75t_L g12897 ( 
.A(n_11975),
.Y(n_12897)
);

AND2x2_ASAP7_75t_L g12898 ( 
.A(n_12312),
.B(n_1379),
.Y(n_12898)
);

AOI22xp5_ASAP7_75t_L g12899 ( 
.A1(n_12270),
.A2(n_1382),
.B1(n_1380),
.B2(n_1381),
.Y(n_12899)
);

INVx2_ASAP7_75t_L g12900 ( 
.A(n_11975),
.Y(n_12900)
);

CKINVDCx5p33_ASAP7_75t_R g12901 ( 
.A(n_12462),
.Y(n_12901)
);

INVx1_ASAP7_75t_L g12902 ( 
.A(n_11934),
.Y(n_12902)
);

OAI22xp5_ASAP7_75t_SL g12903 ( 
.A1(n_11801),
.A2(n_11808),
.B1(n_11972),
.B2(n_11973),
.Y(n_12903)
);

NAND2xp5_ASAP7_75t_L g12904 ( 
.A(n_11723),
.B(n_1380),
.Y(n_12904)
);

INVx1_ASAP7_75t_L g12905 ( 
.A(n_11941),
.Y(n_12905)
);

NOR2xp33_ASAP7_75t_SL g12906 ( 
.A(n_12422),
.B(n_1383),
.Y(n_12906)
);

NAND2xp5_ASAP7_75t_SL g12907 ( 
.A(n_12302),
.B(n_1384),
.Y(n_12907)
);

A2O1A1Ixp33_ASAP7_75t_L g12908 ( 
.A1(n_11782),
.A2(n_1386),
.B(n_1384),
.C(n_1385),
.Y(n_12908)
);

CKINVDCx5p33_ASAP7_75t_R g12909 ( 
.A(n_12462),
.Y(n_12909)
);

INVxp67_ASAP7_75t_L g12910 ( 
.A(n_11668),
.Y(n_12910)
);

INVx2_ASAP7_75t_L g12911 ( 
.A(n_11977),
.Y(n_12911)
);

AND2x4_ASAP7_75t_L g12912 ( 
.A(n_11737),
.B(n_1385),
.Y(n_12912)
);

INVx4_ASAP7_75t_L g12913 ( 
.A(n_11977),
.Y(n_12913)
);

NAND2xp5_ASAP7_75t_SL g12914 ( 
.A(n_11622),
.B(n_1386),
.Y(n_12914)
);

INVx1_ASAP7_75t_L g12915 ( 
.A(n_11944),
.Y(n_12915)
);

INVx1_ASAP7_75t_L g12916 ( 
.A(n_11956),
.Y(n_12916)
);

OAI22xp5_ASAP7_75t_L g12917 ( 
.A1(n_11909),
.A2(n_11914),
.B1(n_12488),
.B2(n_12446),
.Y(n_12917)
);

NOR2xp67_ASAP7_75t_L g12918 ( 
.A(n_11744),
.B(n_11770),
.Y(n_12918)
);

BUFx4f_ASAP7_75t_L g12919 ( 
.A(n_12508),
.Y(n_12919)
);

NAND2xp5_ASAP7_75t_L g12920 ( 
.A(n_11716),
.B(n_1387),
.Y(n_12920)
);

NAND2xp5_ASAP7_75t_L g12921 ( 
.A(n_12219),
.B(n_1388),
.Y(n_12921)
);

NAND2xp5_ASAP7_75t_L g12922 ( 
.A(n_11764),
.B(n_1388),
.Y(n_12922)
);

INVx1_ASAP7_75t_L g12923 ( 
.A(n_11963),
.Y(n_12923)
);

INVx2_ASAP7_75t_L g12924 ( 
.A(n_11966),
.Y(n_12924)
);

AND2x4_ASAP7_75t_L g12925 ( 
.A(n_12375),
.B(n_1389),
.Y(n_12925)
);

AND2x2_ASAP7_75t_L g12926 ( 
.A(n_12465),
.B(n_1389),
.Y(n_12926)
);

INVx2_ASAP7_75t_L g12927 ( 
.A(n_11971),
.Y(n_12927)
);

AND2x2_ASAP7_75t_L g12928 ( 
.A(n_12006),
.B(n_1390),
.Y(n_12928)
);

AND2x2_ASAP7_75t_L g12929 ( 
.A(n_11713),
.B(n_1390),
.Y(n_12929)
);

A2O1A1Ixp33_ASAP7_75t_L g12930 ( 
.A1(n_11733),
.A2(n_1393),
.B(n_1391),
.C(n_1392),
.Y(n_12930)
);

INVx1_ASAP7_75t_L g12931 ( 
.A(n_11993),
.Y(n_12931)
);

BUFx2_ASAP7_75t_L g12932 ( 
.A(n_12508),
.Y(n_12932)
);

OAI21x1_ASAP7_75t_L g12933 ( 
.A1(n_12216),
.A2(n_1391),
.B(n_1393),
.Y(n_12933)
);

NAND2xp5_ASAP7_75t_L g12934 ( 
.A(n_12253),
.B(n_1394),
.Y(n_12934)
);

INVx1_ASAP7_75t_L g12935 ( 
.A(n_12000),
.Y(n_12935)
);

INVx1_ASAP7_75t_L g12936 ( 
.A(n_12005),
.Y(n_12936)
);

INVx1_ASAP7_75t_L g12937 ( 
.A(n_12008),
.Y(n_12937)
);

INVx1_ASAP7_75t_L g12938 ( 
.A(n_12012),
.Y(n_12938)
);

AND2x2_ASAP7_75t_L g12939 ( 
.A(n_11648),
.B(n_1394),
.Y(n_12939)
);

AOI22xp33_ASAP7_75t_L g12940 ( 
.A1(n_12281),
.A2(n_11835),
.B1(n_11848),
.B2(n_11992),
.Y(n_12940)
);

INVx1_ASAP7_75t_L g12941 ( 
.A(n_12017),
.Y(n_12941)
);

INVx1_ASAP7_75t_L g12942 ( 
.A(n_12130),
.Y(n_12942)
);

NAND2xp5_ASAP7_75t_L g12943 ( 
.A(n_12022),
.B(n_1395),
.Y(n_12943)
);

NOR2xp33_ASAP7_75t_R g12944 ( 
.A(n_11807),
.B(n_1395),
.Y(n_12944)
);

NAND2xp5_ASAP7_75t_L g12945 ( 
.A(n_12025),
.B(n_1396),
.Y(n_12945)
);

INVx1_ASAP7_75t_L g12946 ( 
.A(n_12051),
.Y(n_12946)
);

INVxp67_ASAP7_75t_SL g12947 ( 
.A(n_12286),
.Y(n_12947)
);

NOR2xp33_ASAP7_75t_L g12948 ( 
.A(n_11817),
.B(n_1397),
.Y(n_12948)
);

AND2x2_ASAP7_75t_L g12949 ( 
.A(n_11728),
.B(n_1397),
.Y(n_12949)
);

AND2x2_ASAP7_75t_L g12950 ( 
.A(n_12244),
.B(n_1398),
.Y(n_12950)
);

INVx2_ASAP7_75t_L g12951 ( 
.A(n_11826),
.Y(n_12951)
);

INVx2_ASAP7_75t_L g12952 ( 
.A(n_11869),
.Y(n_12952)
);

OAI21xp5_ASAP7_75t_L g12953 ( 
.A1(n_12321),
.A2(n_12348),
.B(n_12344),
.Y(n_12953)
);

AND2x2_ASAP7_75t_L g12954 ( 
.A(n_12228),
.B(n_1398),
.Y(n_12954)
);

INVxp67_ASAP7_75t_L g12955 ( 
.A(n_11929),
.Y(n_12955)
);

OAI22xp5_ASAP7_75t_SL g12956 ( 
.A1(n_11960),
.A2(n_1401),
.B1(n_1399),
.B2(n_1400),
.Y(n_12956)
);

NAND2xp5_ASAP7_75t_L g12957 ( 
.A(n_12028),
.B(n_1399),
.Y(n_12957)
);

NOR2xp67_ASAP7_75t_L g12958 ( 
.A(n_12089),
.B(n_1400),
.Y(n_12958)
);

NAND2xp5_ASAP7_75t_L g12959 ( 
.A(n_12030),
.B(n_1401),
.Y(n_12959)
);

OAI22xp5_ASAP7_75t_SL g12960 ( 
.A1(n_11964),
.A2(n_12040),
.B1(n_11987),
.B2(n_12210),
.Y(n_12960)
);

AND2x2_ASAP7_75t_L g12961 ( 
.A(n_12085),
.B(n_1402),
.Y(n_12961)
);

AOI22xp33_ASAP7_75t_L g12962 ( 
.A1(n_11605),
.A2(n_1404),
.B1(n_1402),
.B2(n_1403),
.Y(n_12962)
);

NOR2xp33_ASAP7_75t_L g12963 ( 
.A(n_11851),
.B(n_1403),
.Y(n_12963)
);

INVx1_ASAP7_75t_SL g12964 ( 
.A(n_11819),
.Y(n_12964)
);

NAND2xp5_ASAP7_75t_SL g12965 ( 
.A(n_12191),
.B(n_1404),
.Y(n_12965)
);

NOR2xp33_ASAP7_75t_L g12966 ( 
.A(n_12240),
.B(n_1405),
.Y(n_12966)
);

AOI22xp33_ASAP7_75t_SL g12967 ( 
.A1(n_11843),
.A2(n_1407),
.B1(n_1405),
.B2(n_1406),
.Y(n_12967)
);

INVx2_ASAP7_75t_L g12968 ( 
.A(n_11947),
.Y(n_12968)
);

INVx3_ASAP7_75t_L g12969 ( 
.A(n_11981),
.Y(n_12969)
);

INVx2_ASAP7_75t_L g12970 ( 
.A(n_11844),
.Y(n_12970)
);

OAI22xp5_ASAP7_75t_L g12971 ( 
.A1(n_11818),
.A2(n_1409),
.B1(n_1406),
.B2(n_1408),
.Y(n_12971)
);

BUFx8_ASAP7_75t_L g12972 ( 
.A(n_12126),
.Y(n_12972)
);

NAND2xp5_ASAP7_75t_L g12973 ( 
.A(n_12038),
.B(n_1408),
.Y(n_12973)
);

INVx3_ASAP7_75t_L g12974 ( 
.A(n_11797),
.Y(n_12974)
);

NAND2x1p5_ASAP7_75t_L g12975 ( 
.A(n_12293),
.B(n_11694),
.Y(n_12975)
);

OAI22xp5_ASAP7_75t_SL g12976 ( 
.A1(n_12175),
.A2(n_1411),
.B1(n_1409),
.B2(n_1410),
.Y(n_12976)
);

AND2x2_ASAP7_75t_L g12977 ( 
.A(n_12108),
.B(n_1410),
.Y(n_12977)
);

CKINVDCx5p33_ASAP7_75t_R g12978 ( 
.A(n_12237),
.Y(n_12978)
);

NAND2xp5_ASAP7_75t_SL g12979 ( 
.A(n_12259),
.B(n_1412),
.Y(n_12979)
);

NAND2xp5_ASAP7_75t_L g12980 ( 
.A(n_12047),
.B(n_1412),
.Y(n_12980)
);

INVx2_ASAP7_75t_SL g12981 ( 
.A(n_12043),
.Y(n_12981)
);

AND2x2_ASAP7_75t_L g12982 ( 
.A(n_12113),
.B(n_12121),
.Y(n_12982)
);

NAND2xp5_ASAP7_75t_L g12983 ( 
.A(n_12050),
.B(n_1413),
.Y(n_12983)
);

AND2x6_ASAP7_75t_L g12984 ( 
.A(n_12296),
.B(n_1413),
.Y(n_12984)
);

NAND3xp33_ASAP7_75t_SL g12985 ( 
.A(n_11997),
.B(n_1414),
.C(n_1415),
.Y(n_12985)
);

AOI22xp5_ASAP7_75t_L g12986 ( 
.A1(n_11831),
.A2(n_1417),
.B1(n_1415),
.B2(n_1416),
.Y(n_12986)
);

INVx1_ASAP7_75t_L g12987 ( 
.A(n_11980),
.Y(n_12987)
);

INVx3_ASAP7_75t_L g12988 ( 
.A(n_12126),
.Y(n_12988)
);

INVx2_ASAP7_75t_L g12989 ( 
.A(n_12342),
.Y(n_12989)
);

BUFx6f_ASAP7_75t_L g12990 ( 
.A(n_12160),
.Y(n_12990)
);

AND3x1_ASAP7_75t_SL g12991 ( 
.A(n_11858),
.B(n_1418),
.C(n_1419),
.Y(n_12991)
);

AND2x2_ASAP7_75t_L g12992 ( 
.A(n_12187),
.B(n_1419),
.Y(n_12992)
);

OR2x6_ASAP7_75t_SL g12993 ( 
.A(n_11729),
.B(n_1420),
.Y(n_12993)
);

NAND2x1p5_ASAP7_75t_L g12994 ( 
.A(n_11714),
.B(n_1421),
.Y(n_12994)
);

BUFx6f_ASAP7_75t_L g12995 ( 
.A(n_12183),
.Y(n_12995)
);

NAND2xp5_ASAP7_75t_L g12996 ( 
.A(n_12076),
.B(n_1421),
.Y(n_12996)
);

NAND2xp5_ASAP7_75t_L g12997 ( 
.A(n_12090),
.B(n_12092),
.Y(n_12997)
);

INVx1_ASAP7_75t_L g12998 ( 
.A(n_11775),
.Y(n_12998)
);

AOI22xp5_ASAP7_75t_L g12999 ( 
.A1(n_11692),
.A2(n_11646),
.B1(n_12109),
.B2(n_12300),
.Y(n_12999)
);

NAND2xp5_ASAP7_75t_L g13000 ( 
.A(n_12093),
.B(n_1422),
.Y(n_13000)
);

AOI22xp5_ASAP7_75t_L g13001 ( 
.A1(n_12180),
.A2(n_1424),
.B1(n_1422),
.B2(n_1423),
.Y(n_13001)
);

NAND2xp5_ASAP7_75t_SL g13002 ( 
.A(n_11923),
.B(n_12360),
.Y(n_13002)
);

AND2x2_ASAP7_75t_L g13003 ( 
.A(n_12205),
.B(n_1423),
.Y(n_13003)
);

NAND2xp5_ASAP7_75t_L g13004 ( 
.A(n_12118),
.B(n_1424),
.Y(n_13004)
);

INVx1_ASAP7_75t_L g13005 ( 
.A(n_11950),
.Y(n_13005)
);

NAND2xp5_ASAP7_75t_L g13006 ( 
.A(n_12127),
.B(n_1425),
.Y(n_13006)
);

NAND2xp5_ASAP7_75t_L g13007 ( 
.A(n_12134),
.B(n_1425),
.Y(n_13007)
);

OAI22xp5_ASAP7_75t_SL g13008 ( 
.A1(n_11884),
.A2(n_1428),
.B1(n_1426),
.B2(n_1427),
.Y(n_13008)
);

HB1xp67_ASAP7_75t_L g13009 ( 
.A(n_12271),
.Y(n_13009)
);

AO22x1_ASAP7_75t_L g13010 ( 
.A1(n_12126),
.A2(n_1429),
.B1(n_1426),
.B2(n_1428),
.Y(n_13010)
);

AND2x2_ASAP7_75t_L g13011 ( 
.A(n_11760),
.B(n_11877),
.Y(n_13011)
);

INVx2_ASAP7_75t_L g13012 ( 
.A(n_11752),
.Y(n_13012)
);

INVx2_ASAP7_75t_L g13013 ( 
.A(n_11787),
.Y(n_13013)
);

NAND2xp5_ASAP7_75t_L g13014 ( 
.A(n_12138),
.B(n_1429),
.Y(n_13014)
);

INVxp67_ASAP7_75t_L g13015 ( 
.A(n_12147),
.Y(n_13015)
);

NOR2xp33_ASAP7_75t_L g13016 ( 
.A(n_12242),
.B(n_1430),
.Y(n_13016)
);

NAND2xp5_ASAP7_75t_L g13017 ( 
.A(n_12150),
.B(n_1430),
.Y(n_13017)
);

AND2x2_ASAP7_75t_L g13018 ( 
.A(n_11892),
.B(n_1431),
.Y(n_13018)
);

NAND2xp5_ASAP7_75t_L g13019 ( 
.A(n_12151),
.B(n_1431),
.Y(n_13019)
);

BUFx6f_ASAP7_75t_L g13020 ( 
.A(n_12169),
.Y(n_13020)
);

NAND2xp5_ASAP7_75t_L g13021 ( 
.A(n_12152),
.B(n_1432),
.Y(n_13021)
);

AND2x4_ASAP7_75t_L g13022 ( 
.A(n_12169),
.B(n_1432),
.Y(n_13022)
);

AND3x1_ASAP7_75t_SL g13023 ( 
.A(n_12455),
.B(n_1433),
.C(n_1434),
.Y(n_13023)
);

AND2x2_ASAP7_75t_L g13024 ( 
.A(n_11899),
.B(n_1433),
.Y(n_13024)
);

NAND2xp5_ASAP7_75t_L g13025 ( 
.A(n_12155),
.B(n_1434),
.Y(n_13025)
);

NAND2xp5_ASAP7_75t_L g13026 ( 
.A(n_12156),
.B(n_1435),
.Y(n_13026)
);

BUFx4f_ASAP7_75t_L g13027 ( 
.A(n_12178),
.Y(n_13027)
);

AND2x2_ASAP7_75t_L g13028 ( 
.A(n_11902),
.B(n_1435),
.Y(n_13028)
);

NAND2xp5_ASAP7_75t_L g13029 ( 
.A(n_12158),
.B(n_1436),
.Y(n_13029)
);

NAND2xp5_ASAP7_75t_L g13030 ( 
.A(n_12164),
.B(n_1436),
.Y(n_13030)
);

CKINVDCx20_ASAP7_75t_R g13031 ( 
.A(n_11735),
.Y(n_13031)
);

BUFx2_ASAP7_75t_L g13032 ( 
.A(n_12303),
.Y(n_13032)
);

AOI22xp33_ASAP7_75t_L g13033 ( 
.A1(n_11836),
.A2(n_1439),
.B1(n_1437),
.B2(n_1438),
.Y(n_13033)
);

INVx2_ASAP7_75t_L g13034 ( 
.A(n_12059),
.Y(n_13034)
);

INVxp67_ASAP7_75t_L g13035 ( 
.A(n_12245),
.Y(n_13035)
);

INVx1_ASAP7_75t_L g13036 ( 
.A(n_12310),
.Y(n_13036)
);

NOR2xp33_ASAP7_75t_R g13037 ( 
.A(n_12491),
.B(n_1437),
.Y(n_13037)
);

INVx2_ASAP7_75t_L g13038 ( 
.A(n_11996),
.Y(n_13038)
);

NAND2xp5_ASAP7_75t_L g13039 ( 
.A(n_12170),
.B(n_1439),
.Y(n_13039)
);

AND3x1_ASAP7_75t_SL g13040 ( 
.A(n_11837),
.B(n_1440),
.C(n_1441),
.Y(n_13040)
);

NOR2xp33_ASAP7_75t_L g13041 ( 
.A(n_11999),
.B(n_1440),
.Y(n_13041)
);

AND2x2_ASAP7_75t_L g13042 ( 
.A(n_11759),
.B(n_1442),
.Y(n_13042)
);

OAI21x1_ASAP7_75t_L g13043 ( 
.A1(n_12024),
.A2(n_1442),
.B(n_1443),
.Y(n_13043)
);

NAND2xp5_ASAP7_75t_L g13044 ( 
.A(n_12192),
.B(n_1443),
.Y(n_13044)
);

AND2x2_ASAP7_75t_L g13045 ( 
.A(n_11978),
.B(n_1444),
.Y(n_13045)
);

OAI22xp5_ASAP7_75t_L g13046 ( 
.A1(n_11968),
.A2(n_1446),
.B1(n_1444),
.B2(n_1445),
.Y(n_13046)
);

HB1xp67_ASAP7_75t_L g13047 ( 
.A(n_12328),
.Y(n_13047)
);

INVx2_ASAP7_75t_L g13048 ( 
.A(n_11825),
.Y(n_13048)
);

OAI22xp5_ASAP7_75t_L g13049 ( 
.A1(n_11781),
.A2(n_1448),
.B1(n_1446),
.B2(n_1447),
.Y(n_13049)
);

INVxp33_ASAP7_75t_L g13050 ( 
.A(n_12065),
.Y(n_13050)
);

NAND2xp5_ASAP7_75t_L g13051 ( 
.A(n_12195),
.B(n_1447),
.Y(n_13051)
);

OAI22xp5_ASAP7_75t_SL g13052 ( 
.A1(n_11908),
.A2(n_1450),
.B1(n_1448),
.B2(n_1449),
.Y(n_13052)
);

NAND2xp5_ASAP7_75t_SL g13053 ( 
.A(n_12317),
.B(n_1449),
.Y(n_13053)
);

BUFx3_ASAP7_75t_L g13054 ( 
.A(n_11678),
.Y(n_13054)
);

INVx2_ASAP7_75t_L g13055 ( 
.A(n_12410),
.Y(n_13055)
);

INVx2_ASAP7_75t_L g13056 ( 
.A(n_11984),
.Y(n_13056)
);

INVx3_ASAP7_75t_L g13057 ( 
.A(n_12178),
.Y(n_13057)
);

BUFx3_ASAP7_75t_L g13058 ( 
.A(n_11679),
.Y(n_13058)
);

INVx2_ASAP7_75t_L g13059 ( 
.A(n_12282),
.Y(n_13059)
);

INVx1_ASAP7_75t_L g13060 ( 
.A(n_12001),
.Y(n_13060)
);

NAND2xp5_ASAP7_75t_L g13061 ( 
.A(n_12196),
.B(n_1450),
.Y(n_13061)
);

AND2x2_ASAP7_75t_L g13062 ( 
.A(n_11701),
.B(n_1451),
.Y(n_13062)
);

HB1xp67_ASAP7_75t_L g13063 ( 
.A(n_11901),
.Y(n_13063)
);

OAI22xp5_ASAP7_75t_SL g13064 ( 
.A1(n_12168),
.A2(n_1453),
.B1(n_1451),
.B2(n_1452),
.Y(n_13064)
);

NAND2xp5_ASAP7_75t_L g13065 ( 
.A(n_12202),
.B(n_1452),
.Y(n_13065)
);

INVx2_ASAP7_75t_L g13066 ( 
.A(n_12289),
.Y(n_13066)
);

NAND2x1p5_ASAP7_75t_L g13067 ( 
.A(n_11724),
.B(n_1453),
.Y(n_13067)
);

INVx2_ASAP7_75t_L g13068 ( 
.A(n_12206),
.Y(n_13068)
);

INVx1_ASAP7_75t_L g13069 ( 
.A(n_12001),
.Y(n_13069)
);

OAI21xp5_ASAP7_75t_L g13070 ( 
.A1(n_12350),
.A2(n_1454),
.B(n_1455),
.Y(n_13070)
);

NAND2xp5_ASAP7_75t_L g13071 ( 
.A(n_12212),
.B(n_1455),
.Y(n_13071)
);

INVx1_ASAP7_75t_L g13072 ( 
.A(n_12013),
.Y(n_13072)
);

BUFx6f_ASAP7_75t_L g13073 ( 
.A(n_11709),
.Y(n_13073)
);

CKINVDCx5p33_ASAP7_75t_R g13074 ( 
.A(n_12174),
.Y(n_13074)
);

NAND2xp5_ASAP7_75t_L g13075 ( 
.A(n_12215),
.B(n_1456),
.Y(n_13075)
);

INVx2_ASAP7_75t_L g13076 ( 
.A(n_12220),
.Y(n_13076)
);

INVx1_ASAP7_75t_L g13077 ( 
.A(n_11725),
.Y(n_13077)
);

INVx2_ASAP7_75t_L g13078 ( 
.A(n_12238),
.Y(n_13078)
);

INVxp33_ASAP7_75t_SL g13079 ( 
.A(n_12079),
.Y(n_13079)
);

INVx2_ASAP7_75t_L g13080 ( 
.A(n_12239),
.Y(n_13080)
);

NAND2xp5_ASAP7_75t_L g13081 ( 
.A(n_12243),
.B(n_1456),
.Y(n_13081)
);

CKINVDCx5p33_ASAP7_75t_R g13082 ( 
.A(n_12101),
.Y(n_13082)
);

INVx1_ASAP7_75t_L g13083 ( 
.A(n_11725),
.Y(n_13083)
);

INVx1_ASAP7_75t_L g13084 ( 
.A(n_12456),
.Y(n_13084)
);

INVx1_ASAP7_75t_L g13085 ( 
.A(n_12456),
.Y(n_13085)
);

NAND2xp5_ASAP7_75t_L g13086 ( 
.A(n_12148),
.B(n_1457),
.Y(n_13086)
);

INVx1_ASAP7_75t_L g13087 ( 
.A(n_11889),
.Y(n_13087)
);

NAND2xp5_ASAP7_75t_L g13088 ( 
.A(n_12341),
.B(n_12361),
.Y(n_13088)
);

NAND2xp5_ASAP7_75t_L g13089 ( 
.A(n_12369),
.B(n_1457),
.Y(n_13089)
);

AOI22xp33_ASAP7_75t_L g13090 ( 
.A1(n_11890),
.A2(n_1460),
.B1(n_1458),
.B2(n_1459),
.Y(n_13090)
);

CKINVDCx5p33_ASAP7_75t_R g13091 ( 
.A(n_12129),
.Y(n_13091)
);

NAND2xp5_ASAP7_75t_L g13092 ( 
.A(n_12372),
.B(n_1458),
.Y(n_13092)
);

INVx2_ASAP7_75t_L g13093 ( 
.A(n_11651),
.Y(n_13093)
);

CKINVDCx5p33_ASAP7_75t_R g13094 ( 
.A(n_12163),
.Y(n_13094)
);

OAI21x1_ASAP7_75t_L g13095 ( 
.A1(n_11741),
.A2(n_1459),
.B(n_1460),
.Y(n_13095)
);

HB1xp67_ASAP7_75t_L g13096 ( 
.A(n_11901),
.Y(n_13096)
);

NAND2xp5_ASAP7_75t_L g13097 ( 
.A(n_12379),
.B(n_1461),
.Y(n_13097)
);

NAND2xp5_ASAP7_75t_L g13098 ( 
.A(n_12392),
.B(n_1462),
.Y(n_13098)
);

NAND2xp5_ASAP7_75t_L g13099 ( 
.A(n_12447),
.B(n_1463),
.Y(n_13099)
);

AND3x1_ASAP7_75t_SL g13100 ( 
.A(n_11666),
.B(n_1463),
.C(n_1464),
.Y(n_13100)
);

INVx2_ASAP7_75t_L g13101 ( 
.A(n_12268),
.Y(n_13101)
);

NAND2xp5_ASAP7_75t_L g13102 ( 
.A(n_12477),
.B(n_1464),
.Y(n_13102)
);

INVx3_ASAP7_75t_L g13103 ( 
.A(n_12287),
.Y(n_13103)
);

BUFx2_ASAP7_75t_L g13104 ( 
.A(n_11906),
.Y(n_13104)
);

INVx1_ASAP7_75t_L g13105 ( 
.A(n_11765),
.Y(n_13105)
);

NAND2xp5_ASAP7_75t_SL g13106 ( 
.A(n_12490),
.B(n_1465),
.Y(n_13106)
);

INVx1_ASAP7_75t_L g13107 ( 
.A(n_12499),
.Y(n_13107)
);

NAND2xp5_ASAP7_75t_L g13108 ( 
.A(n_12505),
.B(n_1465),
.Y(n_13108)
);

INVx2_ASAP7_75t_L g13109 ( 
.A(n_11682),
.Y(n_13109)
);

INVx2_ASAP7_75t_L g13110 ( 
.A(n_12516),
.Y(n_13110)
);

A2O1A1Ixp33_ASAP7_75t_L g13111 ( 
.A1(n_11696),
.A2(n_1468),
.B(n_1466),
.C(n_1467),
.Y(n_13111)
);

AOI22xp5_ASAP7_75t_L g13112 ( 
.A1(n_12231),
.A2(n_1470),
.B1(n_1468),
.B2(n_1469),
.Y(n_13112)
);

INVx2_ASAP7_75t_L g13113 ( 
.A(n_12298),
.Y(n_13113)
);

NAND2xp5_ASAP7_75t_L g13114 ( 
.A(n_12072),
.B(n_1469),
.Y(n_13114)
);

AND2x2_ASAP7_75t_SL g13115 ( 
.A(n_12171),
.B(n_1471),
.Y(n_13115)
);

INVx1_ASAP7_75t_L g13116 ( 
.A(n_12167),
.Y(n_13116)
);

NAND2xp5_ASAP7_75t_L g13117 ( 
.A(n_12074),
.B(n_1471),
.Y(n_13117)
);

NOR2xp33_ASAP7_75t_R g13118 ( 
.A(n_12248),
.B(n_1472),
.Y(n_13118)
);

INVx4_ASAP7_75t_L g13119 ( 
.A(n_12287),
.Y(n_13119)
);

INVxp67_ASAP7_75t_L g13120 ( 
.A(n_12265),
.Y(n_13120)
);

NAND2xp5_ASAP7_75t_L g13121 ( 
.A(n_12141),
.B(n_12354),
.Y(n_13121)
);

INVx1_ASAP7_75t_L g13122 ( 
.A(n_12292),
.Y(n_13122)
);

NAND2xp5_ASAP7_75t_SL g13123 ( 
.A(n_11965),
.B(n_1472),
.Y(n_13123)
);

NAND2xp5_ASAP7_75t_L g13124 ( 
.A(n_12356),
.B(n_1473),
.Y(n_13124)
);

INVx2_ASAP7_75t_L g13125 ( 
.A(n_11906),
.Y(n_13125)
);

AND2x4_ASAP7_75t_L g13126 ( 
.A(n_12091),
.B(n_12115),
.Y(n_13126)
);

OAI21x1_ASAP7_75t_L g13127 ( 
.A1(n_12184),
.A2(n_1474),
.B(n_1475),
.Y(n_13127)
);

AOI22xp33_ASAP7_75t_L g13128 ( 
.A1(n_12039),
.A2(n_1478),
.B1(n_1476),
.B2(n_1477),
.Y(n_13128)
);

INVx1_ASAP7_75t_L g13129 ( 
.A(n_12294),
.Y(n_13129)
);

BUFx6f_ASAP7_75t_L g13130 ( 
.A(n_12189),
.Y(n_13130)
);

AND2x4_ASAP7_75t_L g13131 ( 
.A(n_11803),
.B(n_1477),
.Y(n_13131)
);

INVx1_ASAP7_75t_L g13132 ( 
.A(n_12225),
.Y(n_13132)
);

OAI21xp5_ASAP7_75t_L g13133 ( 
.A1(n_12358),
.A2(n_1478),
.B(n_1479),
.Y(n_13133)
);

CKINVDCx12_ASAP7_75t_R g13134 ( 
.A(n_12176),
.Y(n_13134)
);

OAI22xp5_ASAP7_75t_L g13135 ( 
.A1(n_11867),
.A2(n_1482),
.B1(n_1480),
.B2(n_1481),
.Y(n_13135)
);

NAND3xp33_ASAP7_75t_SL g13136 ( 
.A(n_12383),
.B(n_1480),
.C(n_1481),
.Y(n_13136)
);

NAND2xp5_ASAP7_75t_L g13137 ( 
.A(n_12363),
.B(n_1482),
.Y(n_13137)
);

NOR3xp33_ASAP7_75t_L g13138 ( 
.A(n_12049),
.B(n_1483),
.C(n_1484),
.Y(n_13138)
);

OAI22xp5_ASAP7_75t_L g13139 ( 
.A1(n_11903),
.A2(n_1485),
.B1(n_1483),
.B2(n_1484),
.Y(n_13139)
);

AND2x2_ASAP7_75t_L g13140 ( 
.A(n_12197),
.B(n_1486),
.Y(n_13140)
);

INVx1_ASAP7_75t_L g13141 ( 
.A(n_12225),
.Y(n_13141)
);

AOI22xp5_ASAP7_75t_L g13142 ( 
.A1(n_11998),
.A2(n_1488),
.B1(n_1486),
.B2(n_1487),
.Y(n_13142)
);

AOI21xp5_ASAP7_75t_L g13143 ( 
.A1(n_12276),
.A2(n_1487),
.B(n_1488),
.Y(n_13143)
);

NAND2xp5_ASAP7_75t_L g13144 ( 
.A(n_12365),
.B(n_1489),
.Y(n_13144)
);

INVx2_ASAP7_75t_L g13145 ( 
.A(n_11931),
.Y(n_13145)
);

AOI22xp5_ASAP7_75t_L g13146 ( 
.A1(n_11632),
.A2(n_1491),
.B1(n_1489),
.B2(n_1490),
.Y(n_13146)
);

INVx1_ASAP7_75t_L g13147 ( 
.A(n_12190),
.Y(n_13147)
);

NAND2xp5_ASAP7_75t_L g13148 ( 
.A(n_12371),
.B(n_1491),
.Y(n_13148)
);

AND2x2_ASAP7_75t_L g13149 ( 
.A(n_12209),
.B(n_1492),
.Y(n_13149)
);

INVx1_ASAP7_75t_L g13150 ( 
.A(n_12190),
.Y(n_13150)
);

BUFx6f_ASAP7_75t_L g13151 ( 
.A(n_11878),
.Y(n_13151)
);

INVx1_ASAP7_75t_L g13152 ( 
.A(n_12048),
.Y(n_13152)
);

NAND2xp5_ASAP7_75t_L g13153 ( 
.A(n_12391),
.B(n_1492),
.Y(n_13153)
);

NAND2xp5_ASAP7_75t_L g13154 ( 
.A(n_12393),
.B(n_1493),
.Y(n_13154)
);

INVx1_ASAP7_75t_L g13155 ( 
.A(n_12173),
.Y(n_13155)
);

AOI22x1_ASAP7_75t_L g13156 ( 
.A1(n_12399),
.A2(n_1496),
.B1(n_1494),
.B2(n_1495),
.Y(n_13156)
);

AOI22xp33_ASAP7_75t_L g13157 ( 
.A1(n_12119),
.A2(n_1496),
.B1(n_1494),
.B2(n_1495),
.Y(n_13157)
);

INVx1_ASAP7_75t_L g13158 ( 
.A(n_12084),
.Y(n_13158)
);

INVx1_ASAP7_75t_L g13159 ( 
.A(n_12128),
.Y(n_13159)
);

INVx1_ASAP7_75t_L g13160 ( 
.A(n_12273),
.Y(n_13160)
);

INVx1_ASAP7_75t_L g13161 ( 
.A(n_11686),
.Y(n_13161)
);

NAND2xp5_ASAP7_75t_L g13162 ( 
.A(n_12411),
.B(n_1497),
.Y(n_13162)
);

CKINVDCx5p33_ASAP7_75t_R g13163 ( 
.A(n_11883),
.Y(n_13163)
);

INVx2_ASAP7_75t_L g13164 ( 
.A(n_11983),
.Y(n_13164)
);

AOI22xp5_ASAP7_75t_L g13165 ( 
.A1(n_11640),
.A2(n_1501),
.B1(n_1498),
.B2(n_1500),
.Y(n_13165)
);

INVx1_ASAP7_75t_L g13166 ( 
.A(n_12100),
.Y(n_13166)
);

AND2x2_ASAP7_75t_L g13167 ( 
.A(n_11755),
.B(n_1498),
.Y(n_13167)
);

INVx2_ASAP7_75t_L g13168 ( 
.A(n_11985),
.Y(n_13168)
);

AND2x2_ASAP7_75t_L g13169 ( 
.A(n_12269),
.B(n_1500),
.Y(n_13169)
);

NAND2xp5_ASAP7_75t_L g13170 ( 
.A(n_12412),
.B(n_1501),
.Y(n_13170)
);

NAND2xp5_ASAP7_75t_SL g13171 ( 
.A(n_11822),
.B(n_1502),
.Y(n_13171)
);

INVx1_ASAP7_75t_L g13172 ( 
.A(n_12110),
.Y(n_13172)
);

INVx2_ASAP7_75t_L g13173 ( 
.A(n_11768),
.Y(n_13173)
);

INVx2_ASAP7_75t_L g13174 ( 
.A(n_11907),
.Y(n_13174)
);

OR2x2_ASAP7_75t_L g13175 ( 
.A(n_12097),
.B(n_1502),
.Y(n_13175)
);

AND2x2_ASAP7_75t_L g13176 ( 
.A(n_11939),
.B(n_1503),
.Y(n_13176)
);

INVx1_ASAP7_75t_L g13177 ( 
.A(n_12204),
.Y(n_13177)
);

AOI22xp5_ASAP7_75t_L g13178 ( 
.A1(n_11645),
.A2(n_1505),
.B1(n_1503),
.B2(n_1504),
.Y(n_13178)
);

NAND2xp5_ASAP7_75t_SL g13179 ( 
.A(n_11805),
.B(n_1504),
.Y(n_13179)
);

AND2x2_ASAP7_75t_L g13180 ( 
.A(n_11970),
.B(n_1506),
.Y(n_13180)
);

INVx1_ASAP7_75t_L g13181 ( 
.A(n_12272),
.Y(n_13181)
);

NAND2xp5_ASAP7_75t_L g13182 ( 
.A(n_12416),
.B(n_1507),
.Y(n_13182)
);

NAND2xp33_ASAP7_75t_L g13183 ( 
.A(n_12444),
.B(n_1507),
.Y(n_13183)
);

NAND2xp5_ASAP7_75t_L g13184 ( 
.A(n_12425),
.B(n_1508),
.Y(n_13184)
);

AOI22xp5_ASAP7_75t_L g13185 ( 
.A1(n_11649),
.A2(n_1510),
.B1(n_1508),
.B2(n_1509),
.Y(n_13185)
);

INVx2_ASAP7_75t_L g13186 ( 
.A(n_12227),
.Y(n_13186)
);

INVx2_ASAP7_75t_L g13187 ( 
.A(n_12181),
.Y(n_13187)
);

CKINVDCx5p33_ASAP7_75t_R g13188 ( 
.A(n_11611),
.Y(n_13188)
);

NAND2xp5_ASAP7_75t_SL g13189 ( 
.A(n_12429),
.B(n_1509),
.Y(n_13189)
);

NAND2xp5_ASAP7_75t_L g13190 ( 
.A(n_12430),
.B(n_1511),
.Y(n_13190)
);

CKINVDCx5p33_ASAP7_75t_R g13191 ( 
.A(n_12308),
.Y(n_13191)
);

AOI22xp33_ASAP7_75t_L g13192 ( 
.A1(n_12249),
.A2(n_1514),
.B1(n_1512),
.B2(n_1513),
.Y(n_13192)
);

INVx4_ASAP7_75t_SL g13193 ( 
.A(n_11731),
.Y(n_13193)
);

OAI22xp5_ASAP7_75t_L g13194 ( 
.A1(n_12368),
.A2(n_1515),
.B1(n_1512),
.B2(n_1514),
.Y(n_13194)
);

NOR2xp33_ASAP7_75t_SL g13195 ( 
.A(n_11647),
.B(n_1516),
.Y(n_13195)
);

NAND2xp5_ASAP7_75t_L g13196 ( 
.A(n_12448),
.B(n_1517),
.Y(n_13196)
);

INVx1_ASAP7_75t_L g13197 ( 
.A(n_12103),
.Y(n_13197)
);

NAND2xp5_ASAP7_75t_L g13198 ( 
.A(n_12450),
.B(n_1517),
.Y(n_13198)
);

CKINVDCx20_ASAP7_75t_R g13199 ( 
.A(n_11685),
.Y(n_13199)
);

INVx2_ASAP7_75t_L g13200 ( 
.A(n_12280),
.Y(n_13200)
);

AND2x2_ASAP7_75t_L g13201 ( 
.A(n_11809),
.B(n_1518),
.Y(n_13201)
);

INVx2_ASAP7_75t_L g13202 ( 
.A(n_12291),
.Y(n_13202)
);

BUFx2_ASAP7_75t_L g13203 ( 
.A(n_12125),
.Y(n_13203)
);

NAND2xp5_ASAP7_75t_L g13204 ( 
.A(n_12463),
.B(n_1518),
.Y(n_13204)
);

INVxp67_ASAP7_75t_L g13205 ( 
.A(n_12478),
.Y(n_13205)
);

CKINVDCx5p33_ASAP7_75t_R g13206 ( 
.A(n_12339),
.Y(n_13206)
);

CKINVDCx5p33_ASAP7_75t_R g13207 ( 
.A(n_12343),
.Y(n_13207)
);

NAND2xp5_ASAP7_75t_SL g13208 ( 
.A(n_12482),
.B(n_1519),
.Y(n_13208)
);

AOI22xp5_ASAP7_75t_L g13209 ( 
.A1(n_11659),
.A2(n_1521),
.B1(n_1519),
.B2(n_1520),
.Y(n_13209)
);

AND2x2_ASAP7_75t_L g13210 ( 
.A(n_11812),
.B(n_1521),
.Y(n_13210)
);

INVxp33_ASAP7_75t_SL g13211 ( 
.A(n_12351),
.Y(n_13211)
);

AND2x2_ASAP7_75t_L g13212 ( 
.A(n_12264),
.B(n_1522),
.Y(n_13212)
);

AOI221xp5_ASAP7_75t_L g13213 ( 
.A1(n_12179),
.A2(n_1524),
.B1(n_1522),
.B2(n_1523),
.C(n_1525),
.Y(n_13213)
);

NAND2xp5_ASAP7_75t_L g13214 ( 
.A(n_12485),
.B(n_1523),
.Y(n_13214)
);

NOR2xp33_ASAP7_75t_L g13215 ( 
.A(n_12146),
.B(n_12221),
.Y(n_13215)
);

INVx1_ASAP7_75t_L g13216 ( 
.A(n_11790),
.Y(n_13216)
);

NAND2xp5_ASAP7_75t_SL g13217 ( 
.A(n_12486),
.B(n_1525),
.Y(n_13217)
);

AND2x2_ASAP7_75t_L g13218 ( 
.A(n_12067),
.B(n_1526),
.Y(n_13218)
);

NAND2xp5_ASAP7_75t_L g13219 ( 
.A(n_12487),
.B(n_1526),
.Y(n_13219)
);

INVx2_ASAP7_75t_L g13220 ( 
.A(n_12077),
.Y(n_13220)
);

NAND2xp5_ASAP7_75t_SL g13221 ( 
.A(n_12492),
.B(n_1527),
.Y(n_13221)
);

AND2x2_ASAP7_75t_L g13222 ( 
.A(n_12094),
.B(n_1527),
.Y(n_13222)
);

INVx1_ASAP7_75t_L g13223 ( 
.A(n_11792),
.Y(n_13223)
);

BUFx6f_ASAP7_75t_L g13224 ( 
.A(n_12143),
.Y(n_13224)
);

INVx2_ASAP7_75t_L g13225 ( 
.A(n_12320),
.Y(n_13225)
);

NAND2xp5_ASAP7_75t_SL g13226 ( 
.A(n_12494),
.B(n_1528),
.Y(n_13226)
);

AND3x1_ASAP7_75t_SL g13227 ( 
.A(n_12042),
.B(n_1528),
.C(n_1529),
.Y(n_13227)
);

NAND2xp5_ASAP7_75t_L g13228 ( 
.A(n_12503),
.B(n_1530),
.Y(n_13228)
);

AO22x1_ASAP7_75t_L g13229 ( 
.A1(n_12020),
.A2(n_1533),
.B1(n_1530),
.B2(n_1531),
.Y(n_13229)
);

NAND2xp5_ASAP7_75t_SL g13230 ( 
.A(n_12507),
.B(n_1533),
.Y(n_13230)
);

INVx1_ASAP7_75t_L g13231 ( 
.A(n_12382),
.Y(n_13231)
);

OAI22xp5_ASAP7_75t_L g13232 ( 
.A1(n_12473),
.A2(n_1536),
.B1(n_1534),
.B2(n_1535),
.Y(n_13232)
);

INVx2_ASAP7_75t_L g13233 ( 
.A(n_12469),
.Y(n_13233)
);

NAND2x1_ASAP7_75t_L g13234 ( 
.A(n_11683),
.B(n_11712),
.Y(n_13234)
);

AOI22xp33_ASAP7_75t_SL g13235 ( 
.A1(n_11664),
.A2(n_1536),
.B1(n_1534),
.B2(n_1535),
.Y(n_13235)
);

INVx2_ASAP7_75t_L g13236 ( 
.A(n_12199),
.Y(n_13236)
);

CKINVDCx5p33_ASAP7_75t_R g13237 ( 
.A(n_12385),
.Y(n_13237)
);

INVx2_ASAP7_75t_L g13238 ( 
.A(n_12201),
.Y(n_13238)
);

INVx1_ASAP7_75t_L g13239 ( 
.A(n_12510),
.Y(n_13239)
);

AOI22xp5_ASAP7_75t_L g13240 ( 
.A1(n_11810),
.A2(n_1539),
.B1(n_1537),
.B2(n_1538),
.Y(n_13240)
);

INVx1_ASAP7_75t_L g13241 ( 
.A(n_12512),
.Y(n_13241)
);

INVx1_ASAP7_75t_L g13242 ( 
.A(n_12515),
.Y(n_13242)
);

NAND2xp5_ASAP7_75t_SL g13243 ( 
.A(n_12285),
.B(n_1537),
.Y(n_13243)
);

INVx2_ASAP7_75t_L g13244 ( 
.A(n_12213),
.Y(n_13244)
);

BUFx4f_ASAP7_75t_SL g13245 ( 
.A(n_12226),
.Y(n_13245)
);

AND2x2_ASAP7_75t_L g13246 ( 
.A(n_11942),
.B(n_1538),
.Y(n_13246)
);

AND2x4_ASAP7_75t_L g13247 ( 
.A(n_12145),
.B(n_1539),
.Y(n_13247)
);

AND3x1_ASAP7_75t_SL g13248 ( 
.A(n_11863),
.B(n_1540),
.C(n_1541),
.Y(n_13248)
);

INVx1_ASAP7_75t_L g13249 ( 
.A(n_12284),
.Y(n_13249)
);

INVx1_ASAP7_75t_L g13250 ( 
.A(n_11706),
.Y(n_13250)
);

AND2x2_ASAP7_75t_L g13251 ( 
.A(n_12045),
.B(n_1541),
.Y(n_13251)
);

BUFx12f_ASAP7_75t_L g13252 ( 
.A(n_11620),
.Y(n_13252)
);

BUFx2_ASAP7_75t_L g13253 ( 
.A(n_12073),
.Y(n_13253)
);

INVx1_ASAP7_75t_L g13254 ( 
.A(n_12026),
.Y(n_13254)
);

INVx2_ASAP7_75t_L g13255 ( 
.A(n_12236),
.Y(n_13255)
);

AND2x2_ASAP7_75t_L g13256 ( 
.A(n_12087),
.B(n_1542),
.Y(n_13256)
);

INVx1_ASAP7_75t_L g13257 ( 
.A(n_12037),
.Y(n_13257)
);

OAI21xp5_ASAP7_75t_L g13258 ( 
.A1(n_11921),
.A2(n_1543),
.B(n_1544),
.Y(n_13258)
);

NAND2xp5_ASAP7_75t_L g13259 ( 
.A(n_12241),
.B(n_1543),
.Y(n_13259)
);

AND2x2_ASAP7_75t_L g13260 ( 
.A(n_12297),
.B(n_1544),
.Y(n_13260)
);

INVx1_ASAP7_75t_L g13261 ( 
.A(n_12034),
.Y(n_13261)
);

OAI21xp5_ASAP7_75t_L g13262 ( 
.A1(n_11925),
.A2(n_1545),
.B(n_1546),
.Y(n_13262)
);

INVxp67_ASAP7_75t_L g13263 ( 
.A(n_12275),
.Y(n_13263)
);

INVx2_ASAP7_75t_L g13264 ( 
.A(n_12299),
.Y(n_13264)
);

INVx2_ASAP7_75t_L g13265 ( 
.A(n_12304),
.Y(n_13265)
);

OAI22xp5_ASAP7_75t_SL g13266 ( 
.A1(n_12420),
.A2(n_1547),
.B1(n_1545),
.B2(n_1546),
.Y(n_13266)
);

AND2x2_ASAP7_75t_L g13267 ( 
.A(n_12007),
.B(n_1547),
.Y(n_13267)
);

AND2x2_ASAP7_75t_SL g13268 ( 
.A(n_11905),
.B(n_1548),
.Y(n_13268)
);

INVx2_ASAP7_75t_L g13269 ( 
.A(n_12068),
.Y(n_13269)
);

AND2x6_ASAP7_75t_L g13270 ( 
.A(n_11830),
.B(n_1548),
.Y(n_13270)
);

NAND2xp5_ASAP7_75t_L g13271 ( 
.A(n_11954),
.B(n_1549),
.Y(n_13271)
);

NAND2xp5_ASAP7_75t_L g13272 ( 
.A(n_11949),
.B(n_1549),
.Y(n_13272)
);

AND2x2_ASAP7_75t_L g13273 ( 
.A(n_11839),
.B(n_1550),
.Y(n_13273)
);

AND2x6_ASAP7_75t_L g13274 ( 
.A(n_12046),
.B(n_1550),
.Y(n_13274)
);

AND2x2_ASAP7_75t_L g13275 ( 
.A(n_11847),
.B(n_1551),
.Y(n_13275)
);

INVx2_ASAP7_75t_L g13276 ( 
.A(n_12044),
.Y(n_13276)
);

INVx1_ASAP7_75t_L g13277 ( 
.A(n_11864),
.Y(n_13277)
);

INVx1_ASAP7_75t_L g13278 ( 
.A(n_11798),
.Y(n_13278)
);

INVx1_ASAP7_75t_L g13279 ( 
.A(n_12333),
.Y(n_13279)
);

INVx2_ASAP7_75t_L g13280 ( 
.A(n_12435),
.Y(n_13280)
);

OR2x2_ASAP7_75t_L g13281 ( 
.A(n_11918),
.B(n_1551),
.Y(n_13281)
);

INVx1_ASAP7_75t_L g13282 ( 
.A(n_12367),
.Y(n_13282)
);

AOI22xp5_ASAP7_75t_L g13283 ( 
.A1(n_13195),
.A2(n_11697),
.B1(n_11815),
.B2(n_11631),
.Y(n_13283)
);

OAI21x1_ASAP7_75t_L g13284 ( 
.A1(n_12713),
.A2(n_11758),
.B(n_11926),
.Y(n_13284)
);

INVx2_ASAP7_75t_L g13285 ( 
.A(n_12695),
.Y(n_13285)
);

INVx1_ASAP7_75t_L g13286 ( 
.A(n_12661),
.Y(n_13286)
);

AOI21x1_ASAP7_75t_L g13287 ( 
.A1(n_12528),
.A2(n_12546),
.B(n_12783),
.Y(n_13287)
);

OAI21x1_ASAP7_75t_L g13288 ( 
.A1(n_13234),
.A2(n_11935),
.B(n_11932),
.Y(n_13288)
);

AOI21xp5_ASAP7_75t_L g13289 ( 
.A1(n_12953),
.A2(n_13243),
.B(n_13179),
.Y(n_13289)
);

INVx2_ASAP7_75t_SL g13290 ( 
.A(n_12564),
.Y(n_13290)
);

NAND2xp5_ASAP7_75t_L g13291 ( 
.A(n_13009),
.B(n_12029),
.Y(n_13291)
);

INVx3_ASAP7_75t_L g13292 ( 
.A(n_12804),
.Y(n_13292)
);

AO31x2_ASAP7_75t_L g13293 ( 
.A1(n_12691),
.A2(n_11860),
.A3(n_12461),
.B(n_12439),
.Y(n_13293)
);

NOR2xp33_ASAP7_75t_L g13294 ( 
.A(n_12752),
.B(n_13050),
.Y(n_13294)
);

NAND3xp33_ASAP7_75t_L g13295 ( 
.A(n_12559),
.B(n_11962),
.C(n_11959),
.Y(n_13295)
);

BUFx2_ASAP7_75t_L g13296 ( 
.A(n_12632),
.Y(n_13296)
);

CKINVDCx5p33_ASAP7_75t_R g13297 ( 
.A(n_12591),
.Y(n_13297)
);

OA21x2_ASAP7_75t_L g13298 ( 
.A1(n_12614),
.A2(n_11969),
.B(n_11967),
.Y(n_13298)
);

OAI21xp5_ASAP7_75t_L g13299 ( 
.A1(n_13143),
.A2(n_11979),
.B(n_11976),
.Y(n_13299)
);

AND2x2_ASAP7_75t_L g13300 ( 
.A(n_12525),
.B(n_12301),
.Y(n_13300)
);

AND2x2_ASAP7_75t_L g13301 ( 
.A(n_12541),
.B(n_12295),
.Y(n_13301)
);

HB1xp67_ASAP7_75t_L g13302 ( 
.A(n_12539),
.Y(n_13302)
);

AOI21xp5_ASAP7_75t_L g13303 ( 
.A1(n_13123),
.A2(n_11774),
.B(n_11763),
.Y(n_13303)
);

AOI221x1_ASAP7_75t_L g13304 ( 
.A1(n_12872),
.A2(n_11777),
.B1(n_12495),
.B2(n_12468),
.C(n_11700),
.Y(n_13304)
);

AO31x2_ASAP7_75t_L g13305 ( 
.A1(n_12942),
.A2(n_12182),
.A3(n_11991),
.B(n_11994),
.Y(n_13305)
);

AO31x2_ASAP7_75t_L g13306 ( 
.A1(n_12970),
.A2(n_12009),
.A3(n_12011),
.B(n_11982),
.Y(n_13306)
);

INVx1_ASAP7_75t_L g13307 ( 
.A(n_12563),
.Y(n_13307)
);

INVx3_ASAP7_75t_L g13308 ( 
.A(n_12852),
.Y(n_13308)
);

NAND2xp5_ASAP7_75t_L g13309 ( 
.A(n_13202),
.B(n_12016),
.Y(n_13309)
);

NAND2xp5_ASAP7_75t_L g13310 ( 
.A(n_12582),
.B(n_12018),
.Y(n_13310)
);

AO31x2_ASAP7_75t_L g13311 ( 
.A1(n_12998),
.A2(n_12032),
.A3(n_12035),
.B(n_12031),
.Y(n_13311)
);

INVx1_ASAP7_75t_L g13312 ( 
.A(n_12568),
.Y(n_13312)
);

AOI21xp5_ASAP7_75t_L g13313 ( 
.A1(n_12865),
.A2(n_13183),
.B(n_12773),
.Y(n_13313)
);

OAI21x1_ASAP7_75t_L g13314 ( 
.A1(n_13034),
.A2(n_12060),
.B(n_12054),
.Y(n_13314)
);

OAI21x1_ASAP7_75t_L g13315 ( 
.A1(n_13200),
.A2(n_12069),
.B(n_12066),
.Y(n_13315)
);

OAI21xp5_ASAP7_75t_SL g13316 ( 
.A1(n_12917),
.A2(n_11816),
.B(n_12305),
.Y(n_13316)
);

OR2x2_ASAP7_75t_L g13317 ( 
.A(n_12548),
.B(n_12071),
.Y(n_13317)
);

NAND3xp33_ASAP7_75t_SL g13318 ( 
.A(n_13138),
.B(n_12364),
.C(n_12315),
.Y(n_13318)
);

O2A1O1Ixp33_ASAP7_75t_L g13319 ( 
.A1(n_12842),
.A2(n_11618),
.B(n_11922),
.C(n_12437),
.Y(n_13319)
);

OAI21xp5_ASAP7_75t_L g13320 ( 
.A1(n_13166),
.A2(n_12083),
.B(n_12078),
.Y(n_13320)
);

O2A1O1Ixp33_ASAP7_75t_SL g13321 ( 
.A1(n_12979),
.A2(n_11804),
.B(n_12406),
.C(n_12386),
.Y(n_13321)
);

BUFx6f_ASAP7_75t_L g13322 ( 
.A(n_12543),
.Y(n_13322)
);

AO31x2_ASAP7_75t_L g13323 ( 
.A1(n_12946),
.A2(n_12111),
.A3(n_12114),
.B(n_12086),
.Y(n_13323)
);

OAI21x1_ASAP7_75t_L g13324 ( 
.A1(n_13060),
.A2(n_12123),
.B(n_12116),
.Y(n_13324)
);

BUFx5_ASAP7_75t_L g13325 ( 
.A(n_13069),
.Y(n_13325)
);

OAI21x1_ASAP7_75t_L g13326 ( 
.A1(n_13093),
.A2(n_12162),
.B(n_12131),
.Y(n_13326)
);

AND2x4_ASAP7_75t_L g13327 ( 
.A(n_12853),
.B(n_11852),
.Y(n_13327)
);

AOI21xp5_ASAP7_75t_L g13328 ( 
.A1(n_12914),
.A2(n_11604),
.B(n_11715),
.Y(n_13328)
);

INVxp67_ASAP7_75t_L g13329 ( 
.A(n_12747),
.Y(n_13329)
);

OAI21x1_ASAP7_75t_L g13330 ( 
.A1(n_12987),
.A2(n_12166),
.B(n_11795),
.Y(n_13330)
);

OAI21x1_ASAP7_75t_L g13331 ( 
.A1(n_13005),
.A2(n_12193),
.B(n_12185),
.Y(n_13331)
);

INVx1_ASAP7_75t_L g13332 ( 
.A(n_12577),
.Y(n_13332)
);

AND2x4_ASAP7_75t_L g13333 ( 
.A(n_12571),
.B(n_11853),
.Y(n_13333)
);

AO21x2_ASAP7_75t_L g13334 ( 
.A1(n_13036),
.A2(n_12214),
.B(n_12211),
.Y(n_13334)
);

A2O1A1Ixp33_ASAP7_75t_L g13335 ( 
.A1(n_12547),
.A2(n_12457),
.B(n_12513),
.C(n_12449),
.Y(n_13335)
);

NOR2xp33_ASAP7_75t_L g13336 ( 
.A(n_13079),
.B(n_12136),
.Y(n_13336)
);

BUFx2_ASAP7_75t_SL g13337 ( 
.A(n_12810),
.Y(n_13337)
);

OAI21x1_ASAP7_75t_L g13338 ( 
.A1(n_12989),
.A2(n_12223),
.B(n_12217),
.Y(n_13338)
);

OAI22xp33_ASAP7_75t_L g13339 ( 
.A1(n_13158),
.A2(n_13253),
.B1(n_12999),
.B2(n_13165),
.Y(n_13339)
);

INVx2_ASAP7_75t_L g13340 ( 
.A(n_12696),
.Y(n_13340)
);

OAI21x1_ASAP7_75t_L g13341 ( 
.A1(n_13012),
.A2(n_12234),
.B(n_12233),
.Y(n_13341)
);

INVx1_ASAP7_75t_L g13342 ( 
.A(n_12583),
.Y(n_13342)
);

NAND2x1_ASAP7_75t_L g13343 ( 
.A(n_12794),
.B(n_11610),
.Y(n_13343)
);

HB1xp67_ASAP7_75t_L g13344 ( 
.A(n_12558),
.Y(n_13344)
);

AND2x2_ASAP7_75t_L g13345 ( 
.A(n_12600),
.B(n_11856),
.Y(n_13345)
);

AOI22xp5_ASAP7_75t_L g13346 ( 
.A1(n_12617),
.A2(n_11885),
.B1(n_11895),
.B2(n_11675),
.Y(n_13346)
);

AOI21xp5_ASAP7_75t_L g13347 ( 
.A1(n_12816),
.A2(n_12257),
.B(n_12254),
.Y(n_13347)
);

NAND2xp5_ASAP7_75t_L g13348 ( 
.A(n_12567),
.B(n_11726),
.Y(n_13348)
);

AND2x2_ASAP7_75t_L g13349 ( 
.A(n_12580),
.B(n_11857),
.Y(n_13349)
);

HB1xp67_ASAP7_75t_L g13350 ( 
.A(n_12606),
.Y(n_13350)
);

NAND2xp5_ASAP7_75t_L g13351 ( 
.A(n_12684),
.B(n_11739),
.Y(n_13351)
);

INVx3_ASAP7_75t_L g13352 ( 
.A(n_12724),
.Y(n_13352)
);

INVx2_ASAP7_75t_L g13353 ( 
.A(n_12702),
.Y(n_13353)
);

INVx1_ASAP7_75t_L g13354 ( 
.A(n_12592),
.Y(n_13354)
);

INVx1_ASAP7_75t_L g13355 ( 
.A(n_12597),
.Y(n_13355)
);

AOI21xp5_ASAP7_75t_L g13356 ( 
.A1(n_12693),
.A2(n_12262),
.B(n_12261),
.Y(n_13356)
);

CKINVDCx5p33_ASAP7_75t_R g13357 ( 
.A(n_12542),
.Y(n_13357)
);

INVx1_ASAP7_75t_L g13358 ( 
.A(n_12605),
.Y(n_13358)
);

A2O1A1Ixp33_ASAP7_75t_L g13359 ( 
.A1(n_12834),
.A2(n_11928),
.B(n_11927),
.C(n_12057),
.Y(n_13359)
);

BUFx6f_ASAP7_75t_L g13360 ( 
.A(n_12543),
.Y(n_13360)
);

INVx2_ASAP7_75t_L g13361 ( 
.A(n_12647),
.Y(n_13361)
);

AOI21xp5_ASAP7_75t_L g13362 ( 
.A1(n_12779),
.A2(n_12283),
.B(n_12274),
.Y(n_13362)
);

OAI22xp5_ASAP7_75t_L g13363 ( 
.A1(n_13192),
.A2(n_11873),
.B1(n_11974),
.B2(n_12099),
.Y(n_13363)
);

INVx2_ASAP7_75t_SL g13364 ( 
.A(n_12722),
.Y(n_13364)
);

O2A1O1Ixp33_ASAP7_75t_L g13365 ( 
.A1(n_12522),
.A2(n_11641),
.B(n_11874),
.C(n_12246),
.Y(n_13365)
);

INVx1_ASAP7_75t_L g13366 ( 
.A(n_12608),
.Y(n_13366)
);

BUFx2_ASAP7_75t_L g13367 ( 
.A(n_12652),
.Y(n_13367)
);

OAI21xp5_ASAP7_75t_L g13368 ( 
.A1(n_13205),
.A2(n_11717),
.B(n_11865),
.Y(n_13368)
);

INVx1_ASAP7_75t_L g13369 ( 
.A(n_12613),
.Y(n_13369)
);

OAI21x1_ASAP7_75t_L g13370 ( 
.A1(n_13013),
.A2(n_11684),
.B(n_11617),
.Y(n_13370)
);

AOI31xp67_ASAP7_75t_L g13371 ( 
.A1(n_13055),
.A2(n_11814),
.A3(n_11868),
.B(n_11866),
.Y(n_13371)
);

AOI21xp5_ASAP7_75t_L g13372 ( 
.A1(n_13002),
.A2(n_11886),
.B(n_11871),
.Y(n_13372)
);

INVx2_ASAP7_75t_SL g13373 ( 
.A(n_12722),
.Y(n_13373)
);

OA21x2_ASAP7_75t_L g13374 ( 
.A1(n_13109),
.A2(n_11893),
.B(n_11888),
.Y(n_13374)
);

O2A1O1Ixp33_ASAP7_75t_L g13375 ( 
.A1(n_13046),
.A2(n_11779),
.B(n_11910),
.C(n_1554),
.Y(n_13375)
);

NAND2xp5_ASAP7_75t_SL g13376 ( 
.A(n_13126),
.B(n_1552),
.Y(n_13376)
);

AOI21xp5_ASAP7_75t_L g13377 ( 
.A1(n_13121),
.A2(n_1552),
.B(n_1553),
.Y(n_13377)
);

INVx2_ASAP7_75t_L g13378 ( 
.A(n_12649),
.Y(n_13378)
);

AO32x2_ASAP7_75t_L g13379 ( 
.A1(n_12960),
.A2(n_1557),
.A3(n_1555),
.B1(n_1556),
.B2(n_1558),
.Y(n_13379)
);

NAND2x1p5_ASAP7_75t_L g13380 ( 
.A(n_12610),
.B(n_1555),
.Y(n_13380)
);

BUFx6f_ASAP7_75t_L g13381 ( 
.A(n_12552),
.Y(n_13381)
);

OAI21x1_ASAP7_75t_L g13382 ( 
.A1(n_13048),
.A2(n_1556),
.B(n_1557),
.Y(n_13382)
);

NAND2xp5_ASAP7_75t_L g13383 ( 
.A(n_13122),
.B(n_13129),
.Y(n_13383)
);

AOI21xp5_ASAP7_75t_L g13384 ( 
.A1(n_13189),
.A2(n_1558),
.B(n_1559),
.Y(n_13384)
);

OAI21x1_ASAP7_75t_L g13385 ( 
.A1(n_13038),
.A2(n_1559),
.B(n_1560),
.Y(n_13385)
);

NAND2xp5_ASAP7_75t_SL g13386 ( 
.A(n_13151),
.B(n_1560),
.Y(n_13386)
);

AOI221xp5_ASAP7_75t_L g13387 ( 
.A1(n_12579),
.A2(n_1563),
.B1(n_1561),
.B2(n_1562),
.C(n_1564),
.Y(n_13387)
);

INVx2_ASAP7_75t_L g13388 ( 
.A(n_12653),
.Y(n_13388)
);

OAI21x1_ASAP7_75t_L g13389 ( 
.A1(n_13056),
.A2(n_12933),
.B(n_13127),
.Y(n_13389)
);

AOI21xp5_ASAP7_75t_L g13390 ( 
.A1(n_13208),
.A2(n_1561),
.B(n_1562),
.Y(n_13390)
);

AOI21xp5_ASAP7_75t_L g13391 ( 
.A1(n_13217),
.A2(n_1564),
.B(n_1565),
.Y(n_13391)
);

AO31x2_ASAP7_75t_L g13392 ( 
.A1(n_13155),
.A2(n_1567),
.A3(n_1565),
.B(n_1566),
.Y(n_13392)
);

AND2x2_ASAP7_75t_L g13393 ( 
.A(n_12663),
.B(n_1566),
.Y(n_13393)
);

INVx2_ASAP7_75t_L g13394 ( 
.A(n_12662),
.Y(n_13394)
);

INVx2_ASAP7_75t_L g13395 ( 
.A(n_12667),
.Y(n_13395)
);

A2O1A1Ixp33_ASAP7_75t_L g13396 ( 
.A1(n_12768),
.A2(n_1569),
.B(n_1567),
.C(n_1568),
.Y(n_13396)
);

OAI21x1_ASAP7_75t_L g13397 ( 
.A1(n_13043),
.A2(n_1570),
.B(n_1571),
.Y(n_13397)
);

OAI21x1_ASAP7_75t_L g13398 ( 
.A1(n_13095),
.A2(n_1570),
.B(n_1571),
.Y(n_13398)
);

INVx2_ASAP7_75t_L g13399 ( 
.A(n_12629),
.Y(n_13399)
);

INVx2_ASAP7_75t_L g13400 ( 
.A(n_12630),
.Y(n_13400)
);

INVx3_ASAP7_75t_L g13401 ( 
.A(n_12682),
.Y(n_13401)
);

BUFx12f_ASAP7_75t_L g13402 ( 
.A(n_12544),
.Y(n_13402)
);

NAND2xp5_ASAP7_75t_SL g13403 ( 
.A(n_13151),
.B(n_1572),
.Y(n_13403)
);

INVx1_ASAP7_75t_L g13404 ( 
.A(n_12636),
.Y(n_13404)
);

AOI21xp5_ASAP7_75t_L g13405 ( 
.A1(n_13221),
.A2(n_1572),
.B(n_1573),
.Y(n_13405)
);

NAND2xp5_ASAP7_75t_L g13406 ( 
.A(n_12748),
.B(n_1573),
.Y(n_13406)
);

AOI22xp5_ASAP7_75t_L g13407 ( 
.A1(n_13136),
.A2(n_1576),
.B1(n_1574),
.B2(n_1575),
.Y(n_13407)
);

NOR2xp33_ASAP7_75t_L g13408 ( 
.A(n_12745),
.B(n_1574),
.Y(n_13408)
);

AO31x2_ASAP7_75t_L g13409 ( 
.A1(n_13077),
.A2(n_1578),
.A3(n_1576),
.B(n_1577),
.Y(n_13409)
);

OAI21x1_ASAP7_75t_L g13410 ( 
.A1(n_13161),
.A2(n_1579),
.B(n_1580),
.Y(n_13410)
);

A2O1A1Ixp33_ASAP7_75t_L g13411 ( 
.A1(n_12958),
.A2(n_1581),
.B(n_1579),
.C(n_1580),
.Y(n_13411)
);

BUFx3_ASAP7_75t_L g13412 ( 
.A(n_12698),
.Y(n_13412)
);

AOI21xp5_ASAP7_75t_L g13413 ( 
.A1(n_13226),
.A2(n_1582),
.B(n_1583),
.Y(n_13413)
);

AOI21xp5_ASAP7_75t_L g13414 ( 
.A1(n_13230),
.A2(n_1582),
.B(n_1583),
.Y(n_13414)
);

AOI21x1_ASAP7_75t_L g13415 ( 
.A1(n_12602),
.A2(n_1584),
.B(n_1585),
.Y(n_13415)
);

A2O1A1Ixp33_ASAP7_75t_L g13416 ( 
.A1(n_13215),
.A2(n_1586),
.B(n_1584),
.C(n_1585),
.Y(n_13416)
);

NAND2xp5_ASAP7_75t_SL g13417 ( 
.A(n_13224),
.B(n_13119),
.Y(n_13417)
);

OAI21x1_ASAP7_75t_L g13418 ( 
.A1(n_12808),
.A2(n_1586),
.B(n_1587),
.Y(n_13418)
);

O2A1O1Ixp33_ASAP7_75t_L g13419 ( 
.A1(n_12908),
.A2(n_1589),
.B(n_1587),
.C(n_1588),
.Y(n_13419)
);

NAND2xp5_ASAP7_75t_L g13420 ( 
.A(n_12890),
.B(n_1588),
.Y(n_13420)
);

OAI22xp5_ASAP7_75t_L g13421 ( 
.A1(n_13033),
.A2(n_1591),
.B1(n_1589),
.B2(n_1590),
.Y(n_13421)
);

AOI21xp5_ASAP7_75t_L g13422 ( 
.A1(n_12985),
.A2(n_1590),
.B(n_1592),
.Y(n_13422)
);

HB1xp67_ASAP7_75t_SL g13423 ( 
.A(n_12737),
.Y(n_13423)
);

AOI22xp5_ASAP7_75t_L g13424 ( 
.A1(n_13252),
.A2(n_1594),
.B1(n_1592),
.B2(n_1593),
.Y(n_13424)
);

NAND2xp5_ASAP7_75t_L g13425 ( 
.A(n_13113),
.B(n_1593),
.Y(n_13425)
);

A2O1A1Ixp33_ASAP7_75t_L g13426 ( 
.A1(n_13027),
.A2(n_12520),
.B(n_12685),
.C(n_12609),
.Y(n_13426)
);

NAND2xp5_ASAP7_75t_L g13427 ( 
.A(n_12694),
.B(n_1594),
.Y(n_13427)
);

NAND2xp5_ASAP7_75t_L g13428 ( 
.A(n_12714),
.B(n_1595),
.Y(n_13428)
);

OAI221xp5_ASAP7_75t_L g13429 ( 
.A1(n_12699),
.A2(n_1597),
.B1(n_1595),
.B2(n_1596),
.C(n_1598),
.Y(n_13429)
);

INVx1_ASAP7_75t_L g13430 ( 
.A(n_12641),
.Y(n_13430)
);

OAI21x1_ASAP7_75t_L g13431 ( 
.A1(n_13216),
.A2(n_1596),
.B(n_1597),
.Y(n_13431)
);

OAI21x1_ASAP7_75t_L g13432 ( 
.A1(n_13223),
.A2(n_1598),
.B(n_1599),
.Y(n_13432)
);

NAND2xp5_ASAP7_75t_L g13433 ( 
.A(n_12717),
.B(n_1599),
.Y(n_13433)
);

BUFx2_ASAP7_75t_L g13434 ( 
.A(n_13063),
.Y(n_13434)
);

NAND2xp5_ASAP7_75t_L g13435 ( 
.A(n_12725),
.B(n_1600),
.Y(n_13435)
);

BUFx3_ASAP7_75t_L g13436 ( 
.A(n_12537),
.Y(n_13436)
);

BUFx12f_ASAP7_75t_L g13437 ( 
.A(n_12657),
.Y(n_13437)
);

NAND2xp5_ASAP7_75t_L g13438 ( 
.A(n_12744),
.B(n_1600),
.Y(n_13438)
);

OAI21xp5_ASAP7_75t_L g13439 ( 
.A1(n_12883),
.A2(n_1601),
.B(n_1602),
.Y(n_13439)
);

OR2x6_ASAP7_75t_L g13440 ( 
.A(n_12710),
.B(n_1602),
.Y(n_13440)
);

OAI22xp5_ASAP7_75t_L g13441 ( 
.A1(n_13090),
.A2(n_1605),
.B1(n_1603),
.B2(n_1604),
.Y(n_13441)
);

AOI21xp5_ASAP7_75t_L g13442 ( 
.A1(n_13258),
.A2(n_1603),
.B(n_1604),
.Y(n_13442)
);

OAI21xp5_ASAP7_75t_L g13443 ( 
.A1(n_12800),
.A2(n_1606),
.B(n_1607),
.Y(n_13443)
);

NAND2xp5_ASAP7_75t_L g13444 ( 
.A(n_12762),
.B(n_1606),
.Y(n_13444)
);

INVx1_ASAP7_75t_L g13445 ( 
.A(n_12646),
.Y(n_13445)
);

INVx2_ASAP7_75t_SL g13446 ( 
.A(n_12710),
.Y(n_13446)
);

NAND2xp5_ASAP7_75t_L g13447 ( 
.A(n_12774),
.B(n_1608),
.Y(n_13447)
);

INVx1_ASAP7_75t_L g13448 ( 
.A(n_12654),
.Y(n_13448)
);

INVx2_ASAP7_75t_SL g13449 ( 
.A(n_12616),
.Y(n_13449)
);

AOI21xp5_ASAP7_75t_L g13450 ( 
.A1(n_13262),
.A2(n_1609),
.B(n_1610),
.Y(n_13450)
);

AOI211x1_ASAP7_75t_L g13451 ( 
.A1(n_12672),
.A2(n_13010),
.B(n_12851),
.C(n_13229),
.Y(n_13451)
);

AOI221x1_ASAP7_75t_L g13452 ( 
.A1(n_12706),
.A2(n_1612),
.B1(n_1609),
.B2(n_1611),
.C(n_1613),
.Y(n_13452)
);

A2O1A1Ixp33_ASAP7_75t_L g13453 ( 
.A1(n_12711),
.A2(n_1613),
.B(n_1611),
.C(n_1612),
.Y(n_13453)
);

AOI221x1_ASAP7_75t_L g13454 ( 
.A1(n_12731),
.A2(n_1616),
.B1(n_1614),
.B2(n_1615),
.C(n_1617),
.Y(n_13454)
);

AOI21xp5_ASAP7_75t_L g13455 ( 
.A1(n_12566),
.A2(n_1614),
.B(n_1615),
.Y(n_13455)
);

INVx1_ASAP7_75t_L g13456 ( 
.A(n_12659),
.Y(n_13456)
);

CKINVDCx5p33_ASAP7_75t_R g13457 ( 
.A(n_12523),
.Y(n_13457)
);

INVx2_ASAP7_75t_L g13458 ( 
.A(n_12668),
.Y(n_13458)
);

NOR2xp33_ASAP7_75t_L g13459 ( 
.A(n_13035),
.B(n_1616),
.Y(n_13459)
);

INVx1_ASAP7_75t_L g13460 ( 
.A(n_12669),
.Y(n_13460)
);

INVx2_ASAP7_75t_L g13461 ( 
.A(n_12660),
.Y(n_13461)
);

OAI21x1_ASAP7_75t_L g13462 ( 
.A1(n_13059),
.A2(n_1617),
.B(n_1618),
.Y(n_13462)
);

AO31x2_ASAP7_75t_L g13463 ( 
.A1(n_13083),
.A2(n_1620),
.A3(n_1618),
.B(n_1619),
.Y(n_13463)
);

OAI22xp5_ASAP7_75t_L g13464 ( 
.A1(n_13128),
.A2(n_1621),
.B1(n_1619),
.B2(n_1620),
.Y(n_13464)
);

OAI22xp33_ASAP7_75t_L g13465 ( 
.A1(n_13146),
.A2(n_1623),
.B1(n_1621),
.B2(n_1622),
.Y(n_13465)
);

BUFx10_ASAP7_75t_L g13466 ( 
.A(n_12574),
.Y(n_13466)
);

NAND2xp5_ASAP7_75t_L g13467 ( 
.A(n_12788),
.B(n_1622),
.Y(n_13467)
);

INVx1_ASAP7_75t_L g13468 ( 
.A(n_12527),
.Y(n_13468)
);

AND2x4_ASAP7_75t_L g13469 ( 
.A(n_13125),
.B(n_1623),
.Y(n_13469)
);

AND2x4_ASAP7_75t_L g13470 ( 
.A(n_12812),
.B(n_1624),
.Y(n_13470)
);

NAND2xp5_ASAP7_75t_L g13471 ( 
.A(n_12707),
.B(n_1624),
.Y(n_13471)
);

AND2x2_ASAP7_75t_L g13472 ( 
.A(n_12697),
.B(n_1625),
.Y(n_13472)
);

NAND3xp33_ASAP7_75t_L g13473 ( 
.A(n_13249),
.B(n_1625),
.C(n_1626),
.Y(n_13473)
);

INVx1_ASAP7_75t_L g13474 ( 
.A(n_12540),
.Y(n_13474)
);

INVx2_ASAP7_75t_SL g13475 ( 
.A(n_12755),
.Y(n_13475)
);

NOR2xp33_ASAP7_75t_L g13476 ( 
.A(n_13015),
.B(n_1627),
.Y(n_13476)
);

INVx1_ASAP7_75t_L g13477 ( 
.A(n_12557),
.Y(n_13477)
);

BUFx6f_ASAP7_75t_L g13478 ( 
.A(n_12552),
.Y(n_13478)
);

O2A1O1Ixp5_ASAP7_75t_SL g13479 ( 
.A1(n_13047),
.A2(n_1629),
.B(n_1627),
.C(n_1628),
.Y(n_13479)
);

AO31x2_ASAP7_75t_L g13480 ( 
.A1(n_13084),
.A2(n_1631),
.A3(n_1628),
.B(n_1629),
.Y(n_13480)
);

OAI21xp5_ASAP7_75t_L g13481 ( 
.A1(n_13178),
.A2(n_1632),
.B(n_1633),
.Y(n_13481)
);

OA21x2_ASAP7_75t_L g13482 ( 
.A1(n_13085),
.A2(n_1632),
.B(n_1633),
.Y(n_13482)
);

OAI21xp5_ASAP7_75t_L g13483 ( 
.A1(n_13185),
.A2(n_1635),
.B(n_1636),
.Y(n_13483)
);

AND2x4_ASAP7_75t_L g13484 ( 
.A(n_12819),
.B(n_1636),
.Y(n_13484)
);

A2O1A1Ixp33_ASAP7_75t_L g13485 ( 
.A1(n_12835),
.A2(n_1639),
.B(n_1637),
.C(n_1638),
.Y(n_13485)
);

NAND2xp5_ASAP7_75t_SL g13486 ( 
.A(n_13224),
.B(n_1638),
.Y(n_13486)
);

INVx2_ASAP7_75t_SL g13487 ( 
.A(n_12651),
.Y(n_13487)
);

OAI21x1_ASAP7_75t_L g13488 ( 
.A1(n_13066),
.A2(n_13160),
.B(n_13239),
.Y(n_13488)
);

AOI21xp5_ASAP7_75t_L g13489 ( 
.A1(n_12754),
.A2(n_1640),
.B(n_1641),
.Y(n_13489)
);

AOI22xp5_ASAP7_75t_L g13490 ( 
.A1(n_12976),
.A2(n_13274),
.B1(n_13270),
.B2(n_12971),
.Y(n_13490)
);

NAND2xp5_ASAP7_75t_L g13491 ( 
.A(n_12715),
.B(n_1640),
.Y(n_13491)
);

NOR2xp33_ASAP7_75t_L g13492 ( 
.A(n_13120),
.B(n_1641),
.Y(n_13492)
);

OAI21x1_ASAP7_75t_L g13493 ( 
.A1(n_13241),
.A2(n_1642),
.B(n_1643),
.Y(n_13493)
);

INVx1_ASAP7_75t_L g13494 ( 
.A(n_12561),
.Y(n_13494)
);

BUFx10_ASAP7_75t_L g13495 ( 
.A(n_12735),
.Y(n_13495)
);

AND2x2_ASAP7_75t_SL g13496 ( 
.A(n_12727),
.B(n_1642),
.Y(n_13496)
);

AOI21xp5_ASAP7_75t_L g13497 ( 
.A1(n_13070),
.A2(n_1643),
.B(n_1644),
.Y(n_13497)
);

OAI21x1_ASAP7_75t_L g13498 ( 
.A1(n_13242),
.A2(n_1644),
.B(n_1645),
.Y(n_13498)
);

INVx1_ASAP7_75t_L g13499 ( 
.A(n_12581),
.Y(n_13499)
);

AOI22xp33_ASAP7_75t_L g13500 ( 
.A1(n_13274),
.A2(n_1647),
.B1(n_1645),
.B2(n_1646),
.Y(n_13500)
);

O2A1O1Ixp33_ASAP7_75t_SL g13501 ( 
.A1(n_12907),
.A2(n_1649),
.B(n_1647),
.C(n_1648),
.Y(n_13501)
);

A2O1A1Ixp33_ASAP7_75t_L g13502 ( 
.A1(n_13133),
.A2(n_1650),
.B(n_1648),
.C(n_1649),
.Y(n_13502)
);

BUFx3_ASAP7_75t_L g13503 ( 
.A(n_12633),
.Y(n_13503)
);

INVxp67_ASAP7_75t_SL g13504 ( 
.A(n_12947),
.Y(n_13504)
);

O2A1O1Ixp5_ASAP7_75t_L g13505 ( 
.A1(n_12887),
.A2(n_1652),
.B(n_1650),
.C(n_1651),
.Y(n_13505)
);

INVxp67_ASAP7_75t_SL g13506 ( 
.A(n_12681),
.Y(n_13506)
);

INVx2_ASAP7_75t_L g13507 ( 
.A(n_12703),
.Y(n_13507)
);

NOR2xp33_ASAP7_75t_L g13508 ( 
.A(n_13032),
.B(n_1651),
.Y(n_13508)
);

AO31x2_ASAP7_75t_L g13509 ( 
.A1(n_13147),
.A2(n_1654),
.A3(n_1652),
.B(n_1653),
.Y(n_13509)
);

CKINVDCx5p33_ASAP7_75t_R g13510 ( 
.A(n_12680),
.Y(n_13510)
);

BUFx3_ASAP7_75t_L g13511 ( 
.A(n_12676),
.Y(n_13511)
);

AND2x2_ASAP7_75t_L g13512 ( 
.A(n_12700),
.B(n_1653),
.Y(n_13512)
);

OAI21x1_ASAP7_75t_L g13513 ( 
.A1(n_13116),
.A2(n_1654),
.B(n_1655),
.Y(n_13513)
);

OAI21x1_ASAP7_75t_L g13514 ( 
.A1(n_13152),
.A2(n_1656),
.B(n_1657),
.Y(n_13514)
);

A2O1A1Ixp33_ASAP7_75t_L g13515 ( 
.A1(n_13001),
.A2(n_1658),
.B(n_1656),
.C(n_1657),
.Y(n_13515)
);

AOI21xp5_ASAP7_75t_L g13516 ( 
.A1(n_13111),
.A2(n_1659),
.B(n_1660),
.Y(n_13516)
);

AOI21xp5_ASAP7_75t_L g13517 ( 
.A1(n_12930),
.A2(n_1659),
.B(n_1660),
.Y(n_13517)
);

BUFx12f_ASAP7_75t_L g13518 ( 
.A(n_12671),
.Y(n_13518)
);

INVx1_ASAP7_75t_L g13519 ( 
.A(n_12590),
.Y(n_13519)
);

INVx1_ASAP7_75t_SL g13520 ( 
.A(n_12746),
.Y(n_13520)
);

AOI21xp5_ASAP7_75t_L g13521 ( 
.A1(n_13171),
.A2(n_1661),
.B(n_1662),
.Y(n_13521)
);

HB1xp67_ASAP7_75t_L g13522 ( 
.A(n_12705),
.Y(n_13522)
);

OAI21x1_ASAP7_75t_L g13523 ( 
.A1(n_12975),
.A2(n_1661),
.B(n_1662),
.Y(n_13523)
);

O2A1O1Ixp33_ASAP7_75t_L g13524 ( 
.A1(n_13135),
.A2(n_1665),
.B(n_1663),
.C(n_1664),
.Y(n_13524)
);

OR2x2_ASAP7_75t_L g13525 ( 
.A(n_12594),
.B(n_1663),
.Y(n_13525)
);

BUFx4f_ASAP7_75t_L g13526 ( 
.A(n_12818),
.Y(n_13526)
);

OAI22xp5_ASAP7_75t_L g13527 ( 
.A1(n_13157),
.A2(n_1666),
.B1(n_1664),
.B2(n_1665),
.Y(n_13527)
);

AOI21xp5_ASAP7_75t_L g13528 ( 
.A1(n_12826),
.A2(n_12940),
.B(n_12806),
.Y(n_13528)
);

NAND2xp5_ASAP7_75t_L g13529 ( 
.A(n_12723),
.B(n_1666),
.Y(n_13529)
);

NOR2xp33_ASAP7_75t_L g13530 ( 
.A(n_12997),
.B(n_1667),
.Y(n_13530)
);

CKINVDCx20_ASAP7_75t_R g13531 ( 
.A(n_12576),
.Y(n_13531)
);

OAI21x1_ASAP7_75t_L g13532 ( 
.A1(n_13231),
.A2(n_1667),
.B(n_1668),
.Y(n_13532)
);

INVxp67_ASAP7_75t_SL g13533 ( 
.A(n_12655),
.Y(n_13533)
);

AOI21xp5_ASAP7_75t_L g13534 ( 
.A1(n_13088),
.A2(n_1668),
.B(n_1669),
.Y(n_13534)
);

NOR2xp33_ASAP7_75t_L g13535 ( 
.A(n_12782),
.B(n_1669),
.Y(n_13535)
);

OAI22x1_ASAP7_75t_L g13536 ( 
.A1(n_13104),
.A2(n_1672),
.B1(n_1670),
.B2(n_1671),
.Y(n_13536)
);

INVx2_ASAP7_75t_L g13537 ( 
.A(n_12595),
.Y(n_13537)
);

INVx1_ASAP7_75t_SL g13538 ( 
.A(n_12570),
.Y(n_13538)
);

NOR2xp33_ASAP7_75t_L g13539 ( 
.A(n_12766),
.B(n_1670),
.Y(n_13539)
);

AO31x2_ASAP7_75t_L g13540 ( 
.A1(n_13150),
.A2(n_1674),
.A3(n_1671),
.B(n_1673),
.Y(n_13540)
);

AND2x2_ASAP7_75t_L g13541 ( 
.A(n_12797),
.B(n_1673),
.Y(n_13541)
);

AOI21xp5_ASAP7_75t_L g13542 ( 
.A1(n_13053),
.A2(n_13106),
.B(n_13139),
.Y(n_13542)
);

INVx1_ASAP7_75t_L g13543 ( 
.A(n_12604),
.Y(n_13543)
);

INVx3_ASAP7_75t_L g13544 ( 
.A(n_12793),
.Y(n_13544)
);

OAI21x1_ASAP7_75t_L g13545 ( 
.A1(n_13225),
.A2(n_1674),
.B(n_1675),
.Y(n_13545)
);

OAI22xp5_ASAP7_75t_L g13546 ( 
.A1(n_12678),
.A2(n_1677),
.B1(n_1675),
.B2(n_1676),
.Y(n_13546)
);

OAI21x1_ASAP7_75t_L g13547 ( 
.A1(n_13233),
.A2(n_1676),
.B(n_1677),
.Y(n_13547)
);

NAND2xp5_ASAP7_75t_L g13548 ( 
.A(n_12758),
.B(n_1678),
.Y(n_13548)
);

OR2x6_ASAP7_75t_L g13549 ( 
.A(n_12555),
.B(n_1679),
.Y(n_13549)
);

OAI21xp5_ASAP7_75t_L g13550 ( 
.A1(n_13209),
.A2(n_13137),
.B(n_13124),
.Y(n_13550)
);

INVx1_ASAP7_75t_SL g13551 ( 
.A(n_12767),
.Y(n_13551)
);

AOI21xp5_ASAP7_75t_L g13552 ( 
.A1(n_13087),
.A2(n_1680),
.B(n_1681),
.Y(n_13552)
);

AO31x2_ASAP7_75t_L g13553 ( 
.A1(n_13132),
.A2(n_1682),
.A3(n_1680),
.B(n_1681),
.Y(n_13553)
);

NAND2xp5_ASAP7_75t_L g13554 ( 
.A(n_12770),
.B(n_1682),
.Y(n_13554)
);

AOI21xp5_ASAP7_75t_L g13555 ( 
.A1(n_13272),
.A2(n_1683),
.B(n_1684),
.Y(n_13555)
);

NAND2xp5_ASAP7_75t_L g13556 ( 
.A(n_12771),
.B(n_1685),
.Y(n_13556)
);

AO31x2_ASAP7_75t_L g13557 ( 
.A1(n_13141),
.A2(n_1687),
.A3(n_1685),
.B(n_1686),
.Y(n_13557)
);

AOI21xp5_ASAP7_75t_L g13558 ( 
.A1(n_12644),
.A2(n_1686),
.B(n_1687),
.Y(n_13558)
);

NOR4xp25_ASAP7_75t_L g13559 ( 
.A(n_12549),
.B(n_13177),
.C(n_13159),
.D(n_13212),
.Y(n_13559)
);

AO21x2_ASAP7_75t_L g13560 ( 
.A1(n_12584),
.A2(n_1688),
.B(n_1689),
.Y(n_13560)
);

OAI21xp5_ASAP7_75t_L g13561 ( 
.A1(n_13144),
.A2(n_1688),
.B(n_1689),
.Y(n_13561)
);

O2A1O1Ixp5_ASAP7_75t_L g13562 ( 
.A1(n_13250),
.A2(n_1692),
.B(n_1690),
.C(n_1691),
.Y(n_13562)
);

NAND2xp5_ASAP7_75t_L g13563 ( 
.A(n_13101),
.B(n_1690),
.Y(n_13563)
);

OAI21x1_ASAP7_75t_L g13564 ( 
.A1(n_12687),
.A2(n_1691),
.B(n_1692),
.Y(n_13564)
);

AND2x2_ASAP7_75t_L g13565 ( 
.A(n_12701),
.B(n_1693),
.Y(n_13565)
);

AO31x2_ASAP7_75t_L g13566 ( 
.A1(n_13105),
.A2(n_1695),
.A3(n_1693),
.B(n_1694),
.Y(n_13566)
);

AOI21xp5_ASAP7_75t_L g13567 ( 
.A1(n_13148),
.A2(n_1694),
.B(n_1695),
.Y(n_13567)
);

OA21x2_ASAP7_75t_L g13568 ( 
.A1(n_12588),
.A2(n_1696),
.B(n_1697),
.Y(n_13568)
);

INVx2_ASAP7_75t_L g13569 ( 
.A(n_12623),
.Y(n_13569)
);

NAND2xp5_ASAP7_75t_L g13570 ( 
.A(n_12924),
.B(n_1696),
.Y(n_13570)
);

INVx2_ASAP7_75t_L g13571 ( 
.A(n_12624),
.Y(n_13571)
);

INVx1_ASAP7_75t_L g13572 ( 
.A(n_12625),
.Y(n_13572)
);

AND2x2_ASAP7_75t_L g13573 ( 
.A(n_12740),
.B(n_1697),
.Y(n_13573)
);

INVx3_ASAP7_75t_L g13574 ( 
.A(n_12913),
.Y(n_13574)
);

NAND3xp33_ASAP7_75t_L g13575 ( 
.A(n_13235),
.B(n_1698),
.C(n_1699),
.Y(n_13575)
);

A2O1A1Ixp33_ASAP7_75t_L g13576 ( 
.A1(n_12778),
.A2(n_1700),
.B(n_1698),
.C(n_1699),
.Y(n_13576)
);

NAND2xp5_ASAP7_75t_L g13577 ( 
.A(n_12927),
.B(n_1700),
.Y(n_13577)
);

INVx3_ASAP7_75t_SL g13578 ( 
.A(n_12978),
.Y(n_13578)
);

AOI221x1_ASAP7_75t_L g13579 ( 
.A1(n_13172),
.A2(n_1703),
.B1(n_1701),
.B2(n_1702),
.C(n_1704),
.Y(n_13579)
);

INVx1_ASAP7_75t_L g13580 ( 
.A(n_12627),
.Y(n_13580)
);

AO21x1_ASAP7_75t_L g13581 ( 
.A1(n_12638),
.A2(n_1701),
.B(n_1703),
.Y(n_13581)
);

NAND2xp5_ASAP7_75t_L g13582 ( 
.A(n_12820),
.B(n_1704),
.Y(n_13582)
);

A2O1A1Ixp33_ASAP7_75t_L g13583 ( 
.A1(n_12899),
.A2(n_1707),
.B(n_1705),
.C(n_1706),
.Y(n_13583)
);

INVx4_ASAP7_75t_L g13584 ( 
.A(n_12553),
.Y(n_13584)
);

AOI22xp5_ASAP7_75t_L g13585 ( 
.A1(n_13274),
.A2(n_1708),
.B1(n_1705),
.B2(n_1706),
.Y(n_13585)
);

AOI221x1_ASAP7_75t_L g13586 ( 
.A1(n_12573),
.A2(n_1711),
.B1(n_1709),
.B2(n_1710),
.C(n_1712),
.Y(n_13586)
);

O2A1O1Ixp33_ASAP7_75t_SL g13587 ( 
.A1(n_13211),
.A2(n_1711),
.B(n_1709),
.C(n_1710),
.Y(n_13587)
);

AOI22xp5_ASAP7_75t_L g13588 ( 
.A1(n_13270),
.A2(n_1714),
.B1(n_1712),
.B2(n_1713),
.Y(n_13588)
);

O2A1O1Ixp33_ASAP7_75t_SL g13589 ( 
.A1(n_12965),
.A2(n_1716),
.B(n_1713),
.C(n_1715),
.Y(n_13589)
);

AND2x2_ASAP7_75t_L g13590 ( 
.A(n_12932),
.B(n_1715),
.Y(n_13590)
);

NOR2xp67_ASAP7_75t_L g13591 ( 
.A(n_12780),
.B(n_1716),
.Y(n_13591)
);

OR2x2_ASAP7_75t_L g13592 ( 
.A(n_12620),
.B(n_1717),
.Y(n_13592)
);

NOR2xp33_ASAP7_75t_L g13593 ( 
.A(n_12843),
.B(n_1717),
.Y(n_13593)
);

INVx1_ASAP7_75t_L g13594 ( 
.A(n_12628),
.Y(n_13594)
);

A2O1A1Ixp33_ASAP7_75t_L g13595 ( 
.A1(n_12524),
.A2(n_1720),
.B(n_1718),
.C(n_1719),
.Y(n_13595)
);

A2O1A1Ixp33_ASAP7_75t_L g13596 ( 
.A1(n_12665),
.A2(n_12831),
.B(n_13257),
.C(n_13254),
.Y(n_13596)
);

INVx1_ASAP7_75t_L g13597 ( 
.A(n_12631),
.Y(n_13597)
);

NAND2xp5_ASAP7_75t_L g13598 ( 
.A(n_12821),
.B(n_1719),
.Y(n_13598)
);

BUFx6f_ASAP7_75t_L g13599 ( 
.A(n_12585),
.Y(n_13599)
);

A2O1A1Ixp33_ASAP7_75t_L g13600 ( 
.A1(n_13271),
.A2(n_1723),
.B(n_1721),
.C(n_1722),
.Y(n_13600)
);

AOI22xp5_ASAP7_75t_L g13601 ( 
.A1(n_13270),
.A2(n_1723),
.B1(n_1721),
.B2(n_1722),
.Y(n_13601)
);

NOR2xp33_ASAP7_75t_L g13602 ( 
.A(n_12903),
.B(n_1724),
.Y(n_13602)
);

OAI21xp5_ASAP7_75t_L g13603 ( 
.A1(n_13153),
.A2(n_13162),
.B(n_13154),
.Y(n_13603)
);

AO32x2_ASAP7_75t_L g13604 ( 
.A1(n_13008),
.A2(n_1727),
.A3(n_1725),
.B1(n_1726),
.B2(n_1728),
.Y(n_13604)
);

AOI22xp5_ASAP7_75t_L g13605 ( 
.A1(n_12739),
.A2(n_12984),
.B1(n_12873),
.B2(n_13064),
.Y(n_13605)
);

OAI22x1_ASAP7_75t_L g13606 ( 
.A1(n_13096),
.A2(n_1727),
.B1(n_1725),
.B2(n_1726),
.Y(n_13606)
);

AOI21xp5_ASAP7_75t_L g13607 ( 
.A1(n_13170),
.A2(n_13184),
.B(n_13182),
.Y(n_13607)
);

INVx3_ASAP7_75t_L g13608 ( 
.A(n_12585),
.Y(n_13608)
);

NOR2xp33_ASAP7_75t_L g13609 ( 
.A(n_12531),
.B(n_1728),
.Y(n_13609)
);

OAI21xp5_ASAP7_75t_L g13610 ( 
.A1(n_13190),
.A2(n_1729),
.B(n_1730),
.Y(n_13610)
);

NAND2xp5_ASAP7_75t_L g13611 ( 
.A(n_12830),
.B(n_1729),
.Y(n_13611)
);

BUFx8_ASAP7_75t_SL g13612 ( 
.A(n_12757),
.Y(n_13612)
);

OAI21xp5_ASAP7_75t_L g13613 ( 
.A1(n_13196),
.A2(n_1730),
.B(n_1731),
.Y(n_13613)
);

BUFx6f_ASAP7_75t_L g13614 ( 
.A(n_12716),
.Y(n_13614)
);

AOI21xp5_ASAP7_75t_L g13615 ( 
.A1(n_13198),
.A2(n_1732),
.B(n_1733),
.Y(n_13615)
);

AOI21x1_ASAP7_75t_L g13616 ( 
.A1(n_12918),
.A2(n_1732),
.B(n_1734),
.Y(n_13616)
);

OAI21xp5_ASAP7_75t_L g13617 ( 
.A1(n_13204),
.A2(n_13219),
.B(n_13214),
.Y(n_13617)
);

AND2x2_ASAP7_75t_L g13618 ( 
.A(n_12586),
.B(n_1734),
.Y(n_13618)
);

AOI21xp5_ASAP7_75t_L g13619 ( 
.A1(n_13228),
.A2(n_1735),
.B(n_1736),
.Y(n_13619)
);

O2A1O1Ixp5_ASAP7_75t_L g13620 ( 
.A1(n_13173),
.A2(n_1737),
.B(n_1735),
.C(n_1736),
.Y(n_13620)
);

AO31x2_ASAP7_75t_L g13621 ( 
.A1(n_13203),
.A2(n_1739),
.A3(n_1737),
.B(n_1738),
.Y(n_13621)
);

NOR2xp33_ASAP7_75t_SL g13622 ( 
.A(n_12634),
.B(n_1738),
.Y(n_13622)
);

OAI21x1_ASAP7_75t_L g13623 ( 
.A1(n_13197),
.A2(n_1739),
.B(n_1740),
.Y(n_13623)
);

NAND2x1_ASAP7_75t_L g13624 ( 
.A(n_12683),
.B(n_1741),
.Y(n_13624)
);

OAI21x1_ASAP7_75t_L g13625 ( 
.A1(n_13103),
.A2(n_1741),
.B(n_1742),
.Y(n_13625)
);

OAI21x1_ASAP7_75t_L g13626 ( 
.A1(n_12556),
.A2(n_1742),
.B(n_1743),
.Y(n_13626)
);

OAI21x1_ASAP7_75t_L g13627 ( 
.A1(n_13255),
.A2(n_1744),
.B(n_1745),
.Y(n_13627)
);

AOI21xp5_ASAP7_75t_L g13628 ( 
.A1(n_12679),
.A2(n_1744),
.B(n_1746),
.Y(n_13628)
);

AO32x2_ASAP7_75t_L g13629 ( 
.A1(n_12956),
.A2(n_12789),
.A3(n_12769),
.B1(n_12596),
.B2(n_13266),
.Y(n_13629)
);

NOR2xp33_ASAP7_75t_L g13630 ( 
.A(n_12876),
.B(n_1746),
.Y(n_13630)
);

AOI21xp5_ASAP7_75t_L g13631 ( 
.A1(n_12833),
.A2(n_1747),
.B(n_1748),
.Y(n_13631)
);

OAI21xp5_ASAP7_75t_L g13632 ( 
.A1(n_13263),
.A2(n_1748),
.B(n_1749),
.Y(n_13632)
);

AOI21xp5_ASAP7_75t_L g13633 ( 
.A1(n_12857),
.A2(n_1750),
.B(n_1751),
.Y(n_13633)
);

NAND2xp5_ASAP7_75t_SL g13634 ( 
.A(n_13110),
.B(n_1750),
.Y(n_13634)
);

BUFx6f_ASAP7_75t_L g13635 ( 
.A(n_12716),
.Y(n_13635)
);

OAI22xp5_ASAP7_75t_L g13636 ( 
.A1(n_12635),
.A2(n_1753),
.B1(n_1751),
.B2(n_1752),
.Y(n_13636)
);

OAI21xp5_ASAP7_75t_L g13637 ( 
.A1(n_12966),
.A2(n_1752),
.B(n_1753),
.Y(n_13637)
);

INVx2_ASAP7_75t_L g13638 ( 
.A(n_12849),
.Y(n_13638)
);

AOI21x1_ASAP7_75t_L g13639 ( 
.A1(n_12551),
.A2(n_1754),
.B(n_1755),
.Y(n_13639)
);

AOI21xp5_ASAP7_75t_L g13640 ( 
.A1(n_13259),
.A2(n_1754),
.B(n_1756),
.Y(n_13640)
);

AO22x2_ASAP7_75t_L g13641 ( 
.A1(n_13072),
.A2(n_1758),
.B1(n_1756),
.B2(n_1757),
.Y(n_13641)
);

NOR2xp67_ASAP7_75t_SL g13642 ( 
.A(n_12729),
.B(n_1757),
.Y(n_13642)
);

INVx1_ASAP7_75t_L g13643 ( 
.A(n_12832),
.Y(n_13643)
);

AO31x2_ASAP7_75t_L g13644 ( 
.A1(n_13181),
.A2(n_1760),
.A3(n_1758),
.B(n_1759),
.Y(n_13644)
);

OAI21x1_ASAP7_75t_L g13645 ( 
.A1(n_13264),
.A2(n_1759),
.B(n_1760),
.Y(n_13645)
);

AO31x2_ASAP7_75t_L g13646 ( 
.A1(n_13278),
.A2(n_1763),
.A3(n_1761),
.B(n_1762),
.Y(n_13646)
);

A2O1A1Ixp33_ASAP7_75t_L g13647 ( 
.A1(n_13213),
.A2(n_1763),
.B(n_1761),
.C(n_1762),
.Y(n_13647)
);

AND2x4_ASAP7_75t_L g13648 ( 
.A(n_12854),
.B(n_1764),
.Y(n_13648)
);

CKINVDCx16_ASAP7_75t_R g13649 ( 
.A(n_12615),
.Y(n_13649)
);

AND2x2_ASAP7_75t_L g13650 ( 
.A(n_12785),
.B(n_1764),
.Y(n_13650)
);

AND2x2_ASAP7_75t_L g13651 ( 
.A(n_12798),
.B(n_12897),
.Y(n_13651)
);

BUFx2_ASAP7_75t_L g13652 ( 
.A(n_12860),
.Y(n_13652)
);

OAI21x1_ASAP7_75t_L g13653 ( 
.A1(n_12598),
.A2(n_1765),
.B(n_1766),
.Y(n_13653)
);

NOR2x1_ASAP7_75t_SL g13654 ( 
.A(n_13130),
.B(n_1765),
.Y(n_13654)
);

AOI21xp5_ASAP7_75t_L g13655 ( 
.A1(n_13114),
.A2(n_1766),
.B(n_1767),
.Y(n_13655)
);

BUFx3_ASAP7_75t_L g13656 ( 
.A(n_12756),
.Y(n_13656)
);

OAI21x1_ASAP7_75t_L g13657 ( 
.A1(n_12599),
.A2(n_1767),
.B(n_1768),
.Y(n_13657)
);

AO31x2_ASAP7_75t_L g13658 ( 
.A1(n_13277),
.A2(n_13282),
.A3(n_13279),
.B(n_12848),
.Y(n_13658)
);

AO31x2_ASAP7_75t_L g13659 ( 
.A1(n_12838),
.A2(n_1771),
.A3(n_1769),
.B(n_1770),
.Y(n_13659)
);

BUFx3_ASAP7_75t_L g13660 ( 
.A(n_12751),
.Y(n_13660)
);

INVx1_ASAP7_75t_L g13661 ( 
.A(n_12859),
.Y(n_13661)
);

INVx1_ASAP7_75t_L g13662 ( 
.A(n_12874),
.Y(n_13662)
);

NAND2xp5_ASAP7_75t_L g13663 ( 
.A(n_12879),
.B(n_1769),
.Y(n_13663)
);

AOI221x1_ASAP7_75t_L g13664 ( 
.A1(n_13107),
.A2(n_1772),
.B1(n_1770),
.B2(n_1771),
.C(n_1773),
.Y(n_13664)
);

AOI22xp5_ASAP7_75t_L g13665 ( 
.A1(n_12984),
.A2(n_1774),
.B1(n_1772),
.B2(n_1773),
.Y(n_13665)
);

O2A1O1Ixp33_ASAP7_75t_SL g13666 ( 
.A1(n_12988),
.A2(n_1776),
.B(n_1774),
.C(n_1775),
.Y(n_13666)
);

A2O1A1Ixp33_ASAP7_75t_L g13667 ( 
.A1(n_12986),
.A2(n_1777),
.B(n_1775),
.C(n_1776),
.Y(n_13667)
);

INVx2_ASAP7_75t_L g13668 ( 
.A(n_12862),
.Y(n_13668)
);

A2O1A1Ixp33_ASAP7_75t_L g13669 ( 
.A1(n_13251),
.A2(n_1780),
.B(n_1778),
.C(n_1779),
.Y(n_13669)
);

A2O1A1Ixp33_ASAP7_75t_L g13670 ( 
.A1(n_13256),
.A2(n_1782),
.B(n_1779),
.C(n_1781),
.Y(n_13670)
);

OAI21x1_ASAP7_75t_L g13671 ( 
.A1(n_12601),
.A2(n_1781),
.B(n_1782),
.Y(n_13671)
);

INVx1_ASAP7_75t_L g13672 ( 
.A(n_12885),
.Y(n_13672)
);

NAND2xp5_ASAP7_75t_L g13673 ( 
.A(n_12886),
.B(n_1784),
.Y(n_13673)
);

NAND2x1p5_ASAP7_75t_L g13674 ( 
.A(n_12619),
.B(n_1784),
.Y(n_13674)
);

AOI21x1_ASAP7_75t_L g13675 ( 
.A1(n_13260),
.A2(n_1785),
.B(n_1787),
.Y(n_13675)
);

OAI21xp5_ASAP7_75t_L g13676 ( 
.A1(n_13016),
.A2(n_1785),
.B(n_1787),
.Y(n_13676)
);

INVx1_ASAP7_75t_L g13677 ( 
.A(n_12892),
.Y(n_13677)
);

OAI21xp5_ASAP7_75t_L g13678 ( 
.A1(n_12593),
.A2(n_1788),
.B(n_1789),
.Y(n_13678)
);

INVx3_ASAP7_75t_L g13679 ( 
.A(n_12730),
.Y(n_13679)
);

OAI21x1_ASAP7_75t_L g13680 ( 
.A1(n_12607),
.A2(n_1788),
.B(n_1789),
.Y(n_13680)
);

NOR2xp33_ASAP7_75t_L g13681 ( 
.A(n_12910),
.B(n_1790),
.Y(n_13681)
);

OAI21xp5_ASAP7_75t_L g13682 ( 
.A1(n_13117),
.A2(n_1791),
.B(n_1792),
.Y(n_13682)
);

NAND2xp5_ASAP7_75t_L g13683 ( 
.A(n_12893),
.B(n_1791),
.Y(n_13683)
);

OA21x2_ASAP7_75t_L g13684 ( 
.A1(n_12530),
.A2(n_1793),
.B(n_1794),
.Y(n_13684)
);

A2O1A1Ixp33_ASAP7_75t_L g13685 ( 
.A1(n_13267),
.A2(n_1795),
.B(n_1793),
.C(n_1794),
.Y(n_13685)
);

AOI21xp5_ASAP7_75t_L g13686 ( 
.A1(n_12790),
.A2(n_1795),
.B(n_1796),
.Y(n_13686)
);

AOI21xp5_ASAP7_75t_L g13687 ( 
.A1(n_12880),
.A2(n_1796),
.B(n_1797),
.Y(n_13687)
);

CKINVDCx11_ASAP7_75t_R g13688 ( 
.A(n_13031),
.Y(n_13688)
);

INVx1_ASAP7_75t_SL g13689 ( 
.A(n_13054),
.Y(n_13689)
);

BUFx6f_ASAP7_75t_L g13690 ( 
.A(n_12730),
.Y(n_13690)
);

NOR2xp33_ASAP7_75t_SL g13691 ( 
.A(n_12562),
.B(n_1797),
.Y(n_13691)
);

A2O1A1Ixp33_ASAP7_75t_L g13692 ( 
.A1(n_12948),
.A2(n_1800),
.B(n_1798),
.C(n_1799),
.Y(n_13692)
);

OA21x2_ASAP7_75t_L g13693 ( 
.A1(n_12532),
.A2(n_1798),
.B(n_1799),
.Y(n_13693)
);

INVx1_ASAP7_75t_L g13694 ( 
.A(n_12902),
.Y(n_13694)
);

AOI21xp5_ASAP7_75t_L g13695 ( 
.A1(n_13115),
.A2(n_1800),
.B(n_1801),
.Y(n_13695)
);

INVx1_ASAP7_75t_L g13696 ( 
.A(n_12905),
.Y(n_13696)
);

OR2x2_ASAP7_75t_L g13697 ( 
.A(n_12915),
.B(n_12916),
.Y(n_13697)
);

OAI22xp5_ASAP7_75t_L g13698 ( 
.A1(n_13245),
.A2(n_1803),
.B1(n_1801),
.B2(n_1802),
.Y(n_13698)
);

O2A1O1Ixp5_ASAP7_75t_L g13699 ( 
.A1(n_12622),
.A2(n_1805),
.B(n_1802),
.C(n_1804),
.Y(n_13699)
);

OAI21xp5_ASAP7_75t_L g13700 ( 
.A1(n_12963),
.A2(n_1804),
.B(n_1805),
.Y(n_13700)
);

A2O1A1Ixp33_ASAP7_75t_L g13701 ( 
.A1(n_13112),
.A2(n_1808),
.B(n_1806),
.C(n_1807),
.Y(n_13701)
);

AND2x2_ASAP7_75t_L g13702 ( 
.A(n_13058),
.B(n_1808),
.Y(n_13702)
);

OAI22xp5_ASAP7_75t_L g13703 ( 
.A1(n_12861),
.A2(n_1811),
.B1(n_1809),
.B2(n_1810),
.Y(n_13703)
);

OAI21x1_ASAP7_75t_SL g13704 ( 
.A1(n_12533),
.A2(n_1809),
.B(n_1810),
.Y(n_13704)
);

INVxp67_ASAP7_75t_L g13705 ( 
.A(n_12741),
.Y(n_13705)
);

NAND3xp33_ASAP7_75t_L g13706 ( 
.A(n_13156),
.B(n_1812),
.C(n_1813),
.Y(n_13706)
);

INVx1_ASAP7_75t_SL g13707 ( 
.A(n_12787),
.Y(n_13707)
);

AOI21xp5_ASAP7_75t_L g13708 ( 
.A1(n_13194),
.A2(n_1812),
.B(n_1813),
.Y(n_13708)
);

O2A1O1Ixp33_ASAP7_75t_L g13709 ( 
.A1(n_12719),
.A2(n_1816),
.B(n_1814),
.C(n_1815),
.Y(n_13709)
);

AO31x2_ASAP7_75t_L g13710 ( 
.A1(n_12923),
.A2(n_1816),
.A3(n_1814),
.B(n_1815),
.Y(n_13710)
);

A2O1A1Ixp33_ASAP7_75t_L g13711 ( 
.A1(n_13240),
.A2(n_1819),
.B(n_1817),
.C(n_1818),
.Y(n_13711)
);

AO32x2_ASAP7_75t_L g13712 ( 
.A1(n_13052),
.A2(n_1821),
.A3(n_1819),
.B1(n_1820),
.B2(n_1822),
.Y(n_13712)
);

BUFx2_ASAP7_75t_L g13713 ( 
.A(n_12866),
.Y(n_13713)
);

AOI21xp33_ASAP7_75t_L g13714 ( 
.A1(n_13281),
.A2(n_1820),
.B(n_1822),
.Y(n_13714)
);

AOI21xp5_ASAP7_75t_L g13715 ( 
.A1(n_13232),
.A2(n_1823),
.B(n_1824),
.Y(n_13715)
);

NOR2xp33_ASAP7_75t_SL g13716 ( 
.A(n_12603),
.B(n_1823),
.Y(n_13716)
);

NOR2x1_ASAP7_75t_SL g13717 ( 
.A(n_13130),
.B(n_1824),
.Y(n_13717)
);

AND2x2_ASAP7_75t_L g13718 ( 
.A(n_12982),
.B(n_12814),
.Y(n_13718)
);

A2O1A1Ixp33_ASAP7_75t_L g13719 ( 
.A1(n_13142),
.A2(n_1827),
.B(n_1825),
.C(n_1826),
.Y(n_13719)
);

NAND2xp5_ASAP7_75t_L g13720 ( 
.A(n_12931),
.B(n_12935),
.Y(n_13720)
);

AOI21xp5_ASAP7_75t_L g13721 ( 
.A1(n_13049),
.A2(n_1825),
.B(n_1826),
.Y(n_13721)
);

AOI221xp5_ASAP7_75t_SL g13722 ( 
.A1(n_13041),
.A2(n_1830),
.B1(n_1828),
.B2(n_1829),
.C(n_1831),
.Y(n_13722)
);

NOR2xp33_ASAP7_75t_L g13723 ( 
.A(n_12825),
.B(n_12936),
.Y(n_13723)
);

OR2x2_ASAP7_75t_L g13724 ( 
.A(n_12937),
.B(n_1828),
.Y(n_13724)
);

AO21x2_ASAP7_75t_L g13725 ( 
.A1(n_12560),
.A2(n_1829),
.B(n_1830),
.Y(n_13725)
);

AND2x2_ASAP7_75t_L g13726 ( 
.A(n_12964),
.B(n_1831),
.Y(n_13726)
);

OR2x2_ASAP7_75t_L g13727 ( 
.A(n_12938),
.B(n_1832),
.Y(n_13727)
);

AO31x2_ASAP7_75t_L g13728 ( 
.A1(n_12941),
.A2(n_1834),
.A3(n_1832),
.B(n_1833),
.Y(n_13728)
);

NAND2xp5_ASAP7_75t_L g13729 ( 
.A(n_13068),
.B(n_1833),
.Y(n_13729)
);

AO21x2_ASAP7_75t_L g13730 ( 
.A1(n_12554),
.A2(n_1834),
.B(n_1835),
.Y(n_13730)
);

AOI21xp5_ASAP7_75t_L g13731 ( 
.A1(n_13261),
.A2(n_1835),
.B(n_1836),
.Y(n_13731)
);

OR2x2_ASAP7_75t_L g13732 ( 
.A(n_13076),
.B(n_13078),
.Y(n_13732)
);

AOI21xp5_ASAP7_75t_L g13733 ( 
.A1(n_12962),
.A2(n_1837),
.B(n_1838),
.Y(n_13733)
);

INVx2_ASAP7_75t_L g13734 ( 
.A(n_12881),
.Y(n_13734)
);

NOR2xp33_ASAP7_75t_L g13735 ( 
.A(n_13080),
.B(n_1837),
.Y(n_13735)
);

OAI21xp5_ASAP7_75t_L g13736 ( 
.A1(n_12984),
.A2(n_1839),
.B(n_1840),
.Y(n_13736)
);

INVx8_ASAP7_75t_L g13737 ( 
.A(n_12925),
.Y(n_13737)
);

AOI22xp5_ASAP7_75t_L g13738 ( 
.A1(n_12565),
.A2(n_1841),
.B1(n_1839),
.B2(n_1840),
.Y(n_13738)
);

A2O1A1Ixp33_ASAP7_75t_L g13739 ( 
.A1(n_13273),
.A2(n_1843),
.B(n_1841),
.C(n_1842),
.Y(n_13739)
);

NAND2xp5_ASAP7_75t_L g13740 ( 
.A(n_13174),
.B(n_1842),
.Y(n_13740)
);

BUFx2_ASAP7_75t_L g13741 ( 
.A(n_12811),
.Y(n_13741)
);

A2O1A1Ixp33_ASAP7_75t_L g13742 ( 
.A1(n_13275),
.A2(n_1845),
.B(n_1843),
.C(n_1844),
.Y(n_13742)
);

INVx1_ASAP7_75t_L g13743 ( 
.A(n_12536),
.Y(n_13743)
);

INVx2_ASAP7_75t_L g13744 ( 
.A(n_12900),
.Y(n_13744)
);

CKINVDCx20_ASAP7_75t_R g13745 ( 
.A(n_12777),
.Y(n_13745)
);

AOI21xp5_ASAP7_75t_L g13746 ( 
.A1(n_13089),
.A2(n_1845),
.B(n_1846),
.Y(n_13746)
);

INVx4_ASAP7_75t_L g13747 ( 
.A(n_12791),
.Y(n_13747)
);

AO31x2_ASAP7_75t_L g13748 ( 
.A1(n_13236),
.A2(n_1848),
.A3(n_1846),
.B(n_1847),
.Y(n_13748)
);

NOR2xp33_ASAP7_75t_L g13749 ( 
.A(n_13073),
.B(n_12955),
.Y(n_13749)
);

OAI21x1_ASAP7_75t_L g13750 ( 
.A1(n_13220),
.A2(n_1847),
.B(n_1848),
.Y(n_13750)
);

AOI21xp5_ASAP7_75t_L g13751 ( 
.A1(n_13092),
.A2(n_1849),
.B(n_1850),
.Y(n_13751)
);

OA21x2_ASAP7_75t_L g13752 ( 
.A1(n_12534),
.A2(n_1849),
.B(n_1850),
.Y(n_13752)
);

INVx2_ASAP7_75t_SL g13753 ( 
.A(n_12850),
.Y(n_13753)
);

NOR4xp25_ASAP7_75t_L g13754 ( 
.A(n_12920),
.B(n_1853),
.C(n_1851),
.D(n_1852),
.Y(n_13754)
);

NOR2xp33_ASAP7_75t_SL g13755 ( 
.A(n_12972),
.B(n_12772),
.Y(n_13755)
);

AOI21xp5_ASAP7_75t_L g13756 ( 
.A1(n_13097),
.A2(n_1851),
.B(n_1853),
.Y(n_13756)
);

INVx4_ASAP7_75t_L g13757 ( 
.A(n_12901),
.Y(n_13757)
);

CKINVDCx5p33_ASAP7_75t_R g13758 ( 
.A(n_12728),
.Y(n_13758)
);

BUFx12f_ASAP7_75t_L g13759 ( 
.A(n_12909),
.Y(n_13759)
);

INVx2_ASAP7_75t_L g13760 ( 
.A(n_12911),
.Y(n_13760)
);

OAI21x1_ASAP7_75t_L g13761 ( 
.A1(n_13238),
.A2(n_1854),
.B(n_1855),
.Y(n_13761)
);

OAI22xp5_ASAP7_75t_L g13762 ( 
.A1(n_12967),
.A2(n_1856),
.B1(n_1854),
.B2(n_1855),
.Y(n_13762)
);

AOI21xp5_ASAP7_75t_L g13763 ( 
.A1(n_13098),
.A2(n_1856),
.B(n_1857),
.Y(n_13763)
);

INVx3_ASAP7_75t_SL g13764 ( 
.A(n_13074),
.Y(n_13764)
);

INVx3_ASAP7_75t_L g13765 ( 
.A(n_12796),
.Y(n_13765)
);

AOI21xp5_ASAP7_75t_L g13766 ( 
.A1(n_13099),
.A2(n_1857),
.B(n_1858),
.Y(n_13766)
);

INVx8_ASAP7_75t_L g13767 ( 
.A(n_12759),
.Y(n_13767)
);

INVx2_ASAP7_75t_L g13768 ( 
.A(n_12951),
.Y(n_13768)
);

INVxp67_ASAP7_75t_SL g13769 ( 
.A(n_13164),
.Y(n_13769)
);

O2A1O1Ixp33_ASAP7_75t_SL g13770 ( 
.A1(n_12742),
.A2(n_1860),
.B(n_1858),
.C(n_1859),
.Y(n_13770)
);

INVx1_ASAP7_75t_L g13771 ( 
.A(n_12618),
.Y(n_13771)
);

NOR2xp33_ASAP7_75t_L g13772 ( 
.A(n_13073),
.B(n_1859),
.Y(n_13772)
);

INVx1_ASAP7_75t_SL g13773 ( 
.A(n_12720),
.Y(n_13773)
);

AO31x2_ASAP7_75t_L g13774 ( 
.A1(n_13244),
.A2(n_1862),
.A3(n_1860),
.B(n_1861),
.Y(n_13774)
);

OAI21xp5_ASAP7_75t_L g13775 ( 
.A1(n_12753),
.A2(n_1861),
.B(n_1862),
.Y(n_13775)
);

INVx3_ASAP7_75t_SL g13776 ( 
.A(n_13082),
.Y(n_13776)
);

AOI21x1_ASAP7_75t_L g13777 ( 
.A1(n_12621),
.A2(n_1863),
.B(n_1864),
.Y(n_13777)
);

OR2x6_ASAP7_75t_L g13778 ( 
.A(n_13020),
.B(n_1863),
.Y(n_13778)
);

OAI22xp5_ASAP7_75t_L g13779 ( 
.A1(n_13163),
.A2(n_13191),
.B1(n_13206),
.B2(n_13188),
.Y(n_13779)
);

NAND2xp5_ASAP7_75t_L g13780 ( 
.A(n_13168),
.B(n_1864),
.Y(n_13780)
);

NAND2xp5_ASAP7_75t_L g13781 ( 
.A(n_13186),
.B(n_1865),
.Y(n_13781)
);

AOI21x1_ASAP7_75t_L g13782 ( 
.A1(n_12626),
.A2(n_1865),
.B(n_1866),
.Y(n_13782)
);

O2A1O1Ixp33_ASAP7_75t_L g13783 ( 
.A1(n_13102),
.A2(n_13108),
.B(n_12856),
.C(n_12839),
.Y(n_13783)
);

AO21x1_ASAP7_75t_L g13784 ( 
.A1(n_12526),
.A2(n_1866),
.B(n_1867),
.Y(n_13784)
);

A2O1A1Ixp33_ASAP7_75t_L g13785 ( 
.A1(n_13201),
.A2(n_1869),
.B(n_1867),
.C(n_1868),
.Y(n_13785)
);

OAI22xp5_ASAP7_75t_L g13786 ( 
.A1(n_13207),
.A2(n_13237),
.B1(n_12803),
.B2(n_12993),
.Y(n_13786)
);

AOI31xp67_ASAP7_75t_L g13787 ( 
.A1(n_13145),
.A2(n_1870),
.A3(n_1868),
.B(n_1869),
.Y(n_13787)
);

NOR2xp33_ASAP7_75t_L g13788 ( 
.A(n_13091),
.B(n_13094),
.Y(n_13788)
);

NAND2xp5_ASAP7_75t_L g13789 ( 
.A(n_13187),
.B(n_1871),
.Y(n_13789)
);

NAND2xp5_ASAP7_75t_L g13790 ( 
.A(n_12569),
.B(n_1871),
.Y(n_13790)
);

A2O1A1Ixp33_ASAP7_75t_L g13791 ( 
.A1(n_13210),
.A2(n_1875),
.B(n_1872),
.C(n_1873),
.Y(n_13791)
);

A2O1A1Ixp33_ASAP7_75t_L g13792 ( 
.A1(n_12906),
.A2(n_1875),
.B(n_1872),
.C(n_1873),
.Y(n_13792)
);

OAI21x1_ASAP7_75t_L g13793 ( 
.A1(n_12535),
.A2(n_12538),
.B(n_12643),
.Y(n_13793)
);

AO31x2_ASAP7_75t_L g13794 ( 
.A1(n_13265),
.A2(n_1878),
.A3(n_1876),
.B(n_1877),
.Y(n_13794)
);

AOI22xp33_ASAP7_75t_L g13795 ( 
.A1(n_13268),
.A2(n_13269),
.B1(n_12575),
.B2(n_13037),
.Y(n_13795)
);

CKINVDCx5p33_ASAP7_75t_R g13796 ( 
.A(n_12796),
.Y(n_13796)
);

OR2x2_ASAP7_75t_L g13797 ( 
.A(n_12952),
.B(n_1876),
.Y(n_13797)
);

BUFx2_ASAP7_75t_L g13798 ( 
.A(n_12969),
.Y(n_13798)
);

AOI221xp5_ASAP7_75t_L g13799 ( 
.A1(n_13246),
.A2(n_1879),
.B1(n_1877),
.B2(n_1878),
.C(n_1880),
.Y(n_13799)
);

OR2x2_ASAP7_75t_L g13800 ( 
.A(n_12968),
.B(n_1879),
.Y(n_13800)
);

AO31x2_ASAP7_75t_L g13801 ( 
.A1(n_13280),
.A2(n_1882),
.A3(n_1880),
.B(n_1881),
.Y(n_13801)
);

AOI21xp5_ASAP7_75t_L g13802 ( 
.A1(n_13086),
.A2(n_13247),
.B(n_13175),
.Y(n_13802)
);

AOI22xp33_ASAP7_75t_L g13803 ( 
.A1(n_12575),
.A2(n_1883),
.B1(n_1881),
.B2(n_1882),
.Y(n_13803)
);

INVx1_ASAP7_75t_L g13804 ( 
.A(n_12578),
.Y(n_13804)
);

BUFx12f_ASAP7_75t_L g13805 ( 
.A(n_12827),
.Y(n_13805)
);

BUFx3_ASAP7_75t_L g13806 ( 
.A(n_12990),
.Y(n_13806)
);

AOI21xp5_ASAP7_75t_L g13807 ( 
.A1(n_12837),
.A2(n_1883),
.B(n_1884),
.Y(n_13807)
);

O2A1O1Ixp33_ASAP7_75t_SL g13808 ( 
.A1(n_12934),
.A2(n_1886),
.B(n_1884),
.C(n_1885),
.Y(n_13808)
);

AOI221xp5_ASAP7_75t_SL g13809 ( 
.A1(n_12801),
.A2(n_1888),
.B1(n_1885),
.B2(n_1887),
.C(n_1889),
.Y(n_13809)
);

INVx2_ASAP7_75t_SL g13810 ( 
.A(n_12981),
.Y(n_13810)
);

AOI31xp33_ASAP7_75t_L g13811 ( 
.A1(n_12845),
.A2(n_1889),
.A3(n_1887),
.B(n_1888),
.Y(n_13811)
);

AOI21xp5_ASAP7_75t_L g13812 ( 
.A1(n_12664),
.A2(n_1891),
.B(n_1892),
.Y(n_13812)
);

AND2x4_ASAP7_75t_L g13813 ( 
.A(n_12521),
.B(n_1891),
.Y(n_13813)
);

OA21x2_ASAP7_75t_L g13814 ( 
.A1(n_12639),
.A2(n_1892),
.B(n_1893),
.Y(n_13814)
);

OAI21x1_ASAP7_75t_L g13815 ( 
.A1(n_12666),
.A2(n_1894),
.B(n_1895),
.Y(n_13815)
);

INVx1_ASAP7_75t_L g13816 ( 
.A(n_12587),
.Y(n_13816)
);

O2A1O1Ixp33_ASAP7_75t_SL g13817 ( 
.A1(n_12802),
.A2(n_1896),
.B(n_1894),
.C(n_1895),
.Y(n_13817)
);

NAND3xp33_ASAP7_75t_SL g13818 ( 
.A(n_12944),
.B(n_1897),
.C(n_1898),
.Y(n_13818)
);

INVx2_ASAP7_75t_SL g13819 ( 
.A(n_12550),
.Y(n_13819)
);

AO21x1_ASAP7_75t_L g13820 ( 
.A1(n_12645),
.A2(n_1897),
.B(n_1898),
.Y(n_13820)
);

NAND2xp5_ASAP7_75t_L g13821 ( 
.A(n_12589),
.B(n_1899),
.Y(n_13821)
);

NAND2xp5_ASAP7_75t_L g13822 ( 
.A(n_12611),
.B(n_1899),
.Y(n_13822)
);

NAND2xp5_ASAP7_75t_L g13823 ( 
.A(n_12658),
.B(n_1900),
.Y(n_13823)
);

NAND2xp5_ASAP7_75t_L g13824 ( 
.A(n_12708),
.B(n_1900),
.Y(n_13824)
);

BUFx3_ASAP7_75t_L g13825 ( 
.A(n_12990),
.Y(n_13825)
);

A2O1A1Ixp33_ASAP7_75t_L g13826 ( 
.A1(n_13131),
.A2(n_1904),
.B(n_1901),
.C(n_1902),
.Y(n_13826)
);

OAI21xp5_ASAP7_75t_L g13827 ( 
.A1(n_12575),
.A2(n_1901),
.B(n_1905),
.Y(n_13827)
);

BUFx3_ASAP7_75t_L g13828 ( 
.A(n_12995),
.Y(n_13828)
);

AO31x2_ASAP7_75t_L g13829 ( 
.A1(n_13276),
.A2(n_1907),
.A3(n_1905),
.B(n_1906),
.Y(n_13829)
);

OAI22xp5_ASAP7_75t_L g13830 ( 
.A1(n_13199),
.A2(n_1908),
.B1(n_1906),
.B2(n_1907),
.Y(n_13830)
);

BUFx3_ASAP7_75t_L g13831 ( 
.A(n_12995),
.Y(n_13831)
);

BUFx2_ASAP7_75t_L g13832 ( 
.A(n_12871),
.Y(n_13832)
);

BUFx6f_ASAP7_75t_L g13833 ( 
.A(n_12864),
.Y(n_13833)
);

NOR2xp67_ASAP7_75t_L g13834 ( 
.A(n_12786),
.B(n_1908),
.Y(n_13834)
);

AND2x2_ASAP7_75t_SL g13835 ( 
.A(n_13020),
.B(n_13022),
.Y(n_13835)
);

O2A1O1Ixp33_ASAP7_75t_L g13836 ( 
.A1(n_12994),
.A2(n_1911),
.B(n_1909),
.C(n_1910),
.Y(n_13836)
);

A2O1A1Ixp33_ASAP7_75t_L g13837 ( 
.A1(n_13218),
.A2(n_1912),
.B(n_1909),
.C(n_1910),
.Y(n_13837)
);

INVxp67_ASAP7_75t_L g13838 ( 
.A(n_12712),
.Y(n_13838)
);

NOR2x1_ASAP7_75t_SL g13839 ( 
.A(n_13287),
.B(n_12529),
.Y(n_13839)
);

NOR2x1_ASAP7_75t_SL g13840 ( 
.A(n_13417),
.B(n_12656),
.Y(n_13840)
);

OAI21x1_ASAP7_75t_L g13841 ( 
.A1(n_13488),
.A2(n_12674),
.B(n_12673),
.Y(n_13841)
);

AND2x4_ASAP7_75t_L g13842 ( 
.A(n_13434),
.B(n_13057),
.Y(n_13842)
);

OAI22xp33_ASAP7_75t_L g13843 ( 
.A1(n_13490),
.A2(n_13067),
.B1(n_12805),
.B2(n_12921),
.Y(n_13843)
);

OAI21x1_ASAP7_75t_L g13844 ( 
.A1(n_13389),
.A2(n_12688),
.B(n_12677),
.Y(n_13844)
);

NOR2xp33_ASAP7_75t_L g13845 ( 
.A(n_13423),
.B(n_12846),
.Y(n_13845)
);

OAI21xp5_ASAP7_75t_L g13846 ( 
.A1(n_13313),
.A2(n_12922),
.B(n_12829),
.Y(n_13846)
);

HB1xp67_ASAP7_75t_L g13847 ( 
.A(n_13658),
.Y(n_13847)
);

OAI21x1_ASAP7_75t_L g13848 ( 
.A1(n_13324),
.A2(n_12692),
.B(n_12689),
.Y(n_13848)
);

AND2x2_ASAP7_75t_L g13849 ( 
.A(n_13367),
.B(n_12974),
.Y(n_13849)
);

OR2x6_ASAP7_75t_L g13850 ( 
.A(n_13337),
.B(n_13289),
.Y(n_13850)
);

INVx1_ASAP7_75t_L g13851 ( 
.A(n_13522),
.Y(n_13851)
);

AND2x4_ASAP7_75t_L g13852 ( 
.A(n_13769),
.B(n_12743),
.Y(n_13852)
);

INVx6_ASAP7_75t_L g13853 ( 
.A(n_13466),
.Y(n_13853)
);

INVx6_ASAP7_75t_L g13854 ( 
.A(n_13759),
.Y(n_13854)
);

OAI21x1_ASAP7_75t_L g13855 ( 
.A1(n_13348),
.A2(n_12726),
.B(n_12718),
.Y(n_13855)
);

OAI21x1_ASAP7_75t_L g13856 ( 
.A1(n_13338),
.A2(n_12750),
.B(n_12738),
.Y(n_13856)
);

HB1xp67_ASAP7_75t_L g13857 ( 
.A(n_13658),
.Y(n_13857)
);

OAI21x1_ASAP7_75t_L g13858 ( 
.A1(n_13341),
.A2(n_13326),
.B(n_13309),
.Y(n_13858)
);

OAI21xp5_ASAP7_75t_L g13859 ( 
.A1(n_13295),
.A2(n_12809),
.B(n_12807),
.Y(n_13859)
);

NAND2xp5_ASAP7_75t_SL g13860 ( 
.A(n_13649),
.B(n_13011),
.Y(n_13860)
);

NOR2xp33_ASAP7_75t_L g13861 ( 
.A(n_13297),
.B(n_12858),
.Y(n_13861)
);

OAI21x1_ASAP7_75t_L g13862 ( 
.A1(n_13351),
.A2(n_12761),
.B(n_12760),
.Y(n_13862)
);

AOI21x1_ASAP7_75t_L g13863 ( 
.A1(n_13291),
.A2(n_12709),
.B(n_12775),
.Y(n_13863)
);

NAND2x1p5_ASAP7_75t_L g13864 ( 
.A(n_13296),
.B(n_12867),
.Y(n_13864)
);

OR2x6_ASAP7_75t_L g13865 ( 
.A(n_13449),
.B(n_12736),
.Y(n_13865)
);

BUFx2_ASAP7_75t_L g13866 ( 
.A(n_13344),
.Y(n_13866)
);

AO22x2_ASAP7_75t_L g13867 ( 
.A1(n_13451),
.A2(n_13193),
.B1(n_12823),
.B2(n_12840),
.Y(n_13867)
);

OAI22xp5_ASAP7_75t_L g13868 ( 
.A1(n_13426),
.A2(n_12828),
.B1(n_12894),
.B2(n_12784),
.Y(n_13868)
);

AND2x4_ASAP7_75t_L g13869 ( 
.A(n_13741),
.B(n_12950),
.Y(n_13869)
);

OAI21x1_ASAP7_75t_L g13870 ( 
.A1(n_13370),
.A2(n_12824),
.B(n_12817),
.Y(n_13870)
);

NOR2xp33_ASAP7_75t_L g13871 ( 
.A(n_13578),
.B(n_12882),
.Y(n_13871)
);

INVx2_ASAP7_75t_L g13872 ( 
.A(n_13325),
.Y(n_13872)
);

OAI21x1_ASAP7_75t_L g13873 ( 
.A1(n_13317),
.A2(n_12813),
.B(n_12904),
.Y(n_13873)
);

INVx1_ASAP7_75t_L g13874 ( 
.A(n_13307),
.Y(n_13874)
);

OAI21x1_ASAP7_75t_L g13875 ( 
.A1(n_13315),
.A2(n_12704),
.B(n_12690),
.Y(n_13875)
);

INVx3_ASAP7_75t_L g13876 ( 
.A(n_13660),
.Y(n_13876)
);

INVx2_ASAP7_75t_L g13877 ( 
.A(n_13325),
.Y(n_13877)
);

BUFx2_ASAP7_75t_L g13878 ( 
.A(n_13302),
.Y(n_13878)
);

INVx2_ASAP7_75t_SL g13879 ( 
.A(n_13436),
.Y(n_13879)
);

OAI22xp5_ASAP7_75t_L g13880 ( 
.A1(n_13283),
.A2(n_12836),
.B1(n_12844),
.B2(n_12841),
.Y(n_13880)
);

O2A1O1Ixp33_ASAP7_75t_SL g13881 ( 
.A1(n_13705),
.A2(n_12870),
.B(n_12877),
.C(n_12869),
.Y(n_13881)
);

BUFx8_ASAP7_75t_L g13882 ( 
.A(n_13437),
.Y(n_13882)
);

INVx1_ASAP7_75t_L g13883 ( 
.A(n_13312),
.Y(n_13883)
);

INVx1_ASAP7_75t_L g13884 ( 
.A(n_13332),
.Y(n_13884)
);

OAI21x1_ASAP7_75t_SL g13885 ( 
.A1(n_13581),
.A2(n_12822),
.B(n_12878),
.Y(n_13885)
);

INVx2_ASAP7_75t_L g13886 ( 
.A(n_13325),
.Y(n_13886)
);

AND2x2_ASAP7_75t_L g13887 ( 
.A(n_13798),
.B(n_12670),
.Y(n_13887)
);

OAI21x1_ASAP7_75t_L g13888 ( 
.A1(n_13331),
.A2(n_13026),
.B(n_13025),
.Y(n_13888)
);

NOR2xp33_ASAP7_75t_L g13889 ( 
.A(n_13764),
.B(n_12943),
.Y(n_13889)
);

NAND2xp5_ASAP7_75t_L g13890 ( 
.A(n_13506),
.B(n_12612),
.Y(n_13890)
);

OR2x2_ASAP7_75t_L g13891 ( 
.A(n_13350),
.B(n_12939),
.Y(n_13891)
);

NOR2xp33_ASAP7_75t_L g13892 ( 
.A(n_13776),
.B(n_12945),
.Y(n_13892)
);

INVx1_ASAP7_75t_L g13893 ( 
.A(n_13342),
.Y(n_13893)
);

OAI21x1_ASAP7_75t_L g13894 ( 
.A1(n_13310),
.A2(n_13030),
.B(n_13029),
.Y(n_13894)
);

NAND2x1p5_ASAP7_75t_L g13895 ( 
.A(n_13832),
.B(n_12875),
.Y(n_13895)
);

OAI21x1_ASAP7_75t_L g13896 ( 
.A1(n_13284),
.A2(n_13044),
.B(n_13039),
.Y(n_13896)
);

INVx2_ASAP7_75t_L g13897 ( 
.A(n_13325),
.Y(n_13897)
);

OAI21x1_ASAP7_75t_L g13898 ( 
.A1(n_13330),
.A2(n_13383),
.B(n_13314),
.Y(n_13898)
);

INVx1_ASAP7_75t_SL g13899 ( 
.A(n_13688),
.Y(n_13899)
);

NOR2xp67_ASAP7_75t_L g13900 ( 
.A(n_13364),
.B(n_13373),
.Y(n_13900)
);

NAND2xp5_ASAP7_75t_L g13901 ( 
.A(n_13533),
.B(n_13723),
.Y(n_13901)
);

INVx1_ASAP7_75t_L g13902 ( 
.A(n_13354),
.Y(n_13902)
);

AOI21x1_ASAP7_75t_L g13903 ( 
.A1(n_13528),
.A2(n_13061),
.B(n_13051),
.Y(n_13903)
);

AO31x2_ASAP7_75t_L g13904 ( 
.A1(n_13784),
.A2(n_12895),
.A3(n_12891),
.B(n_13065),
.Y(n_13904)
);

INVxp67_ASAP7_75t_SL g13905 ( 
.A(n_13504),
.Y(n_13905)
);

OAI21x1_ASAP7_75t_L g13906 ( 
.A1(n_13793),
.A2(n_13075),
.B(n_13071),
.Y(n_13906)
);

OA21x2_ASAP7_75t_L g13907 ( 
.A1(n_13720),
.A2(n_13081),
.B(n_12959),
.Y(n_13907)
);

AND2x4_ASAP7_75t_L g13908 ( 
.A(n_13327),
.B(n_12640),
.Y(n_13908)
);

AND2x2_ASAP7_75t_L g13909 ( 
.A(n_13401),
.B(n_12637),
.Y(n_13909)
);

INVx1_ASAP7_75t_L g13910 ( 
.A(n_13355),
.Y(n_13910)
);

AND2x2_ASAP7_75t_L g13911 ( 
.A(n_13718),
.B(n_12675),
.Y(n_13911)
);

OAI21x1_ASAP7_75t_SL g13912 ( 
.A1(n_13654),
.A2(n_12973),
.B(n_12957),
.Y(n_13912)
);

AO21x1_ASAP7_75t_L g13913 ( 
.A1(n_13811),
.A2(n_12572),
.B(n_12980),
.Y(n_13913)
);

OAI21x1_ASAP7_75t_L g13914 ( 
.A1(n_13288),
.A2(n_13222),
.B(n_12996),
.Y(n_13914)
);

NAND2xp5_ASAP7_75t_L g13915 ( 
.A(n_13771),
.B(n_12733),
.Y(n_13915)
);

BUFx4f_ASAP7_75t_SL g13916 ( 
.A(n_13531),
.Y(n_13916)
);

BUFx12f_ASAP7_75t_L g13917 ( 
.A(n_13510),
.Y(n_13917)
);

CKINVDCx5p33_ASAP7_75t_R g13918 ( 
.A(n_13457),
.Y(n_13918)
);

NAND2xp5_ASAP7_75t_L g13919 ( 
.A(n_13349),
.B(n_13607),
.Y(n_13919)
);

OAI21x1_ASAP7_75t_L g13920 ( 
.A1(n_13431),
.A2(n_13000),
.B(n_12983),
.Y(n_13920)
);

NOR2xp33_ASAP7_75t_L g13921 ( 
.A(n_13520),
.B(n_13004),
.Y(n_13921)
);

OAI221xp5_ASAP7_75t_L g13922 ( 
.A1(n_13316),
.A2(n_13006),
.B1(n_13017),
.B2(n_13014),
.C(n_13007),
.Y(n_13922)
);

OAI21x1_ASAP7_75t_L g13923 ( 
.A1(n_13432),
.A2(n_13021),
.B(n_13019),
.Y(n_13923)
);

OAI221xp5_ASAP7_75t_L g13924 ( 
.A1(n_13559),
.A2(n_13169),
.B1(n_13180),
.B2(n_13176),
.C(n_13167),
.Y(n_13924)
);

INVx2_ASAP7_75t_L g13925 ( 
.A(n_13399),
.Y(n_13925)
);

INVx1_ASAP7_75t_L g13926 ( 
.A(n_13358),
.Y(n_13926)
);

AND2x4_ASAP7_75t_L g13927 ( 
.A(n_13329),
.B(n_13544),
.Y(n_13927)
);

INVxp67_ASAP7_75t_L g13928 ( 
.A(n_13301),
.Y(n_13928)
);

OAI21x1_ASAP7_75t_L g13929 ( 
.A1(n_13343),
.A2(n_12642),
.B(n_12650),
.Y(n_13929)
);

CKINVDCx5p33_ASAP7_75t_R g13930 ( 
.A(n_13612),
.Y(n_13930)
);

INVx1_ASAP7_75t_L g13931 ( 
.A(n_13366),
.Y(n_13931)
);

BUFx3_ASAP7_75t_L g13932 ( 
.A(n_13402),
.Y(n_13932)
);

INVx3_ASAP7_75t_L g13933 ( 
.A(n_13574),
.Y(n_13933)
);

AND2x2_ASAP7_75t_L g13934 ( 
.A(n_13651),
.B(n_12776),
.Y(n_13934)
);

NOR2xp33_ASAP7_75t_L g13935 ( 
.A(n_13584),
.B(n_13134),
.Y(n_13935)
);

BUFx8_ASAP7_75t_L g13936 ( 
.A(n_13518),
.Y(n_13936)
);

INVx1_ASAP7_75t_L g13937 ( 
.A(n_13369),
.Y(n_13937)
);

OAI21x1_ASAP7_75t_SL g13938 ( 
.A1(n_13717),
.A2(n_12734),
.B(n_12721),
.Y(n_13938)
);

OAI21x1_ASAP7_75t_L g13939 ( 
.A1(n_13697),
.A2(n_12749),
.B(n_12732),
.Y(n_13939)
);

INVx1_ASAP7_75t_L g13940 ( 
.A(n_13404),
.Y(n_13940)
);

CKINVDCx5p33_ASAP7_75t_R g13941 ( 
.A(n_13357),
.Y(n_13941)
);

BUFx2_ASAP7_75t_L g13942 ( 
.A(n_13333),
.Y(n_13942)
);

INVx2_ASAP7_75t_SL g13943 ( 
.A(n_13526),
.Y(n_13943)
);

OAI21xp5_ASAP7_75t_L g13944 ( 
.A1(n_13362),
.A2(n_13042),
.B(n_13140),
.Y(n_13944)
);

BUFx2_ASAP7_75t_L g13945 ( 
.A(n_13652),
.Y(n_13945)
);

AO31x2_ASAP7_75t_L g13946 ( 
.A1(n_13820),
.A2(n_13248),
.A3(n_13100),
.B(n_12686),
.Y(n_13946)
);

INVx1_ASAP7_75t_L g13947 ( 
.A(n_13430),
.Y(n_13947)
);

AND2x4_ASAP7_75t_L g13948 ( 
.A(n_13768),
.B(n_12954),
.Y(n_13948)
);

INVx1_ASAP7_75t_L g13949 ( 
.A(n_13445),
.Y(n_13949)
);

AOI22xp33_ASAP7_75t_L g13950 ( 
.A1(n_13318),
.A2(n_13193),
.B1(n_13149),
.B2(n_13018),
.Y(n_13950)
);

NAND2x1p5_ASAP7_75t_L g13951 ( 
.A(n_13689),
.B(n_12919),
.Y(n_13951)
);

AOI21x1_ASAP7_75t_L g13952 ( 
.A1(n_13616),
.A2(n_12764),
.B(n_12763),
.Y(n_13952)
);

AO21x2_ASAP7_75t_L g13953 ( 
.A1(n_13406),
.A2(n_13118),
.B(n_12949),
.Y(n_13953)
);

BUFx6f_ASAP7_75t_L g13954 ( 
.A(n_13412),
.Y(n_13954)
);

NAND2x1p5_ASAP7_75t_L g13955 ( 
.A(n_13551),
.B(n_12648),
.Y(n_13955)
);

BUFx3_ASAP7_75t_L g13956 ( 
.A(n_13503),
.Y(n_13956)
);

INVx2_ASAP7_75t_L g13957 ( 
.A(n_13400),
.Y(n_13957)
);

OAI21xp5_ASAP7_75t_L g13958 ( 
.A1(n_13372),
.A2(n_13028),
.B(n_13024),
.Y(n_13958)
);

INVx2_ASAP7_75t_L g13959 ( 
.A(n_13458),
.Y(n_13959)
);

INVx1_ASAP7_75t_L g13960 ( 
.A(n_13448),
.Y(n_13960)
);

INVx2_ASAP7_75t_L g13961 ( 
.A(n_13507),
.Y(n_13961)
);

AO21x2_ASAP7_75t_L g13962 ( 
.A1(n_13420),
.A2(n_12929),
.B(n_12765),
.Y(n_13962)
);

AOI222xp33_ASAP7_75t_L g13963 ( 
.A1(n_13443),
.A2(n_13676),
.B1(n_13700),
.B2(n_13637),
.C1(n_13682),
.C2(n_13363),
.Y(n_13963)
);

BUFx12f_ASAP7_75t_L g13964 ( 
.A(n_13495),
.Y(n_13964)
);

NOR2xp33_ASAP7_75t_L g13965 ( 
.A(n_13511),
.B(n_12888),
.Y(n_13965)
);

OAI21x1_ASAP7_75t_L g13966 ( 
.A1(n_13643),
.A2(n_12898),
.B(n_12889),
.Y(n_13966)
);

OR2x2_ASAP7_75t_L g13967 ( 
.A(n_13732),
.B(n_13743),
.Y(n_13967)
);

NAND2xp5_ASAP7_75t_SL g13968 ( 
.A(n_13294),
.B(n_13045),
.Y(n_13968)
);

AND2x4_ASAP7_75t_L g13969 ( 
.A(n_13819),
.B(n_12926),
.Y(n_13969)
);

AOI22xp33_ASAP7_75t_L g13970 ( 
.A1(n_13339),
.A2(n_13062),
.B1(n_12961),
.B2(n_12977),
.Y(n_13970)
);

INVx2_ASAP7_75t_L g13971 ( 
.A(n_13286),
.Y(n_13971)
);

INVx2_ASAP7_75t_L g13972 ( 
.A(n_13361),
.Y(n_13972)
);

INVx5_ASAP7_75t_L g13973 ( 
.A(n_13440),
.Y(n_13973)
);

NOR2xp33_ASAP7_75t_R g13974 ( 
.A(n_13745),
.B(n_12884),
.Y(n_13974)
);

AOI22xp33_ASAP7_75t_L g13975 ( 
.A1(n_13429),
.A2(n_12992),
.B1(n_13003),
.B2(n_12928),
.Y(n_13975)
);

NAND2xp5_ASAP7_75t_L g13976 ( 
.A(n_13661),
.B(n_12781),
.Y(n_13976)
);

INVx6_ASAP7_75t_L g13977 ( 
.A(n_13747),
.Y(n_13977)
);

OAI21x1_ASAP7_75t_L g13978 ( 
.A1(n_13662),
.A2(n_12795),
.B(n_12799),
.Y(n_13978)
);

OR2x2_ASAP7_75t_L g13979 ( 
.A(n_13461),
.B(n_12815),
.Y(n_13979)
);

NAND2xp5_ASAP7_75t_L g13980 ( 
.A(n_13672),
.B(n_13677),
.Y(n_13980)
);

OA21x2_ASAP7_75t_L g13981 ( 
.A1(n_13456),
.A2(n_12868),
.B(n_12863),
.Y(n_13981)
);

NAND2xp5_ASAP7_75t_L g13982 ( 
.A(n_13694),
.B(n_12847),
.Y(n_13982)
);

INVx2_ASAP7_75t_L g13983 ( 
.A(n_13378),
.Y(n_13983)
);

INVx2_ASAP7_75t_L g13984 ( 
.A(n_13388),
.Y(n_13984)
);

OAI21x1_ASAP7_75t_L g13985 ( 
.A1(n_13696),
.A2(n_12545),
.B(n_13040),
.Y(n_13985)
);

OA21x2_ASAP7_75t_L g13986 ( 
.A1(n_13460),
.A2(n_12912),
.B(n_12991),
.Y(n_13986)
);

INVx6_ASAP7_75t_L g13987 ( 
.A(n_13757),
.Y(n_13987)
);

CKINVDCx11_ASAP7_75t_R g13988 ( 
.A(n_13833),
.Y(n_13988)
);

BUFx3_ASAP7_75t_L g13989 ( 
.A(n_13656),
.Y(n_13989)
);

INVx1_ASAP7_75t_L g13990 ( 
.A(n_13468),
.Y(n_13990)
);

OR2x2_ASAP7_75t_L g13991 ( 
.A(n_13569),
.B(n_1912),
.Y(n_13991)
);

OA21x2_ASAP7_75t_L g13992 ( 
.A1(n_13603),
.A2(n_12855),
.B(n_12792),
.Y(n_13992)
);

BUFx6f_ASAP7_75t_L g13993 ( 
.A(n_13322),
.Y(n_13993)
);

AOI21x1_ASAP7_75t_L g13994 ( 
.A1(n_13591),
.A2(n_13023),
.B(n_12896),
.Y(n_13994)
);

INVx1_ASAP7_75t_L g13995 ( 
.A(n_13474),
.Y(n_13995)
);

INVx2_ASAP7_75t_L g13996 ( 
.A(n_13394),
.Y(n_13996)
);

OAI22xp5_ASAP7_75t_L g13997 ( 
.A1(n_13335),
.A2(n_13605),
.B1(n_13359),
.B2(n_13738),
.Y(n_13997)
);

AOI21x1_ASAP7_75t_L g13998 ( 
.A1(n_13415),
.A2(n_13227),
.B(n_1913),
.Y(n_13998)
);

INVx1_ASAP7_75t_L g13999 ( 
.A(n_13477),
.Y(n_13999)
);

NAND2xp5_ASAP7_75t_L g14000 ( 
.A(n_13345),
.B(n_1913),
.Y(n_14000)
);

INVx1_ASAP7_75t_L g14001 ( 
.A(n_13494),
.Y(n_14001)
);

INVx2_ASAP7_75t_L g14002 ( 
.A(n_13395),
.Y(n_14002)
);

INVx1_ASAP7_75t_L g14003 ( 
.A(n_13499),
.Y(n_14003)
);

NAND2xp5_ASAP7_75t_L g14004 ( 
.A(n_13617),
.B(n_13838),
.Y(n_14004)
);

OAI21xp5_ASAP7_75t_L g14005 ( 
.A1(n_13356),
.A2(n_13347),
.B(n_13550),
.Y(n_14005)
);

HB1xp67_ASAP7_75t_L g14006 ( 
.A(n_13519),
.Y(n_14006)
);

NAND2x1p5_ASAP7_75t_L g14007 ( 
.A(n_13352),
.B(n_1914),
.Y(n_14007)
);

NAND2xp5_ASAP7_75t_L g14008 ( 
.A(n_13285),
.B(n_1915),
.Y(n_14008)
);

AO21x2_ASAP7_75t_L g14009 ( 
.A1(n_13834),
.A2(n_13827),
.B(n_13704),
.Y(n_14009)
);

INVx1_ASAP7_75t_L g14010 ( 
.A(n_13543),
.Y(n_14010)
);

AND2x2_ASAP7_75t_L g14011 ( 
.A(n_13713),
.B(n_1915),
.Y(n_14011)
);

OA21x2_ASAP7_75t_L g14012 ( 
.A1(n_13802),
.A2(n_1916),
.B(n_1917),
.Y(n_14012)
);

CKINVDCx20_ASAP7_75t_R g14013 ( 
.A(n_13758),
.Y(n_14013)
);

INVx1_ASAP7_75t_L g14014 ( 
.A(n_13572),
.Y(n_14014)
);

INVx2_ASAP7_75t_L g14015 ( 
.A(n_13340),
.Y(n_14015)
);

INVx6_ASAP7_75t_L g14016 ( 
.A(n_13805),
.Y(n_14016)
);

OA21x2_ASAP7_75t_L g14017 ( 
.A1(n_13580),
.A2(n_1918),
.B(n_1919),
.Y(n_14017)
);

INVx1_ASAP7_75t_L g14018 ( 
.A(n_13594),
.Y(n_14018)
);

INVx2_ASAP7_75t_L g14019 ( 
.A(n_13353),
.Y(n_14019)
);

OA21x2_ASAP7_75t_L g14020 ( 
.A1(n_13597),
.A2(n_1918),
.B(n_1919),
.Y(n_14020)
);

OAI21x1_ASAP7_75t_L g14021 ( 
.A1(n_13532),
.A2(n_1920),
.B(n_1921),
.Y(n_14021)
);

AND2x4_ASAP7_75t_L g14022 ( 
.A(n_13292),
.B(n_1920),
.Y(n_14022)
);

AOI22xp33_ASAP7_75t_L g14023 ( 
.A1(n_13299),
.A2(n_1923),
.B1(n_1921),
.B2(n_1922),
.Y(n_14023)
);

OA21x2_ASAP7_75t_L g14024 ( 
.A1(n_13571),
.A2(n_13537),
.B(n_13638),
.Y(n_14024)
);

NAND2xp5_ASAP7_75t_L g14025 ( 
.A(n_13734),
.B(n_13744),
.Y(n_14025)
);

AOI21x1_ASAP7_75t_L g14026 ( 
.A1(n_13482),
.A2(n_1922),
.B(n_1923),
.Y(n_14026)
);

AOI22xp33_ASAP7_75t_L g14027 ( 
.A1(n_13481),
.A2(n_13483),
.B1(n_13320),
.B2(n_13298),
.Y(n_14027)
);

NOR2xp33_ASAP7_75t_L g14028 ( 
.A(n_13475),
.B(n_1924),
.Y(n_14028)
);

INVx1_ASAP7_75t_L g14029 ( 
.A(n_13668),
.Y(n_14029)
);

INVx3_ASAP7_75t_L g14030 ( 
.A(n_13322),
.Y(n_14030)
);

OA21x2_ASAP7_75t_L g14031 ( 
.A1(n_13760),
.A2(n_1925),
.B(n_1926),
.Y(n_14031)
);

O2A1O1Ixp33_ASAP7_75t_L g14032 ( 
.A1(n_13321),
.A2(n_1927),
.B(n_1925),
.C(n_1926),
.Y(n_14032)
);

O2A1O1Ixp33_ASAP7_75t_L g14033 ( 
.A1(n_13416),
.A2(n_13396),
.B(n_13587),
.C(n_13485),
.Y(n_14033)
);

OAI21x1_ASAP7_75t_L g14034 ( 
.A1(n_13513),
.A2(n_1928),
.B(n_1929),
.Y(n_14034)
);

INVx1_ASAP7_75t_L g14035 ( 
.A(n_13804),
.Y(n_14035)
);

CKINVDCx5p33_ASAP7_75t_R g14036 ( 
.A(n_13796),
.Y(n_14036)
);

OAI21x1_ASAP7_75t_L g14037 ( 
.A1(n_13514),
.A2(n_1928),
.B(n_1929),
.Y(n_14037)
);

O2A1O1Ixp33_ASAP7_75t_SL g14038 ( 
.A1(n_13376),
.A2(n_1932),
.B(n_1930),
.C(n_1931),
.Y(n_14038)
);

OAI21x1_ASAP7_75t_L g14039 ( 
.A1(n_13368),
.A2(n_1931),
.B(n_1932),
.Y(n_14039)
);

A2O1A1Ixp33_ASAP7_75t_L g14040 ( 
.A1(n_13442),
.A2(n_1935),
.B(n_1933),
.C(n_1934),
.Y(n_14040)
);

INVx1_ASAP7_75t_SL g14041 ( 
.A(n_13773),
.Y(n_14041)
);

INVx2_ASAP7_75t_L g14042 ( 
.A(n_13525),
.Y(n_14042)
);

OR3x4_ASAP7_75t_SL g14043 ( 
.A(n_13629),
.B(n_1934),
.C(n_1935),
.Y(n_14043)
);

AND2x2_ASAP7_75t_L g14044 ( 
.A(n_13810),
.B(n_1936),
.Y(n_14044)
);

HB1xp67_ASAP7_75t_L g14045 ( 
.A(n_13816),
.Y(n_14045)
);

HB1xp67_ASAP7_75t_L g14046 ( 
.A(n_13684),
.Y(n_14046)
);

OR2x2_ASAP7_75t_L g14047 ( 
.A(n_13592),
.B(n_1936),
.Y(n_14047)
);

NAND2x1p5_ASAP7_75t_L g14048 ( 
.A(n_13308),
.B(n_1937),
.Y(n_14048)
);

OAI21x1_ASAP7_75t_L g14049 ( 
.A1(n_13418),
.A2(n_13493),
.B(n_13410),
.Y(n_14049)
);

INVx1_ASAP7_75t_L g14050 ( 
.A(n_13427),
.Y(n_14050)
);

AND2x2_ASAP7_75t_L g14051 ( 
.A(n_13487),
.B(n_1938),
.Y(n_14051)
);

AOI22xp33_ASAP7_75t_L g14052 ( 
.A1(n_13439),
.A2(n_1940),
.B1(n_1938),
.B2(n_1939),
.Y(n_14052)
);

AO21x2_ASAP7_75t_L g14053 ( 
.A1(n_13471),
.A2(n_1940),
.B(n_1941),
.Y(n_14053)
);

CKINVDCx5p33_ASAP7_75t_R g14054 ( 
.A(n_13538),
.Y(n_14054)
);

OAI21x1_ASAP7_75t_L g14055 ( 
.A1(n_13498),
.A2(n_1941),
.B(n_1942),
.Y(n_14055)
);

O2A1O1Ixp33_ASAP7_75t_SL g14056 ( 
.A1(n_13624),
.A2(n_1945),
.B(n_1943),
.C(n_1944),
.Y(n_14056)
);

OAI21xp5_ASAP7_75t_L g14057 ( 
.A1(n_13450),
.A2(n_1943),
.B(n_1945),
.Y(n_14057)
);

INVx1_ASAP7_75t_SL g14058 ( 
.A(n_13707),
.Y(n_14058)
);

INVx2_ASAP7_75t_L g14059 ( 
.A(n_13797),
.Y(n_14059)
);

INVx8_ASAP7_75t_L g14060 ( 
.A(n_13440),
.Y(n_14060)
);

AO21x2_ASAP7_75t_L g14061 ( 
.A1(n_13491),
.A2(n_1947),
.B(n_1948),
.Y(n_14061)
);

OAI21xp5_ASAP7_75t_L g14062 ( 
.A1(n_13497),
.A2(n_1947),
.B(n_1948),
.Y(n_14062)
);

NOR2xp33_ASAP7_75t_L g14063 ( 
.A(n_13446),
.B(n_1949),
.Y(n_14063)
);

CKINVDCx11_ASAP7_75t_R g14064 ( 
.A(n_13833),
.Y(n_14064)
);

OA21x2_ASAP7_75t_L g14065 ( 
.A1(n_13529),
.A2(n_1949),
.B(n_1950),
.Y(n_14065)
);

NOR2xp33_ASAP7_75t_L g14066 ( 
.A(n_13336),
.B(n_1950),
.Y(n_14066)
);

AND2x2_ASAP7_75t_L g14067 ( 
.A(n_13300),
.B(n_1951),
.Y(n_14067)
);

INVx1_ASAP7_75t_L g14068 ( 
.A(n_13409),
.Y(n_14068)
);

OAI21x1_ASAP7_75t_L g14069 ( 
.A1(n_13385),
.A2(n_1951),
.B(n_1952),
.Y(n_14069)
);

INVx1_ASAP7_75t_L g14070 ( 
.A(n_13409),
.Y(n_14070)
);

OAI222xp33_ASAP7_75t_L g14071 ( 
.A1(n_13585),
.A2(n_1954),
.B1(n_1956),
.B2(n_1952),
.C1(n_1953),
.C2(n_1955),
.Y(n_14071)
);

INVx2_ASAP7_75t_L g14072 ( 
.A(n_13800),
.Y(n_14072)
);

OAI221xp5_ASAP7_75t_L g14073 ( 
.A1(n_13678),
.A2(n_1955),
.B1(n_1953),
.B2(n_1954),
.C(n_1956),
.Y(n_14073)
);

AOI21x1_ASAP7_75t_L g14074 ( 
.A1(n_13675),
.A2(n_1957),
.B(n_1958),
.Y(n_14074)
);

AND2x4_ASAP7_75t_L g14075 ( 
.A(n_13290),
.B(n_1957),
.Y(n_14075)
);

AOI22xp33_ASAP7_75t_L g14076 ( 
.A1(n_13602),
.A2(n_1960),
.B1(n_1958),
.B2(n_1959),
.Y(n_14076)
);

OAI21x1_ASAP7_75t_L g14077 ( 
.A1(n_13545),
.A2(n_1959),
.B(n_1960),
.Y(n_14077)
);

INVx1_ASAP7_75t_SL g14078 ( 
.A(n_13835),
.Y(n_14078)
);

NAND2xp5_ASAP7_75t_L g14079 ( 
.A(n_13535),
.B(n_1961),
.Y(n_14079)
);

OAI22xp5_ASAP7_75t_L g14080 ( 
.A1(n_13588),
.A2(n_1964),
.B1(n_1962),
.B2(n_1963),
.Y(n_14080)
);

HB1xp67_ASAP7_75t_L g14081 ( 
.A(n_13693),
.Y(n_14081)
);

INVx2_ASAP7_75t_L g14082 ( 
.A(n_13724),
.Y(n_14082)
);

OAI21x1_ASAP7_75t_L g14083 ( 
.A1(n_13547),
.A2(n_1964),
.B(n_1965),
.Y(n_14083)
);

AOI21x1_ASAP7_75t_L g14084 ( 
.A1(n_13548),
.A2(n_1966),
.B(n_1967),
.Y(n_14084)
);

INVx1_ASAP7_75t_L g14085 ( 
.A(n_13463),
.Y(n_14085)
);

OAI21x1_ASAP7_75t_L g14086 ( 
.A1(n_13382),
.A2(n_1966),
.B(n_1967),
.Y(n_14086)
);

OAI22xp33_ASAP7_75t_L g14087 ( 
.A1(n_13304),
.A2(n_1970),
.B1(n_1968),
.B2(n_1969),
.Y(n_14087)
);

AOI22xp33_ASAP7_75t_L g14088 ( 
.A1(n_13328),
.A2(n_1971),
.B1(n_1968),
.B2(n_1970),
.Y(n_14088)
);

OAI21x1_ASAP7_75t_L g14089 ( 
.A1(n_13462),
.A2(n_13623),
.B(n_13397),
.Y(n_14089)
);

NAND3xp33_ASAP7_75t_L g14090 ( 
.A(n_13377),
.B(n_1971),
.C(n_1972),
.Y(n_14090)
);

INVxp67_ASAP7_75t_L g14091 ( 
.A(n_13814),
.Y(n_14091)
);

AOI21xp5_ASAP7_75t_L g14092 ( 
.A1(n_13303),
.A2(n_1972),
.B(n_1973),
.Y(n_14092)
);

BUFx3_ASAP7_75t_L g14093 ( 
.A(n_13806),
.Y(n_14093)
);

OAI22xp5_ASAP7_75t_L g14094 ( 
.A1(n_13601),
.A2(n_1975),
.B1(n_1973),
.B2(n_1974),
.Y(n_14094)
);

OAI21x1_ASAP7_75t_L g14095 ( 
.A1(n_13398),
.A2(n_1974),
.B(n_1976),
.Y(n_14095)
);

HB1xp67_ASAP7_75t_L g14096 ( 
.A(n_13568),
.Y(n_14096)
);

AOI21xp5_ASAP7_75t_L g14097 ( 
.A1(n_13319),
.A2(n_1977),
.B(n_1980),
.Y(n_14097)
);

BUFx2_ASAP7_75t_SL g14098 ( 
.A(n_13753),
.Y(n_14098)
);

NOR2xp67_ASAP7_75t_L g14099 ( 
.A(n_13788),
.B(n_13818),
.Y(n_14099)
);

NOR2xp67_ASAP7_75t_L g14100 ( 
.A(n_13727),
.B(n_1980),
.Y(n_14100)
);

NAND2xp5_ASAP7_75t_L g14101 ( 
.A(n_13530),
.B(n_1981),
.Y(n_14101)
);

BUFx2_ASAP7_75t_L g14102 ( 
.A(n_13825),
.Y(n_14102)
);

INVx2_ASAP7_75t_L g14103 ( 
.A(n_13828),
.Y(n_14103)
);

OAI21x1_ASAP7_75t_L g14104 ( 
.A1(n_13523),
.A2(n_13645),
.B(n_13627),
.Y(n_14104)
);

OAI21x1_ASAP7_75t_SL g14105 ( 
.A1(n_13736),
.A2(n_1981),
.B(n_1982),
.Y(n_14105)
);

OA21x2_ASAP7_75t_L g14106 ( 
.A1(n_13554),
.A2(n_1982),
.B(n_1983),
.Y(n_14106)
);

OAI21x1_ASAP7_75t_SL g14107 ( 
.A1(n_13775),
.A2(n_13639),
.B(n_13777),
.Y(n_14107)
);

AND2x4_ASAP7_75t_L g14108 ( 
.A(n_13831),
.B(n_1983),
.Y(n_14108)
);

OAI21x1_ASAP7_75t_L g14109 ( 
.A1(n_13750),
.A2(n_1984),
.B(n_1985),
.Y(n_14109)
);

OAI22xp5_ASAP7_75t_L g14110 ( 
.A1(n_13407),
.A2(n_1986),
.B1(n_1984),
.B2(n_1985),
.Y(n_14110)
);

NAND2xp5_ASAP7_75t_L g14111 ( 
.A(n_13752),
.B(n_1986),
.Y(n_14111)
);

INVxp67_ASAP7_75t_L g14112 ( 
.A(n_13725),
.Y(n_14112)
);

AOI22x1_ASAP7_75t_L g14113 ( 
.A1(n_13536),
.A2(n_1989),
.B1(n_1987),
.B2(n_1988),
.Y(n_14113)
);

BUFx6f_ASAP7_75t_L g14114 ( 
.A(n_13360),
.Y(n_14114)
);

CKINVDCx8_ASAP7_75t_R g14115 ( 
.A(n_13767),
.Y(n_14115)
);

NAND2xp5_ASAP7_75t_L g14116 ( 
.A(n_13735),
.B(n_1988),
.Y(n_14116)
);

BUFx3_ASAP7_75t_L g14117 ( 
.A(n_13737),
.Y(n_14117)
);

NOR2xp67_ASAP7_75t_SL g14118 ( 
.A(n_13473),
.B(n_1989),
.Y(n_14118)
);

BUFx8_ASAP7_75t_SL g14119 ( 
.A(n_13549),
.Y(n_14119)
);

AOI22xp5_ASAP7_75t_L g14120 ( 
.A1(n_13722),
.A2(n_1992),
.B1(n_1990),
.B2(n_1991),
.Y(n_14120)
);

BUFx6f_ASAP7_75t_L g14121 ( 
.A(n_13360),
.Y(n_14121)
);

AO21x2_ASAP7_75t_L g14122 ( 
.A1(n_13556),
.A2(n_1990),
.B(n_1991),
.Y(n_14122)
);

AOI22xp33_ASAP7_75t_L g14123 ( 
.A1(n_13575),
.A2(n_1994),
.B1(n_1992),
.B2(n_1993),
.Y(n_14123)
);

INVx2_ASAP7_75t_L g14124 ( 
.A(n_13608),
.Y(n_14124)
);

AO21x2_ASAP7_75t_L g14125 ( 
.A1(n_13582),
.A2(n_1993),
.B(n_1994),
.Y(n_14125)
);

AND2x2_ASAP7_75t_L g14126 ( 
.A(n_13679),
.B(n_1995),
.Y(n_14126)
);

OAI21x1_ASAP7_75t_L g14127 ( 
.A1(n_13761),
.A2(n_1995),
.B(n_1996),
.Y(n_14127)
);

NAND2xp5_ASAP7_75t_L g14128 ( 
.A(n_13472),
.B(n_1996),
.Y(n_14128)
);

OAI21x1_ASAP7_75t_L g14129 ( 
.A1(n_13782),
.A2(n_1997),
.B(n_1998),
.Y(n_14129)
);

OAI21x1_ASAP7_75t_L g14130 ( 
.A1(n_13815),
.A2(n_1997),
.B(n_1998),
.Y(n_14130)
);

AO21x2_ASAP7_75t_L g14131 ( 
.A1(n_13598),
.A2(n_1999),
.B(n_2000),
.Y(n_14131)
);

OA21x2_ASAP7_75t_L g14132 ( 
.A1(n_13749),
.A2(n_2001),
.B(n_2002),
.Y(n_14132)
);

OAI21xp33_ASAP7_75t_SL g14133 ( 
.A1(n_13496),
.A2(n_2001),
.B(n_2002),
.Y(n_14133)
);

INVxp67_ASAP7_75t_SL g14134 ( 
.A(n_13425),
.Y(n_14134)
);

AO21x1_ASAP7_75t_L g14135 ( 
.A1(n_13786),
.A2(n_2003),
.B(n_2004),
.Y(n_14135)
);

CKINVDCx5p33_ASAP7_75t_R g14136 ( 
.A(n_13381),
.Y(n_14136)
);

OAI21xp5_ASAP7_75t_L g14137 ( 
.A1(n_13555),
.A2(n_13615),
.B(n_13567),
.Y(n_14137)
);

INVx2_ASAP7_75t_L g14138 ( 
.A(n_13765),
.Y(n_14138)
);

OAI21x1_ASAP7_75t_L g14139 ( 
.A1(n_13625),
.A2(n_2003),
.B(n_2004),
.Y(n_14139)
);

BUFx2_ASAP7_75t_L g14140 ( 
.A(n_13381),
.Y(n_14140)
);

OAI21x1_ASAP7_75t_L g14141 ( 
.A1(n_13626),
.A2(n_2005),
.B(n_2006),
.Y(n_14141)
);

INVx1_ASAP7_75t_L g14142 ( 
.A(n_13463),
.Y(n_14142)
);

XNOR2xp5_ASAP7_75t_L g14143 ( 
.A(n_13779),
.B(n_2005),
.Y(n_14143)
);

OAI21x1_ASAP7_75t_L g14144 ( 
.A1(n_13653),
.A2(n_2007),
.B(n_2008),
.Y(n_14144)
);

BUFx2_ASAP7_75t_L g14145 ( 
.A(n_13478),
.Y(n_14145)
);

NAND2xp5_ASAP7_75t_L g14146 ( 
.A(n_13512),
.B(n_2007),
.Y(n_14146)
);

NAND2x1p5_ASAP7_75t_L g14147 ( 
.A(n_13642),
.B(n_2008),
.Y(n_14147)
);

OAI21x1_ASAP7_75t_L g14148 ( 
.A1(n_13657),
.A2(n_2009),
.B(n_2010),
.Y(n_14148)
);

OAI21x1_ASAP7_75t_L g14149 ( 
.A1(n_13671),
.A2(n_2009),
.B(n_2010),
.Y(n_14149)
);

A2O1A1Ixp33_ASAP7_75t_L g14150 ( 
.A1(n_13419),
.A2(n_2013),
.B(n_2011),
.C(n_2012),
.Y(n_14150)
);

OA21x2_ASAP7_75t_L g14151 ( 
.A1(n_13611),
.A2(n_13673),
.B(n_13663),
.Y(n_14151)
);

AO31x2_ASAP7_75t_L g14152 ( 
.A1(n_13454),
.A2(n_2015),
.A3(n_2012),
.B(n_2014),
.Y(n_14152)
);

AOI22xp33_ASAP7_75t_L g14153 ( 
.A1(n_13387),
.A2(n_2017),
.B1(n_2015),
.B2(n_2016),
.Y(n_14153)
);

OAI21x1_ASAP7_75t_L g14154 ( 
.A1(n_13680),
.A2(n_2016),
.B(n_2017),
.Y(n_14154)
);

BUFx3_ASAP7_75t_L g14155 ( 
.A(n_13737),
.Y(n_14155)
);

NAND2xp5_ASAP7_75t_L g14156 ( 
.A(n_13539),
.B(n_2019),
.Y(n_14156)
);

AND2x2_ASAP7_75t_L g14157 ( 
.A(n_13478),
.B(n_2020),
.Y(n_14157)
);

OAI21x1_ASAP7_75t_L g14158 ( 
.A1(n_13563),
.A2(n_2020),
.B(n_2021),
.Y(n_14158)
);

OAI22xp5_ASAP7_75t_L g14159 ( 
.A1(n_13795),
.A2(n_2023),
.B1(n_2021),
.B2(n_2022),
.Y(n_14159)
);

INVx2_ASAP7_75t_L g14160 ( 
.A(n_13480),
.Y(n_14160)
);

AND2x4_ASAP7_75t_L g14161 ( 
.A(n_13599),
.B(n_2022),
.Y(n_14161)
);

CKINVDCx20_ASAP7_75t_R g14162 ( 
.A(n_13767),
.Y(n_14162)
);

INVx1_ASAP7_75t_L g14163 ( 
.A(n_13480),
.Y(n_14163)
);

AND2x2_ASAP7_75t_L g14164 ( 
.A(n_13599),
.B(n_2023),
.Y(n_14164)
);

BUFx3_ASAP7_75t_L g14165 ( 
.A(n_13614),
.Y(n_14165)
);

AND2x2_ASAP7_75t_L g14166 ( 
.A(n_13614),
.B(n_2024),
.Y(n_14166)
);

OA21x2_ASAP7_75t_L g14167 ( 
.A1(n_13683),
.A2(n_2024),
.B(n_2025),
.Y(n_14167)
);

OA21x2_ASAP7_75t_L g14168 ( 
.A1(n_13428),
.A2(n_2025),
.B(n_2026),
.Y(n_14168)
);

INVx1_ASAP7_75t_L g14169 ( 
.A(n_13509),
.Y(n_14169)
);

OAI21x1_ASAP7_75t_L g14170 ( 
.A1(n_13374),
.A2(n_2026),
.B(n_2027),
.Y(n_14170)
);

INVx1_ASAP7_75t_L g14171 ( 
.A(n_13509),
.Y(n_14171)
);

INVx2_ASAP7_75t_L g14172 ( 
.A(n_13565),
.Y(n_14172)
);

OAI21x1_ASAP7_75t_L g14173 ( 
.A1(n_13783),
.A2(n_13380),
.B(n_13433),
.Y(n_14173)
);

OAI21x1_ASAP7_75t_L g14174 ( 
.A1(n_13435),
.A2(n_2027),
.B(n_2028),
.Y(n_14174)
);

OAI21xp5_ASAP7_75t_L g14175 ( 
.A1(n_13619),
.A2(n_2028),
.B(n_2029),
.Y(n_14175)
);

OAI21x1_ASAP7_75t_SL g14176 ( 
.A1(n_13836),
.A2(n_2029),
.B(n_2030),
.Y(n_14176)
);

INVx3_ASAP7_75t_L g14177 ( 
.A(n_13635),
.Y(n_14177)
);

OAI21x1_ASAP7_75t_L g14178 ( 
.A1(n_13438),
.A2(n_2031),
.B(n_2032),
.Y(n_14178)
);

OAI21x1_ASAP7_75t_L g14179 ( 
.A1(n_13444),
.A2(n_2031),
.B(n_2032),
.Y(n_14179)
);

AOI22xp5_ASAP7_75t_L g14180 ( 
.A1(n_13809),
.A2(n_2035),
.B1(n_2033),
.B2(n_2034),
.Y(n_14180)
);

BUFx3_ASAP7_75t_L g14181 ( 
.A(n_13635),
.Y(n_14181)
);

NAND2x1p5_ASAP7_75t_L g14182 ( 
.A(n_13486),
.B(n_2033),
.Y(n_14182)
);

NAND2xp5_ASAP7_75t_L g14183 ( 
.A(n_13593),
.B(n_2034),
.Y(n_14183)
);

INVx1_ASAP7_75t_L g14184 ( 
.A(n_13540),
.Y(n_14184)
);

OAI22xp33_ASAP7_75t_L g14185 ( 
.A1(n_13586),
.A2(n_13346),
.B1(n_13579),
.B2(n_13664),
.Y(n_14185)
);

OAI21x1_ASAP7_75t_L g14186 ( 
.A1(n_13447),
.A2(n_2035),
.B(n_2036),
.Y(n_14186)
);

OAI21x1_ASAP7_75t_L g14187 ( 
.A1(n_13467),
.A2(n_2036),
.B(n_2037),
.Y(n_14187)
);

CKINVDCx5p33_ASAP7_75t_R g14188 ( 
.A(n_13690),
.Y(n_14188)
);

AOI21xp5_ASAP7_75t_L g14189 ( 
.A1(n_13516),
.A2(n_2037),
.B(n_2038),
.Y(n_14189)
);

AOI22xp33_ASAP7_75t_L g14190 ( 
.A1(n_13609),
.A2(n_2041),
.B1(n_2039),
.B2(n_2040),
.Y(n_14190)
);

AND2x4_ASAP7_75t_L g14191 ( 
.A(n_13690),
.B(n_2039),
.Y(n_14191)
);

INVx3_ASAP7_75t_L g14192 ( 
.A(n_13470),
.Y(n_14192)
);

OAI22xp5_ASAP7_75t_L g14193 ( 
.A1(n_13453),
.A2(n_2042),
.B1(n_2040),
.B2(n_2041),
.Y(n_14193)
);

HB1xp67_ASAP7_75t_L g14194 ( 
.A(n_13334),
.Y(n_14194)
);

O2A1O1Ixp33_ASAP7_75t_SL g14195 ( 
.A1(n_13792),
.A2(n_2044),
.B(n_2042),
.C(n_2043),
.Y(n_14195)
);

OAI21x1_ASAP7_75t_L g14196 ( 
.A1(n_13570),
.A2(n_13577),
.B(n_13564),
.Y(n_14196)
);

NOR2xp33_ASAP7_75t_L g14197 ( 
.A(n_13823),
.B(n_2043),
.Y(n_14197)
);

NAND2xp5_ASAP7_75t_L g14198 ( 
.A(n_13408),
.B(n_13630),
.Y(n_14198)
);

AOI21xp5_ASAP7_75t_L g14199 ( 
.A1(n_13517),
.A2(n_2044),
.B(n_2045),
.Y(n_14199)
);

NAND2xp5_ASAP7_75t_L g14200 ( 
.A(n_13681),
.B(n_2045),
.Y(n_14200)
);

INVx2_ASAP7_75t_SL g14201 ( 
.A(n_13393),
.Y(n_14201)
);

NAND2x1p5_ASAP7_75t_L g14202 ( 
.A(n_13386),
.B(n_2046),
.Y(n_14202)
);

OAI22xp33_ASAP7_75t_L g14203 ( 
.A1(n_13755),
.A2(n_2048),
.B1(n_2046),
.B2(n_2047),
.Y(n_14203)
);

HB1xp67_ASAP7_75t_L g14204 ( 
.A(n_13560),
.Y(n_14204)
);

A2O1A1Ixp33_ASAP7_75t_L g14205 ( 
.A1(n_13534),
.A2(n_2049),
.B(n_2047),
.C(n_2048),
.Y(n_14205)
);

OAI21x1_ASAP7_75t_L g14206 ( 
.A1(n_13729),
.A2(n_2049),
.B(n_2050),
.Y(n_14206)
);

OAI21x1_ASAP7_75t_L g14207 ( 
.A1(n_13781),
.A2(n_13789),
.B(n_13780),
.Y(n_14207)
);

AND2x2_ASAP7_75t_L g14208 ( 
.A(n_13541),
.B(n_2051),
.Y(n_14208)
);

BUFx2_ASAP7_75t_L g14209 ( 
.A(n_13484),
.Y(n_14209)
);

OAI21x1_ASAP7_75t_L g14210 ( 
.A1(n_13740),
.A2(n_2051),
.B(n_2052),
.Y(n_14210)
);

HB1xp67_ASAP7_75t_L g14211 ( 
.A(n_13730),
.Y(n_14211)
);

NAND2x1p5_ASAP7_75t_L g14212 ( 
.A(n_13403),
.B(n_2052),
.Y(n_14212)
);

NAND2xp5_ASAP7_75t_L g14213 ( 
.A(n_13459),
.B(n_2053),
.Y(n_14213)
);

AND2x4_ASAP7_75t_L g14214 ( 
.A(n_13573),
.B(n_2053),
.Y(n_14214)
);

OAI22xp33_ASAP7_75t_L g14215 ( 
.A1(n_13452),
.A2(n_2056),
.B1(n_2054),
.B2(n_2055),
.Y(n_14215)
);

NAND2xp5_ASAP7_75t_SL g14216 ( 
.A(n_13622),
.B(n_13754),
.Y(n_14216)
);

OAI21x1_ASAP7_75t_L g14217 ( 
.A1(n_13812),
.A2(n_2054),
.B(n_2055),
.Y(n_14217)
);

BUFx3_ASAP7_75t_L g14218 ( 
.A(n_13469),
.Y(n_14218)
);

INVx3_ASAP7_75t_L g14219 ( 
.A(n_13648),
.Y(n_14219)
);

AND2x2_ASAP7_75t_L g14220 ( 
.A(n_13650),
.B(n_2056),
.Y(n_14220)
);

AOI221xp5_ASAP7_75t_L g14221 ( 
.A1(n_13808),
.A2(n_2059),
.B1(n_2057),
.B2(n_2058),
.C(n_2060),
.Y(n_14221)
);

OAI21x1_ASAP7_75t_L g14222 ( 
.A1(n_13746),
.A2(n_13756),
.B(n_13751),
.Y(n_14222)
);

NAND2xp5_ASAP7_75t_L g14223 ( 
.A(n_13476),
.B(n_2057),
.Y(n_14223)
);

OAI22xp5_ASAP7_75t_L g14224 ( 
.A1(n_13502),
.A2(n_2060),
.B1(n_2058),
.B2(n_2059),
.Y(n_14224)
);

BUFx2_ASAP7_75t_L g14225 ( 
.A(n_13590),
.Y(n_14225)
);

OAI21x1_ASAP7_75t_L g14226 ( 
.A1(n_13763),
.A2(n_2061),
.B(n_2062),
.Y(n_14226)
);

NOR2xp33_ASAP7_75t_L g14227 ( 
.A(n_13824),
.B(n_2061),
.Y(n_14227)
);

OAI21x1_ASAP7_75t_L g14228 ( 
.A1(n_13766),
.A2(n_2062),
.B(n_2063),
.Y(n_14228)
);

AND2x4_ASAP7_75t_L g14229 ( 
.A(n_13726),
.B(n_2063),
.Y(n_14229)
);

AOI22x1_ASAP7_75t_L g14230 ( 
.A1(n_13641),
.A2(n_2066),
.B1(n_2064),
.B2(n_2065),
.Y(n_14230)
);

OAI22xp5_ASAP7_75t_L g14231 ( 
.A1(n_13500),
.A2(n_2066),
.B1(n_2064),
.B2(n_2065),
.Y(n_14231)
);

NAND3xp33_ASAP7_75t_L g14232 ( 
.A(n_13552),
.B(n_2067),
.C(n_2068),
.Y(n_14232)
);

OAI21x1_ASAP7_75t_L g14233 ( 
.A1(n_13562),
.A2(n_2068),
.B(n_2069),
.Y(n_14233)
);

AO31x2_ASAP7_75t_L g14234 ( 
.A1(n_13606),
.A2(n_2072),
.A3(n_2070),
.B(n_2071),
.Y(n_14234)
);

OAI21x1_ASAP7_75t_L g14235 ( 
.A1(n_13479),
.A2(n_13542),
.B(n_13640),
.Y(n_14235)
);

OAI221xp5_ASAP7_75t_L g14236 ( 
.A1(n_13561),
.A2(n_2073),
.B1(n_2070),
.B2(n_2071),
.C(n_2074),
.Y(n_14236)
);

AO31x2_ASAP7_75t_L g14237 ( 
.A1(n_13596),
.A2(n_2075),
.A3(n_2073),
.B(n_2074),
.Y(n_14237)
);

A2O1A1Ixp33_ASAP7_75t_L g14238 ( 
.A1(n_13375),
.A2(n_2077),
.B(n_2075),
.C(n_2076),
.Y(n_14238)
);

BUFx4f_ASAP7_75t_SL g14239 ( 
.A(n_13813),
.Y(n_14239)
);

NAND2xp5_ASAP7_75t_L g14240 ( 
.A(n_13618),
.B(n_2077),
.Y(n_14240)
);

AOI22xp5_ASAP7_75t_L g14241 ( 
.A1(n_13465),
.A2(n_2080),
.B1(n_2078),
.B2(n_2079),
.Y(n_14241)
);

AO31x2_ASAP7_75t_L g14242 ( 
.A1(n_13669),
.A2(n_2080),
.A3(n_2078),
.B(n_2079),
.Y(n_14242)
);

INVx3_ASAP7_75t_L g14243 ( 
.A(n_13778),
.Y(n_14243)
);

INVx1_ASAP7_75t_L g14244 ( 
.A(n_13540),
.Y(n_14244)
);

INVx1_ASAP7_75t_L g14245 ( 
.A(n_13553),
.Y(n_14245)
);

INVx1_ASAP7_75t_L g14246 ( 
.A(n_13553),
.Y(n_14246)
);

OAI22xp5_ASAP7_75t_L g14247 ( 
.A1(n_13665),
.A2(n_2083),
.B1(n_2081),
.B2(n_2082),
.Y(n_14247)
);

NOR2xp33_ASAP7_75t_L g14248 ( 
.A(n_13772),
.B(n_2081),
.Y(n_14248)
);

INVx2_ASAP7_75t_L g14249 ( 
.A(n_13557),
.Y(n_14249)
);

HB1xp67_ASAP7_75t_L g14250 ( 
.A(n_13557),
.Y(n_14250)
);

INVx1_ASAP7_75t_L g14251 ( 
.A(n_13566),
.Y(n_14251)
);

AND2x4_ASAP7_75t_L g14252 ( 
.A(n_13801),
.B(n_13748),
.Y(n_14252)
);

NOR2xp33_ASAP7_75t_L g14253 ( 
.A(n_13492),
.B(n_2082),
.Y(n_14253)
);

OAI21xp5_ASAP7_75t_SL g14254 ( 
.A1(n_13424),
.A2(n_2083),
.B(n_2084),
.Y(n_14254)
);

INVx1_ASAP7_75t_L g14255 ( 
.A(n_13566),
.Y(n_14255)
);

OAI21x1_ASAP7_75t_L g14256 ( 
.A1(n_13655),
.A2(n_2084),
.B(n_2085),
.Y(n_14256)
);

OAI21x1_ASAP7_75t_L g14257 ( 
.A1(n_13634),
.A2(n_2085),
.B(n_2086),
.Y(n_14257)
);

AO31x2_ASAP7_75t_L g14258 ( 
.A1(n_13670),
.A2(n_2089),
.A3(n_2087),
.B(n_2088),
.Y(n_14258)
);

BUFx2_ASAP7_75t_L g14259 ( 
.A(n_13379),
.Y(n_14259)
);

AO21x2_ASAP7_75t_L g14260 ( 
.A1(n_13422),
.A2(n_2087),
.B(n_2088),
.Y(n_14260)
);

INVx1_ASAP7_75t_L g14261 ( 
.A(n_13392),
.Y(n_14261)
);

AO31x2_ASAP7_75t_L g14262 ( 
.A1(n_13685),
.A2(n_2091),
.A3(n_2089),
.B(n_2090),
.Y(n_14262)
);

NAND2xp5_ASAP7_75t_L g14263 ( 
.A(n_13621),
.B(n_2090),
.Y(n_14263)
);

OR2x2_ASAP7_75t_L g14264 ( 
.A(n_13790),
.B(n_2091),
.Y(n_14264)
);

NAND2xp5_ASAP7_75t_L g14265 ( 
.A(n_13621),
.B(n_2092),
.Y(n_14265)
);

OA21x2_ASAP7_75t_L g14266 ( 
.A1(n_13620),
.A2(n_2092),
.B(n_2093),
.Y(n_14266)
);

INVx2_ASAP7_75t_SL g14267 ( 
.A(n_13702),
.Y(n_14267)
);

OAI21x1_ASAP7_75t_L g14268 ( 
.A1(n_13731),
.A2(n_2093),
.B(n_2094),
.Y(n_14268)
);

INVx1_ASAP7_75t_L g14269 ( 
.A(n_13392),
.Y(n_14269)
);

NAND2xp5_ASAP7_75t_L g14270 ( 
.A(n_13305),
.B(n_2094),
.Y(n_14270)
);

AO21x2_ASAP7_75t_L g14271 ( 
.A1(n_13610),
.A2(n_13613),
.B(n_13632),
.Y(n_14271)
);

INVx3_ASAP7_75t_SL g14272 ( 
.A(n_13549),
.Y(n_14272)
);

OAI21x1_ASAP7_75t_SL g14273 ( 
.A1(n_13695),
.A2(n_2095),
.B(n_2096),
.Y(n_14273)
);

NAND2x1p5_ASAP7_75t_L g14274 ( 
.A(n_13807),
.B(n_2095),
.Y(n_14274)
);

BUFx2_ASAP7_75t_L g14275 ( 
.A(n_13379),
.Y(n_14275)
);

AND2x4_ASAP7_75t_L g14276 ( 
.A(n_13900),
.B(n_13801),
.Y(n_14276)
);

NAND2xp5_ASAP7_75t_L g14277 ( 
.A(n_13907),
.B(n_13305),
.Y(n_14277)
);

AND2x4_ASAP7_75t_L g14278 ( 
.A(n_13842),
.B(n_13748),
.Y(n_14278)
);

AOI21xp5_ASAP7_75t_L g14279 ( 
.A1(n_14005),
.A2(n_13489),
.B(n_13455),
.Y(n_14279)
);

HB1xp67_ASAP7_75t_L g14280 ( 
.A(n_13866),
.Y(n_14280)
);

INVx1_ASAP7_75t_L g14281 ( 
.A(n_13874),
.Y(n_14281)
);

O2A1O1Ixp5_ASAP7_75t_L g14282 ( 
.A1(n_14216),
.A2(n_13714),
.B(n_13830),
.C(n_13692),
.Y(n_14282)
);

AND2x2_ASAP7_75t_L g14283 ( 
.A(n_13942),
.B(n_14078),
.Y(n_14283)
);

AND2x2_ASAP7_75t_L g14284 ( 
.A(n_13928),
.B(n_13629),
.Y(n_14284)
);

OR2x2_ASAP7_75t_L g14285 ( 
.A(n_13919),
.B(n_13306),
.Y(n_14285)
);

AOI21xp5_ASAP7_75t_L g14286 ( 
.A1(n_14027),
.A2(n_13817),
.B(n_13365),
.Y(n_14286)
);

NAND2xp5_ASAP7_75t_L g14287 ( 
.A(n_14134),
.B(n_13644),
.Y(n_14287)
);

O2A1O1Ixp33_ASAP7_75t_L g14288 ( 
.A1(n_13997),
.A2(n_13515),
.B(n_13411),
.C(n_13600),
.Y(n_14288)
);

CKINVDCx12_ASAP7_75t_R g14289 ( 
.A(n_13850),
.Y(n_14289)
);

OAI21x1_ASAP7_75t_L g14290 ( 
.A1(n_13858),
.A2(n_13674),
.B(n_13821),
.Y(n_14290)
);

AND2x2_ASAP7_75t_L g14291 ( 
.A(n_13945),
.B(n_13508),
.Y(n_14291)
);

INVxp67_ASAP7_75t_L g14292 ( 
.A(n_14046),
.Y(n_14292)
);

NAND2xp5_ASAP7_75t_L g14293 ( 
.A(n_14151),
.B(n_13644),
.Y(n_14293)
);

AND2x2_ASAP7_75t_L g14294 ( 
.A(n_13981),
.B(n_13778),
.Y(n_14294)
);

AND2x2_ASAP7_75t_L g14295 ( 
.A(n_13840),
.B(n_13822),
.Y(n_14295)
);

O2A1O1Ixp33_ASAP7_75t_L g14296 ( 
.A1(n_14032),
.A2(n_13583),
.B(n_13647),
.C(n_13701),
.Y(n_14296)
);

NAND2xp5_ASAP7_75t_L g14297 ( 
.A(n_13894),
.B(n_13774),
.Y(n_14297)
);

A2O1A1Ixp33_ASAP7_75t_SL g14298 ( 
.A1(n_14097),
.A2(n_13524),
.B(n_13709),
.C(n_13803),
.Y(n_14298)
);

NAND2xp33_ASAP7_75t_SL g14299 ( 
.A(n_14259),
.B(n_13698),
.Y(n_14299)
);

INVx1_ASAP7_75t_SL g14300 ( 
.A(n_14119),
.Y(n_14300)
);

OR2x2_ASAP7_75t_L g14301 ( 
.A(n_13967),
.B(n_13306),
.Y(n_14301)
);

NAND2xp5_ASAP7_75t_L g14302 ( 
.A(n_13862),
.B(n_13774),
.Y(n_14302)
);

OAI21x1_ASAP7_75t_SL g14303 ( 
.A1(n_13839),
.A2(n_13633),
.B(n_13631),
.Y(n_14303)
);

NAND2xp5_ASAP7_75t_L g14304 ( 
.A(n_14004),
.B(n_13293),
.Y(n_14304)
);

AND2x2_ASAP7_75t_L g14305 ( 
.A(n_13850),
.B(n_13794),
.Y(n_14305)
);

NAND2x1p5_ASAP7_75t_L g14306 ( 
.A(n_13878),
.B(n_13691),
.Y(n_14306)
);

INVx1_ASAP7_75t_L g14307 ( 
.A(n_13883),
.Y(n_14307)
);

AND2x2_ASAP7_75t_L g14308 ( 
.A(n_13895),
.B(n_13794),
.Y(n_14308)
);

HB1xp67_ASAP7_75t_L g14309 ( 
.A(n_14096),
.Y(n_14309)
);

AND2x2_ASAP7_75t_L g14310 ( 
.A(n_13864),
.B(n_13311),
.Y(n_14310)
);

AND2x2_ASAP7_75t_L g14311 ( 
.A(n_13933),
.B(n_13849),
.Y(n_14311)
);

INVx1_ASAP7_75t_L g14312 ( 
.A(n_13884),
.Y(n_14312)
);

A2O1A1Ixp33_ASAP7_75t_SL g14313 ( 
.A1(n_14118),
.A2(n_13558),
.B(n_13628),
.C(n_13687),
.Y(n_14313)
);

NOR2xp33_ASAP7_75t_L g14314 ( 
.A(n_13964),
.B(n_13716),
.Y(n_14314)
);

HB1xp67_ASAP7_75t_L g14315 ( 
.A(n_14081),
.Y(n_14315)
);

O2A1O1Ixp33_ASAP7_75t_L g14316 ( 
.A1(n_14087),
.A2(n_13837),
.B(n_13739),
.C(n_13742),
.Y(n_14316)
);

NOR2xp33_ASAP7_75t_SL g14317 ( 
.A(n_13930),
.B(n_13826),
.Y(n_14317)
);

NOR2xp33_ASAP7_75t_L g14318 ( 
.A(n_13854),
.B(n_13785),
.Y(n_14318)
);

AND2x2_ASAP7_75t_L g14319 ( 
.A(n_14225),
.B(n_13311),
.Y(n_14319)
);

INVx1_ASAP7_75t_L g14320 ( 
.A(n_13893),
.Y(n_14320)
);

HB1xp67_ASAP7_75t_L g14321 ( 
.A(n_14250),
.Y(n_14321)
);

BUFx6f_ASAP7_75t_L g14322 ( 
.A(n_13988),
.Y(n_14322)
);

O2A1O1Ixp33_ASAP7_75t_L g14323 ( 
.A1(n_14185),
.A2(n_13791),
.B(n_13576),
.C(n_13595),
.Y(n_14323)
);

AND2x4_ASAP7_75t_L g14324 ( 
.A(n_13927),
.B(n_13829),
.Y(n_14324)
);

INVx2_ASAP7_75t_L g14325 ( 
.A(n_13929),
.Y(n_14325)
);

AND2x4_ASAP7_75t_L g14326 ( 
.A(n_14117),
.B(n_13829),
.Y(n_14326)
);

A2O1A1Ixp33_ASAP7_75t_L g14327 ( 
.A1(n_14033),
.A2(n_13799),
.B(n_13721),
.C(n_13719),
.Y(n_14327)
);

AOI21xp5_ASAP7_75t_L g14328 ( 
.A1(n_14137),
.A2(n_13706),
.B(n_13521),
.Y(n_14328)
);

INVx1_ASAP7_75t_L g14329 ( 
.A(n_13902),
.Y(n_14329)
);

AND2x2_ASAP7_75t_L g14330 ( 
.A(n_14102),
.B(n_13323),
.Y(n_14330)
);

AND2x4_ASAP7_75t_L g14331 ( 
.A(n_14155),
.B(n_13293),
.Y(n_14331)
);

OR2x6_ASAP7_75t_SL g14332 ( 
.A(n_14036),
.B(n_13546),
.Y(n_14332)
);

AND2x2_ASAP7_75t_L g14333 ( 
.A(n_14140),
.B(n_14145),
.Y(n_14333)
);

AOI21x1_ASAP7_75t_SL g14334 ( 
.A1(n_14270),
.A2(n_13604),
.B(n_13712),
.Y(n_14334)
);

AND2x2_ASAP7_75t_L g14335 ( 
.A(n_13962),
.B(n_13323),
.Y(n_14335)
);

AND2x2_ASAP7_75t_L g14336 ( 
.A(n_13908),
.B(n_13875),
.Y(n_14336)
);

A2O1A1Ixp33_ASAP7_75t_L g14337 ( 
.A1(n_14254),
.A2(n_14275),
.B(n_14222),
.C(n_14120),
.Y(n_14337)
);

AND2x4_ASAP7_75t_L g14338 ( 
.A(n_13876),
.B(n_13659),
.Y(n_14338)
);

INVx1_ASAP7_75t_L g14339 ( 
.A(n_13910),
.Y(n_14339)
);

OA21x2_ASAP7_75t_L g14340 ( 
.A1(n_14091),
.A2(n_13505),
.B(n_13699),
.Y(n_14340)
);

AOI21xp5_ASAP7_75t_SL g14341 ( 
.A1(n_14012),
.A2(n_13667),
.B(n_13711),
.Y(n_14341)
);

OAI22xp33_ASAP7_75t_L g14342 ( 
.A1(n_14180),
.A2(n_13973),
.B1(n_14073),
.B2(n_14204),
.Y(n_14342)
);

O2A1O1Ixp5_ASAP7_75t_L g14343 ( 
.A1(n_14135),
.A2(n_13913),
.B(n_13860),
.C(n_14057),
.Y(n_14343)
);

AND2x4_ASAP7_75t_L g14344 ( 
.A(n_13879),
.B(n_13659),
.Y(n_14344)
);

AND2x2_ASAP7_75t_L g14345 ( 
.A(n_14124),
.B(n_13710),
.Y(n_14345)
);

AND2x2_ASAP7_75t_L g14346 ( 
.A(n_14138),
.B(n_13710),
.Y(n_14346)
);

AOI21x1_ASAP7_75t_SL g14347 ( 
.A1(n_14111),
.A2(n_13604),
.B(n_13712),
.Y(n_14347)
);

INVx1_ASAP7_75t_L g14348 ( 
.A(n_13926),
.Y(n_14348)
);

INVx1_ASAP7_75t_L g14349 ( 
.A(n_13931),
.Y(n_14349)
);

NAND2xp5_ASAP7_75t_L g14350 ( 
.A(n_13855),
.B(n_13728),
.Y(n_14350)
);

AOI21xp5_ASAP7_75t_L g14351 ( 
.A1(n_14092),
.A2(n_13390),
.B(n_13384),
.Y(n_14351)
);

BUFx6f_ASAP7_75t_L g14352 ( 
.A(n_14064),
.Y(n_14352)
);

INVx1_ASAP7_75t_L g14353 ( 
.A(n_13937),
.Y(n_14353)
);

INVx1_ASAP7_75t_L g14354 ( 
.A(n_13940),
.Y(n_14354)
);

OAI22xp5_ASAP7_75t_L g14355 ( 
.A1(n_13867),
.A2(n_13703),
.B1(n_13715),
.B2(n_13708),
.Y(n_14355)
);

INVxp67_ASAP7_75t_L g14356 ( 
.A(n_14132),
.Y(n_14356)
);

AOI21xp5_ASAP7_75t_L g14357 ( 
.A1(n_13963),
.A2(n_13405),
.B(n_13391),
.Y(n_14357)
);

NAND2xp5_ASAP7_75t_L g14358 ( 
.A(n_13873),
.B(n_13906),
.Y(n_14358)
);

AOI22xp33_ASAP7_75t_L g14359 ( 
.A1(n_14271),
.A2(n_13636),
.B1(n_13686),
.B2(n_13441),
.Y(n_14359)
);

INVx1_ASAP7_75t_L g14360 ( 
.A(n_13947),
.Y(n_14360)
);

AND2x4_ASAP7_75t_L g14361 ( 
.A(n_14042),
.B(n_13728),
.Y(n_14361)
);

AOI211xp5_ASAP7_75t_L g14362 ( 
.A1(n_14215),
.A2(n_13762),
.B(n_13464),
.C(n_13527),
.Y(n_14362)
);

INVx2_ASAP7_75t_L g14363 ( 
.A(n_14024),
.Y(n_14363)
);

A2O1A1Ixp33_ASAP7_75t_L g14364 ( 
.A1(n_14133),
.A2(n_13413),
.B(n_13414),
.C(n_13733),
.Y(n_14364)
);

AOI21xp5_ASAP7_75t_L g14365 ( 
.A1(n_14062),
.A2(n_13666),
.B(n_13501),
.Y(n_14365)
);

NAND2xp5_ASAP7_75t_L g14366 ( 
.A(n_14050),
.B(n_13646),
.Y(n_14366)
);

AND2x2_ASAP7_75t_L g14367 ( 
.A(n_13887),
.B(n_14059),
.Y(n_14367)
);

INVx2_ASAP7_75t_L g14368 ( 
.A(n_13972),
.Y(n_14368)
);

OAI22xp5_ASAP7_75t_SL g14369 ( 
.A1(n_14043),
.A2(n_13421),
.B1(n_13787),
.B2(n_13589),
.Y(n_14369)
);

A2O1A1Ixp33_ASAP7_75t_L g14370 ( 
.A1(n_14066),
.A2(n_13371),
.B(n_13770),
.C(n_13646),
.Y(n_14370)
);

INVx2_ASAP7_75t_L g14371 ( 
.A(n_13983),
.Y(n_14371)
);

INVx1_ASAP7_75t_L g14372 ( 
.A(n_13949),
.Y(n_14372)
);

OR2x2_ASAP7_75t_L g14373 ( 
.A(n_13901),
.B(n_2097),
.Y(n_14373)
);

NOR2xp67_ASAP7_75t_L g14374 ( 
.A(n_13973),
.B(n_2097),
.Y(n_14374)
);

BUFx2_ASAP7_75t_L g14375 ( 
.A(n_14272),
.Y(n_14375)
);

AND2x2_ASAP7_75t_SL g14376 ( 
.A(n_13992),
.B(n_2098),
.Y(n_14376)
);

AND2x2_ASAP7_75t_L g14377 ( 
.A(n_14072),
.B(n_2098),
.Y(n_14377)
);

AOI21xp5_ASAP7_75t_L g14378 ( 
.A1(n_14175),
.A2(n_2099),
.B(n_2100),
.Y(n_14378)
);

INVx2_ASAP7_75t_L g14379 ( 
.A(n_13984),
.Y(n_14379)
);

OR2x2_ASAP7_75t_L g14380 ( 
.A(n_14082),
.B(n_2100),
.Y(n_14380)
);

AOI21xp5_ASAP7_75t_L g14381 ( 
.A1(n_14090),
.A2(n_2101),
.B(n_2103),
.Y(n_14381)
);

AND2x2_ASAP7_75t_L g14382 ( 
.A(n_13939),
.B(n_2103),
.Y(n_14382)
);

AND2x2_ASAP7_75t_L g14383 ( 
.A(n_13869),
.B(n_2104),
.Y(n_14383)
);

INVx1_ASAP7_75t_L g14384 ( 
.A(n_13960),
.Y(n_14384)
);

INVx3_ASAP7_75t_L g14385 ( 
.A(n_14115),
.Y(n_14385)
);

BUFx2_ASAP7_75t_L g14386 ( 
.A(n_13882),
.Y(n_14386)
);

INVx2_ASAP7_75t_L g14387 ( 
.A(n_13996),
.Y(n_14387)
);

BUFx3_ASAP7_75t_L g14388 ( 
.A(n_13917),
.Y(n_14388)
);

NOR2xp33_ASAP7_75t_L g14389 ( 
.A(n_13853),
.B(n_2104),
.Y(n_14389)
);

AND2x4_ASAP7_75t_L g14390 ( 
.A(n_14093),
.B(n_2105),
.Y(n_14390)
);

OR2x2_ASAP7_75t_L g14391 ( 
.A(n_13891),
.B(n_2105),
.Y(n_14391)
);

INVx1_ASAP7_75t_L g14392 ( 
.A(n_14045),
.Y(n_14392)
);

NAND2xp5_ASAP7_75t_L g14393 ( 
.A(n_14112),
.B(n_2106),
.Y(n_14393)
);

OAI22xp5_ASAP7_75t_SL g14394 ( 
.A1(n_13950),
.A2(n_2108),
.B1(n_2106),
.B2(n_2107),
.Y(n_14394)
);

AOI21xp5_ASAP7_75t_SL g14395 ( 
.A1(n_14017),
.A2(n_2107),
.B(n_2108),
.Y(n_14395)
);

AND2x2_ASAP7_75t_L g14396 ( 
.A(n_13934),
.B(n_2109),
.Y(n_14396)
);

NAND2xp5_ASAP7_75t_L g14397 ( 
.A(n_14211),
.B(n_2109),
.Y(n_14397)
);

INVx1_ASAP7_75t_L g14398 ( 
.A(n_13980),
.Y(n_14398)
);

NOR2xp67_ASAP7_75t_L g14399 ( 
.A(n_14194),
.B(n_2110),
.Y(n_14399)
);

O2A1O1Ixp5_ASAP7_75t_L g14400 ( 
.A1(n_13903),
.A2(n_2112),
.B(n_2110),
.C(n_2111),
.Y(n_14400)
);

INVx1_ASAP7_75t_L g14401 ( 
.A(n_13990),
.Y(n_14401)
);

AOI221x1_ASAP7_75t_L g14402 ( 
.A1(n_13885),
.A2(n_2113),
.B1(n_2111),
.B2(n_2112),
.C(n_2114),
.Y(n_14402)
);

OR2x2_ASAP7_75t_L g14403 ( 
.A(n_13905),
.B(n_2113),
.Y(n_14403)
);

A2O1A1Ixp33_ASAP7_75t_L g14404 ( 
.A1(n_14173),
.A2(n_2117),
.B(n_2115),
.C(n_2116),
.Y(n_14404)
);

AND2x2_ASAP7_75t_L g14405 ( 
.A(n_13852),
.B(n_2115),
.Y(n_14405)
);

A2O1A1Ixp33_ASAP7_75t_L g14406 ( 
.A1(n_14235),
.A2(n_2118),
.B(n_2116),
.C(n_2117),
.Y(n_14406)
);

INVx1_ASAP7_75t_L g14407 ( 
.A(n_13995),
.Y(n_14407)
);

AOI21xp5_ASAP7_75t_SL g14408 ( 
.A1(n_14020),
.A2(n_2118),
.B(n_2119),
.Y(n_14408)
);

INVx1_ASAP7_75t_L g14409 ( 
.A(n_13999),
.Y(n_14409)
);

INVx1_ASAP7_75t_L g14410 ( 
.A(n_14001),
.Y(n_14410)
);

INVx1_ASAP7_75t_L g14411 ( 
.A(n_14003),
.Y(n_14411)
);

BUFx6f_ASAP7_75t_L g14412 ( 
.A(n_13954),
.Y(n_14412)
);

O2A1O1Ixp33_ASAP7_75t_L g14413 ( 
.A1(n_14150),
.A2(n_2121),
.B(n_2119),
.C(n_2120),
.Y(n_14413)
);

NAND2xp5_ASAP7_75t_L g14414 ( 
.A(n_13863),
.B(n_2120),
.Y(n_14414)
);

AND2x2_ASAP7_75t_L g14415 ( 
.A(n_13909),
.B(n_2121),
.Y(n_14415)
);

INVxp67_ASAP7_75t_SL g14416 ( 
.A(n_13847),
.Y(n_14416)
);

NOR2xp33_ASAP7_75t_L g14417 ( 
.A(n_13954),
.B(n_2122),
.Y(n_14417)
);

AND2x2_ASAP7_75t_L g14418 ( 
.A(n_13978),
.B(n_2122),
.Y(n_14418)
);

INVx1_ASAP7_75t_L g14419 ( 
.A(n_14010),
.Y(n_14419)
);

AND2x2_ASAP7_75t_L g14420 ( 
.A(n_13911),
.B(n_2123),
.Y(n_14420)
);

OR2x2_ASAP7_75t_L g14421 ( 
.A(n_13890),
.B(n_2123),
.Y(n_14421)
);

AOI21xp5_ASAP7_75t_L g14422 ( 
.A1(n_14040),
.A2(n_2124),
.B(n_2125),
.Y(n_14422)
);

A2O1A1Ixp33_ASAP7_75t_SL g14423 ( 
.A1(n_14236),
.A2(n_2127),
.B(n_2125),
.C(n_2126),
.Y(n_14423)
);

NAND2xp5_ASAP7_75t_L g14424 ( 
.A(n_14196),
.B(n_2128),
.Y(n_14424)
);

O2A1O1Ixp33_ASAP7_75t_L g14425 ( 
.A1(n_14107),
.A2(n_2130),
.B(n_2128),
.C(n_2129),
.Y(n_14425)
);

NAND2xp5_ASAP7_75t_L g14426 ( 
.A(n_13904),
.B(n_13920),
.Y(n_14426)
);

OAI22xp5_ASAP7_75t_L g14427 ( 
.A1(n_14052),
.A2(n_2132),
.B1(n_2129),
.B2(n_2130),
.Y(n_14427)
);

NOR2xp67_ASAP7_75t_L g14428 ( 
.A(n_14243),
.B(n_2132),
.Y(n_14428)
);

AND2x4_ASAP7_75t_L g14429 ( 
.A(n_13989),
.B(n_2133),
.Y(n_14429)
);

INVx1_ASAP7_75t_L g14430 ( 
.A(n_14014),
.Y(n_14430)
);

INVx1_ASAP7_75t_SL g14431 ( 
.A(n_14098),
.Y(n_14431)
);

A2O1A1Ixp33_ASAP7_75t_L g14432 ( 
.A1(n_14238),
.A2(n_2135),
.B(n_2133),
.C(n_2134),
.Y(n_14432)
);

AOI21xp5_ASAP7_75t_L g14433 ( 
.A1(n_14189),
.A2(n_14199),
.B(n_14232),
.Y(n_14433)
);

O2A1O1Ixp33_ASAP7_75t_L g14434 ( 
.A1(n_14205),
.A2(n_2137),
.B(n_2134),
.C(n_2135),
.Y(n_14434)
);

AND2x4_ASAP7_75t_L g14435 ( 
.A(n_14267),
.B(n_2137),
.Y(n_14435)
);

AND2x2_ASAP7_75t_L g14436 ( 
.A(n_14103),
.B(n_2138),
.Y(n_14436)
);

INVx2_ASAP7_75t_L g14437 ( 
.A(n_14002),
.Y(n_14437)
);

AOI21xp5_ASAP7_75t_SL g14438 ( 
.A1(n_13986),
.A2(n_2138),
.B(n_2139),
.Y(n_14438)
);

AND2x2_ASAP7_75t_L g14439 ( 
.A(n_14172),
.B(n_2139),
.Y(n_14439)
);

NOR2xp67_ASAP7_75t_L g14440 ( 
.A(n_13857),
.B(n_2140),
.Y(n_14440)
);

INVx3_ASAP7_75t_L g14441 ( 
.A(n_13932),
.Y(n_14441)
);

INVx5_ASAP7_75t_L g14442 ( 
.A(n_14060),
.Y(n_14442)
);

AOI211xp5_ASAP7_75t_L g14443 ( 
.A1(n_14203),
.A2(n_2142),
.B(n_2140),
.C(n_2141),
.Y(n_14443)
);

AOI21xp5_ASAP7_75t_L g14444 ( 
.A1(n_13881),
.A2(n_2141),
.B(n_2142),
.Y(n_14444)
);

NAND2xp5_ASAP7_75t_L g14445 ( 
.A(n_13904),
.B(n_2143),
.Y(n_14445)
);

NOR2xp67_ASAP7_75t_L g14446 ( 
.A(n_13943),
.B(n_2143),
.Y(n_14446)
);

INVx2_ASAP7_75t_L g14447 ( 
.A(n_14015),
.Y(n_14447)
);

HB1xp67_ASAP7_75t_L g14448 ( 
.A(n_14252),
.Y(n_14448)
);

OA21x2_ASAP7_75t_L g14449 ( 
.A1(n_13958),
.A2(n_2144),
.B(n_2145),
.Y(n_14449)
);

A2O1A1Ixp33_ASAP7_75t_L g14450 ( 
.A1(n_14099),
.A2(n_2146),
.B(n_2144),
.C(n_2145),
.Y(n_14450)
);

INVx2_ASAP7_75t_L g14451 ( 
.A(n_14019),
.Y(n_14451)
);

AOI21xp5_ASAP7_75t_L g14452 ( 
.A1(n_14195),
.A2(n_2146),
.B(n_2147),
.Y(n_14452)
);

AND2x4_ASAP7_75t_L g14453 ( 
.A(n_14165),
.B(n_2148),
.Y(n_14453)
);

AND2x4_ASAP7_75t_L g14454 ( 
.A(n_14181),
.B(n_14201),
.Y(n_14454)
);

A2O1A1Ixp33_ASAP7_75t_SL g14455 ( 
.A1(n_14088),
.A2(n_2151),
.B(n_2149),
.C(n_2150),
.Y(n_14455)
);

INVx1_ASAP7_75t_L g14456 ( 
.A(n_14018),
.Y(n_14456)
);

HB1xp67_ASAP7_75t_L g14457 ( 
.A(n_14006),
.Y(n_14457)
);

NAND2xp5_ASAP7_75t_L g14458 ( 
.A(n_13923),
.B(n_14207),
.Y(n_14458)
);

NAND2xp5_ASAP7_75t_L g14459 ( 
.A(n_13888),
.B(n_2149),
.Y(n_14459)
);

AND2x2_ASAP7_75t_L g14460 ( 
.A(n_13914),
.B(n_2150),
.Y(n_14460)
);

NAND2xp5_ASAP7_75t_L g14461 ( 
.A(n_13851),
.B(n_13856),
.Y(n_14461)
);

INVx2_ASAP7_75t_SL g14462 ( 
.A(n_14060),
.Y(n_14462)
);

INVx2_ASAP7_75t_L g14463 ( 
.A(n_13925),
.Y(n_14463)
);

BUFx2_ASAP7_75t_L g14464 ( 
.A(n_13936),
.Y(n_14464)
);

O2A1O1Ixp5_ASAP7_75t_L g14465 ( 
.A1(n_14263),
.A2(n_2153),
.B(n_2151),
.C(n_2152),
.Y(n_14465)
);

O2A1O1Ixp5_ASAP7_75t_L g14466 ( 
.A1(n_14265),
.A2(n_2154),
.B(n_2152),
.C(n_2153),
.Y(n_14466)
);

A2O1A1Ixp33_ASAP7_75t_L g14467 ( 
.A1(n_14221),
.A2(n_2156),
.B(n_2154),
.C(n_2155),
.Y(n_14467)
);

INVx2_ASAP7_75t_L g14468 ( 
.A(n_13957),
.Y(n_14468)
);

OR2x2_ASAP7_75t_L g14469 ( 
.A(n_13915),
.B(n_2155),
.Y(n_14469)
);

INVx2_ASAP7_75t_L g14470 ( 
.A(n_13959),
.Y(n_14470)
);

INVx1_ASAP7_75t_L g14471 ( 
.A(n_14035),
.Y(n_14471)
);

AND2x2_ASAP7_75t_L g14472 ( 
.A(n_13966),
.B(n_2156),
.Y(n_14472)
);

INVx3_ASAP7_75t_L g14473 ( 
.A(n_14016),
.Y(n_14473)
);

NOR2xp33_ASAP7_75t_SL g14474 ( 
.A(n_13899),
.B(n_2157),
.Y(n_14474)
);

BUFx12f_ASAP7_75t_L g14475 ( 
.A(n_13941),
.Y(n_14475)
);

INVx1_ASAP7_75t_SL g14476 ( 
.A(n_13916),
.Y(n_14476)
);

OA21x2_ASAP7_75t_L g14477 ( 
.A1(n_13898),
.A2(n_2158),
.B(n_2159),
.Y(n_14477)
);

O2A1O1Ixp33_ASAP7_75t_L g14478 ( 
.A1(n_14071),
.A2(n_2162),
.B(n_2159),
.C(n_2161),
.Y(n_14478)
);

AND2x4_ASAP7_75t_SL g14479 ( 
.A(n_14162),
.B(n_2161),
.Y(n_14479)
);

CKINVDCx5p33_ASAP7_75t_R g14480 ( 
.A(n_13918),
.Y(n_14480)
);

AND2x2_ASAP7_75t_L g14481 ( 
.A(n_13969),
.B(n_2162),
.Y(n_14481)
);

OR2x2_ASAP7_75t_L g14482 ( 
.A(n_13971),
.B(n_2163),
.Y(n_14482)
);

AND2x2_ASAP7_75t_L g14483 ( 
.A(n_13948),
.B(n_2163),
.Y(n_14483)
);

AND2x2_ASAP7_75t_L g14484 ( 
.A(n_14030),
.B(n_2164),
.Y(n_14484)
);

A2O1A1Ixp33_ASAP7_75t_L g14485 ( 
.A1(n_13985),
.A2(n_2166),
.B(n_2164),
.C(n_2165),
.Y(n_14485)
);

AND2x4_ASAP7_75t_L g14486 ( 
.A(n_14209),
.B(n_2166),
.Y(n_14486)
);

OAI22xp5_ASAP7_75t_L g14487 ( 
.A1(n_13975),
.A2(n_2169),
.B1(n_2167),
.B2(n_2168),
.Y(n_14487)
);

A2O1A1Ixp33_ASAP7_75t_L g14488 ( 
.A1(n_14241),
.A2(n_2170),
.B(n_2167),
.C(n_2168),
.Y(n_14488)
);

AND2x2_ASAP7_75t_L g14489 ( 
.A(n_14177),
.B(n_2170),
.Y(n_14489)
);

OAI22xp5_ASAP7_75t_SL g14490 ( 
.A1(n_13924),
.A2(n_2173),
.B1(n_2171),
.B2(n_2172),
.Y(n_14490)
);

AND2x4_ASAP7_75t_L g14491 ( 
.A(n_14192),
.B(n_2171),
.Y(n_14491)
);

OR2x2_ASAP7_75t_L g14492 ( 
.A(n_13976),
.B(n_2172),
.Y(n_14492)
);

INVx1_ASAP7_75t_L g14493 ( 
.A(n_14068),
.Y(n_14493)
);

OR2x2_ASAP7_75t_L g14494 ( 
.A(n_14251),
.B(n_2174),
.Y(n_14494)
);

A2O1A1Ixp33_ASAP7_75t_L g14495 ( 
.A1(n_14217),
.A2(n_2176),
.B(n_2174),
.C(n_2175),
.Y(n_14495)
);

NAND2xp5_ASAP7_75t_L g14496 ( 
.A(n_13896),
.B(n_2176),
.Y(n_14496)
);

OA21x2_ASAP7_75t_L g14497 ( 
.A1(n_13870),
.A2(n_2177),
.B(n_2178),
.Y(n_14497)
);

OAI22xp5_ASAP7_75t_SL g14498 ( 
.A1(n_14143),
.A2(n_2179),
.B1(n_2177),
.B2(n_2178),
.Y(n_14498)
);

A2O1A1Ixp33_ASAP7_75t_SL g14499 ( 
.A1(n_14023),
.A2(n_14076),
.B(n_14123),
.C(n_14153),
.Y(n_14499)
);

A2O1A1Ixp33_ASAP7_75t_L g14500 ( 
.A1(n_14226),
.A2(n_2182),
.B(n_2179),
.C(n_2181),
.Y(n_14500)
);

INVx1_ASAP7_75t_L g14501 ( 
.A(n_14070),
.Y(n_14501)
);

AND2x2_ASAP7_75t_L g14502 ( 
.A(n_14219),
.B(n_2181),
.Y(n_14502)
);

NAND2xp5_ASAP7_75t_L g14503 ( 
.A(n_13848),
.B(n_13844),
.Y(n_14503)
);

A2O1A1Ixp33_ASAP7_75t_L g14504 ( 
.A1(n_14228),
.A2(n_2184),
.B(n_2182),
.C(n_2183),
.Y(n_14504)
);

AND2x2_ASAP7_75t_L g14505 ( 
.A(n_13841),
.B(n_13955),
.Y(n_14505)
);

OR2x2_ASAP7_75t_L g14506 ( 
.A(n_14255),
.B(n_2183),
.Y(n_14506)
);

OR2x2_ASAP7_75t_L g14507 ( 
.A(n_14261),
.B(n_2184),
.Y(n_14507)
);

HB1xp67_ASAP7_75t_L g14508 ( 
.A(n_14170),
.Y(n_14508)
);

AND2x2_ASAP7_75t_L g14509 ( 
.A(n_13961),
.B(n_2185),
.Y(n_14509)
);

INVx1_ASAP7_75t_L g14510 ( 
.A(n_14085),
.Y(n_14510)
);

NOR2xp33_ASAP7_75t_SL g14511 ( 
.A(n_13938),
.B(n_2186),
.Y(n_14511)
);

NOR2xp67_ASAP7_75t_L g14512 ( 
.A(n_14269),
.B(n_2186),
.Y(n_14512)
);

AND2x4_ASAP7_75t_L g14513 ( 
.A(n_14218),
.B(n_2187),
.Y(n_14513)
);

A2O1A1Ixp33_ASAP7_75t_L g14514 ( 
.A1(n_14256),
.A2(n_2189),
.B(n_2187),
.C(n_2188),
.Y(n_14514)
);

INVx1_ASAP7_75t_SL g14515 ( 
.A(n_13974),
.Y(n_14515)
);

OA21x2_ASAP7_75t_L g14516 ( 
.A1(n_13872),
.A2(n_13886),
.B(n_13877),
.Y(n_14516)
);

NAND2xp5_ASAP7_75t_L g14517 ( 
.A(n_14000),
.B(n_2188),
.Y(n_14517)
);

OA21x2_ASAP7_75t_L g14518 ( 
.A1(n_13897),
.A2(n_2190),
.B(n_2192),
.Y(n_14518)
);

OR2x2_ASAP7_75t_L g14519 ( 
.A(n_14169),
.B(n_2192),
.Y(n_14519)
);

BUFx2_ASAP7_75t_L g14520 ( 
.A(n_13951),
.Y(n_14520)
);

OA21x2_ASAP7_75t_L g14521 ( 
.A1(n_14142),
.A2(n_2193),
.B(n_2194),
.Y(n_14521)
);

A2O1A1Ixp33_ASAP7_75t_L g14522 ( 
.A1(n_14253),
.A2(n_2196),
.B(n_2194),
.C(n_2195),
.Y(n_14522)
);

INVx5_ASAP7_75t_L g14523 ( 
.A(n_14161),
.Y(n_14523)
);

AOI221xp5_ASAP7_75t_L g14524 ( 
.A1(n_13843),
.A2(n_2197),
.B1(n_2195),
.B2(n_2196),
.C(n_2198),
.Y(n_14524)
);

INVx2_ASAP7_75t_L g14525 ( 
.A(n_14029),
.Y(n_14525)
);

AND2x2_ASAP7_75t_L g14526 ( 
.A(n_13865),
.B(n_2197),
.Y(n_14526)
);

NAND2xp5_ASAP7_75t_L g14527 ( 
.A(n_14011),
.B(n_2198),
.Y(n_14527)
);

NOR2xp33_ASAP7_75t_L g14528 ( 
.A(n_13977),
.B(n_2199),
.Y(n_14528)
);

A2O1A1Ixp33_ASAP7_75t_L g14529 ( 
.A1(n_13944),
.A2(n_2201),
.B(n_2199),
.C(n_2200),
.Y(n_14529)
);

O2A1O1Ixp33_ASAP7_75t_L g14530 ( 
.A1(n_14193),
.A2(n_2202),
.B(n_2200),
.C(n_2201),
.Y(n_14530)
);

NAND2xp5_ASAP7_75t_L g14531 ( 
.A(n_14065),
.B(n_2202),
.Y(n_14531)
);

AND2x2_ASAP7_75t_L g14532 ( 
.A(n_13865),
.B(n_2203),
.Y(n_14532)
);

NOR2xp33_ASAP7_75t_L g14533 ( 
.A(n_13987),
.B(n_2203),
.Y(n_14533)
);

O2A1O1Ixp5_ASAP7_75t_L g14534 ( 
.A1(n_14026),
.A2(n_2206),
.B(n_2204),
.C(n_2205),
.Y(n_14534)
);

AND2x2_ASAP7_75t_L g14535 ( 
.A(n_13953),
.B(n_2204),
.Y(n_14535)
);

NOR2xp33_ASAP7_75t_L g14536 ( 
.A(n_13922),
.B(n_2205),
.Y(n_14536)
);

AND2x2_ASAP7_75t_L g14537 ( 
.A(n_13979),
.B(n_13968),
.Y(n_14537)
);

AOI21xp5_ASAP7_75t_L g14538 ( 
.A1(n_13859),
.A2(n_2207),
.B(n_2208),
.Y(n_14538)
);

AOI21xp5_ASAP7_75t_L g14539 ( 
.A1(n_13846),
.A2(n_2207),
.B(n_2209),
.Y(n_14539)
);

INVx1_ASAP7_75t_L g14540 ( 
.A(n_14163),
.Y(n_14540)
);

NAND2xp5_ASAP7_75t_L g14541 ( 
.A(n_14106),
.B(n_2209),
.Y(n_14541)
);

NAND2xp5_ASAP7_75t_L g14542 ( 
.A(n_14167),
.B(n_2210),
.Y(n_14542)
);

CKINVDCx11_ASAP7_75t_R g14543 ( 
.A(n_14013),
.Y(n_14543)
);

INVx2_ASAP7_75t_SL g14544 ( 
.A(n_13993),
.Y(n_14544)
);

OR2x2_ASAP7_75t_L g14545 ( 
.A(n_14171),
.B(n_2210),
.Y(n_14545)
);

A2O1A1Ixp33_ASAP7_75t_L g14546 ( 
.A1(n_14039),
.A2(n_2213),
.B(n_2211),
.C(n_2212),
.Y(n_14546)
);

OR2x2_ASAP7_75t_L g14547 ( 
.A(n_14184),
.B(n_2212),
.Y(n_14547)
);

AND2x2_ASAP7_75t_L g14548 ( 
.A(n_13993),
.B(n_2213),
.Y(n_14548)
);

INVx2_ASAP7_75t_L g14549 ( 
.A(n_14025),
.Y(n_14549)
);

AOI21xp5_ASAP7_75t_SL g14550 ( 
.A1(n_14031),
.A2(n_2214),
.B(n_2215),
.Y(n_14550)
);

INVx2_ASAP7_75t_L g14551 ( 
.A(n_13952),
.Y(n_14551)
);

INVx3_ASAP7_75t_L g14552 ( 
.A(n_14114),
.Y(n_14552)
);

OAI21x1_ASAP7_75t_SL g14553 ( 
.A1(n_13912),
.A2(n_2215),
.B(n_2216),
.Y(n_14553)
);

AND2x2_ASAP7_75t_L g14554 ( 
.A(n_14114),
.B(n_2216),
.Y(n_14554)
);

AND2x2_ASAP7_75t_L g14555 ( 
.A(n_14121),
.B(n_2217),
.Y(n_14555)
);

AND2x2_ASAP7_75t_L g14556 ( 
.A(n_14121),
.B(n_2217),
.Y(n_14556)
);

INVx2_ASAP7_75t_L g14557 ( 
.A(n_13991),
.Y(n_14557)
);

INVx1_ASAP7_75t_L g14558 ( 
.A(n_14244),
.Y(n_14558)
);

AND2x2_ASAP7_75t_L g14559 ( 
.A(n_14058),
.B(n_2218),
.Y(n_14559)
);

HB1xp67_ASAP7_75t_L g14560 ( 
.A(n_14249),
.Y(n_14560)
);

INVx1_ASAP7_75t_L g14561 ( 
.A(n_14245),
.Y(n_14561)
);

AND2x2_ASAP7_75t_L g14562 ( 
.A(n_13982),
.B(n_2218),
.Y(n_14562)
);

NOR2x2_ASAP7_75t_L g14563 ( 
.A(n_14160),
.B(n_2219),
.Y(n_14563)
);

OR2x2_ASAP7_75t_L g14564 ( 
.A(n_14246),
.B(n_2220),
.Y(n_14564)
);

AND2x2_ASAP7_75t_L g14565 ( 
.A(n_14067),
.B(n_2220),
.Y(n_14565)
);

AND2x2_ASAP7_75t_L g14566 ( 
.A(n_13935),
.B(n_2221),
.Y(n_14566)
);

AND2x4_ASAP7_75t_L g14567 ( 
.A(n_13956),
.B(n_14104),
.Y(n_14567)
);

NAND2xp5_ASAP7_75t_L g14568 ( 
.A(n_14168),
.B(n_2221),
.Y(n_14568)
);

AND2x2_ASAP7_75t_L g14569 ( 
.A(n_14041),
.B(n_2222),
.Y(n_14569)
);

OAI22xp5_ASAP7_75t_L g14570 ( 
.A1(n_13970),
.A2(n_14230),
.B1(n_13998),
.B2(n_14224),
.Y(n_14570)
);

AOI21xp5_ASAP7_75t_L g14571 ( 
.A1(n_13868),
.A2(n_2222),
.B(n_2223),
.Y(n_14571)
);

NAND2xp5_ASAP7_75t_L g14572 ( 
.A(n_14009),
.B(n_2223),
.Y(n_14572)
);

INVx2_ASAP7_75t_L g14573 ( 
.A(n_14089),
.Y(n_14573)
);

OAI22xp5_ASAP7_75t_L g14574 ( 
.A1(n_14190),
.A2(n_2226),
.B1(n_2224),
.B2(n_2225),
.Y(n_14574)
);

A2O1A1Ixp33_ASAP7_75t_SL g14575 ( 
.A1(n_14110),
.A2(n_2226),
.B(n_2224),
.C(n_2225),
.Y(n_14575)
);

AND2x2_ASAP7_75t_L g14576 ( 
.A(n_13889),
.B(n_2227),
.Y(n_14576)
);

INVx1_ASAP7_75t_L g14577 ( 
.A(n_14008),
.Y(n_14577)
);

AND2x2_ASAP7_75t_L g14578 ( 
.A(n_13892),
.B(n_2227),
.Y(n_14578)
);

INVx2_ASAP7_75t_L g14579 ( 
.A(n_14049),
.Y(n_14579)
);

AND2x2_ASAP7_75t_L g14580 ( 
.A(n_14044),
.B(n_2228),
.Y(n_14580)
);

AND2x2_ASAP7_75t_L g14581 ( 
.A(n_14051),
.B(n_2228),
.Y(n_14581)
);

AND2x2_ASAP7_75t_L g14582 ( 
.A(n_13871),
.B(n_14126),
.Y(n_14582)
);

AND2x4_ASAP7_75t_L g14583 ( 
.A(n_14022),
.B(n_14108),
.Y(n_14583)
);

AND2x2_ASAP7_75t_L g14584 ( 
.A(n_14136),
.B(n_14188),
.Y(n_14584)
);

BUFx6f_ASAP7_75t_L g14585 ( 
.A(n_14075),
.Y(n_14585)
);

INVx2_ASAP7_75t_L g14586 ( 
.A(n_14053),
.Y(n_14586)
);

BUFx8_ASAP7_75t_SL g14587 ( 
.A(n_14054),
.Y(n_14587)
);

A2O1A1Ixp33_ASAP7_75t_L g14588 ( 
.A1(n_14100),
.A2(n_2231),
.B(n_2229),
.C(n_2230),
.Y(n_14588)
);

AND2x2_ASAP7_75t_L g14589 ( 
.A(n_13965),
.B(n_2229),
.Y(n_14589)
);

O2A1O1Ixp33_ASAP7_75t_L g14590 ( 
.A1(n_14080),
.A2(n_2232),
.B(n_2230),
.C(n_2231),
.Y(n_14590)
);

AND2x2_ASAP7_75t_L g14591 ( 
.A(n_14220),
.B(n_2232),
.Y(n_14591)
);

BUFx3_ASAP7_75t_L g14592 ( 
.A(n_14239),
.Y(n_14592)
);

INVxp67_ASAP7_75t_L g14593 ( 
.A(n_14061),
.Y(n_14593)
);

OR2x6_ASAP7_75t_L g14594 ( 
.A(n_14007),
.B(n_2233),
.Y(n_14594)
);

OAI22xp5_ASAP7_75t_L g14595 ( 
.A1(n_14113),
.A2(n_2235),
.B1(n_2233),
.B2(n_2234),
.Y(n_14595)
);

INVx2_ASAP7_75t_L g14596 ( 
.A(n_14122),
.Y(n_14596)
);

OAI22xp5_ASAP7_75t_SL g14597 ( 
.A1(n_13845),
.A2(n_2236),
.B1(n_2234),
.B2(n_2235),
.Y(n_14597)
);

CKINVDCx20_ASAP7_75t_R g14598 ( 
.A(n_13861),
.Y(n_14598)
);

A2O1A1Ixp33_ASAP7_75t_L g14599 ( 
.A1(n_14248),
.A2(n_2238),
.B(n_2236),
.C(n_2237),
.Y(n_14599)
);

O2A1O1Ixp33_ASAP7_75t_L g14600 ( 
.A1(n_14094),
.A2(n_2239),
.B(n_2237),
.C(n_2238),
.Y(n_14600)
);

BUFx3_ASAP7_75t_L g14601 ( 
.A(n_14214),
.Y(n_14601)
);

AOI211xp5_ASAP7_75t_L g14602 ( 
.A1(n_14247),
.A2(n_2241),
.B(n_2239),
.C(n_2240),
.Y(n_14602)
);

AND2x2_ASAP7_75t_L g14603 ( 
.A(n_13921),
.B(n_2240),
.Y(n_14603)
);

INVx1_ASAP7_75t_L g14604 ( 
.A(n_14074),
.Y(n_14604)
);

NAND2xp5_ASAP7_75t_L g14605 ( 
.A(n_14125),
.B(n_2241),
.Y(n_14605)
);

NAND2xp5_ASAP7_75t_L g14606 ( 
.A(n_14131),
.B(n_2242),
.Y(n_14606)
);

AND2x2_ASAP7_75t_L g14607 ( 
.A(n_14208),
.B(n_2242),
.Y(n_14607)
);

INVx5_ASAP7_75t_L g14608 ( 
.A(n_14191),
.Y(n_14608)
);

OR2x2_ASAP7_75t_L g14609 ( 
.A(n_14047),
.B(n_2243),
.Y(n_14609)
);

AND2x2_ASAP7_75t_L g14610 ( 
.A(n_14229),
.B(n_2243),
.Y(n_14610)
);

INVx2_ASAP7_75t_L g14611 ( 
.A(n_14084),
.Y(n_14611)
);

AOI21xp5_ASAP7_75t_SL g14612 ( 
.A1(n_14266),
.A2(n_2244),
.B(n_2245),
.Y(n_14612)
);

BUFx12f_ASAP7_75t_L g14613 ( 
.A(n_14264),
.Y(n_14613)
);

O2A1O1Ixp5_ASAP7_75t_L g14614 ( 
.A1(n_13994),
.A2(n_2247),
.B(n_2245),
.C(n_2246),
.Y(n_14614)
);

AND2x2_ASAP7_75t_L g14615 ( 
.A(n_14157),
.B(n_14164),
.Y(n_14615)
);

OAI22xp5_ASAP7_75t_L g14616 ( 
.A1(n_14198),
.A2(n_14202),
.B1(n_14212),
.B2(n_14182),
.Y(n_14616)
);

BUFx12f_ASAP7_75t_L g14617 ( 
.A(n_14048),
.Y(n_14617)
);

AND2x2_ASAP7_75t_L g14618 ( 
.A(n_14166),
.B(n_2246),
.Y(n_14618)
);

A2O1A1Ixp33_ASAP7_75t_SL g14619 ( 
.A1(n_14197),
.A2(n_2249),
.B(n_2247),
.C(n_2248),
.Y(n_14619)
);

NOR2xp33_ASAP7_75t_SL g14620 ( 
.A(n_14147),
.B(n_2249),
.Y(n_14620)
);

NAND2xp5_ASAP7_75t_L g14621 ( 
.A(n_13880),
.B(n_2250),
.Y(n_14621)
);

BUFx2_ASAP7_75t_L g14622 ( 
.A(n_14237),
.Y(n_14622)
);

BUFx6f_ASAP7_75t_L g14623 ( 
.A(n_14139),
.Y(n_14623)
);

INVx3_ASAP7_75t_L g14624 ( 
.A(n_14210),
.Y(n_14624)
);

AND2x2_ASAP7_75t_L g14625 ( 
.A(n_14158),
.B(n_2250),
.Y(n_14625)
);

CKINVDCx5p33_ASAP7_75t_R g14626 ( 
.A(n_14028),
.Y(n_14626)
);

OA21x2_ASAP7_75t_L g14627 ( 
.A1(n_14240),
.A2(n_2251),
.B(n_2252),
.Y(n_14627)
);

O2A1O1Ixp33_ASAP7_75t_L g14628 ( 
.A1(n_14159),
.A2(n_2255),
.B(n_2251),
.C(n_2254),
.Y(n_14628)
);

OR2x2_ASAP7_75t_L g14629 ( 
.A(n_14128),
.B(n_2254),
.Y(n_14629)
);

AOI21xp5_ASAP7_75t_L g14630 ( 
.A1(n_14260),
.A2(n_2255),
.B(n_2256),
.Y(n_14630)
);

AND2x2_ASAP7_75t_L g14631 ( 
.A(n_14174),
.B(n_2256),
.Y(n_14631)
);

AND2x2_ASAP7_75t_L g14632 ( 
.A(n_14178),
.B(n_2258),
.Y(n_14632)
);

BUFx6f_ASAP7_75t_L g14633 ( 
.A(n_14179),
.Y(n_14633)
);

OAI22xp5_ASAP7_75t_L g14634 ( 
.A1(n_14274),
.A2(n_2260),
.B1(n_2258),
.B2(n_2259),
.Y(n_14634)
);

BUFx8_ASAP7_75t_L g14635 ( 
.A(n_14063),
.Y(n_14635)
);

CKINVDCx5p33_ASAP7_75t_R g14636 ( 
.A(n_14227),
.Y(n_14636)
);

HB1xp67_ASAP7_75t_L g14637 ( 
.A(n_14129),
.Y(n_14637)
);

INVx3_ASAP7_75t_L g14638 ( 
.A(n_14186),
.Y(n_14638)
);

NOR2xp33_ASAP7_75t_L g14639 ( 
.A(n_14079),
.B(n_2260),
.Y(n_14639)
);

NOR2xp33_ASAP7_75t_SL g14640 ( 
.A(n_14105),
.B(n_2261),
.Y(n_14640)
);

INVx2_ASAP7_75t_L g14641 ( 
.A(n_14187),
.Y(n_14641)
);

O2A1O1Ixp5_ASAP7_75t_L g14642 ( 
.A1(n_14101),
.A2(n_2263),
.B(n_2261),
.C(n_2262),
.Y(n_14642)
);

AOI21xp5_ASAP7_75t_L g14643 ( 
.A1(n_14056),
.A2(n_2263),
.B(n_2264),
.Y(n_14643)
);

OAI22xp5_ASAP7_75t_L g14644 ( 
.A1(n_14231),
.A2(n_2266),
.B1(n_2264),
.B2(n_2265),
.Y(n_14644)
);

AND2x2_ASAP7_75t_L g14645 ( 
.A(n_14206),
.B(n_2266),
.Y(n_14645)
);

AND2x2_ASAP7_75t_SL g14646 ( 
.A(n_14116),
.B(n_2267),
.Y(n_14646)
);

INVx2_ASAP7_75t_SL g14647 ( 
.A(n_14146),
.Y(n_14647)
);

INVx1_ASAP7_75t_L g14648 ( 
.A(n_14141),
.Y(n_14648)
);

AND2x4_ASAP7_75t_L g14649 ( 
.A(n_14055),
.B(n_2267),
.Y(n_14649)
);

INVx1_ASAP7_75t_L g14650 ( 
.A(n_14144),
.Y(n_14650)
);

INVx2_ASAP7_75t_L g14651 ( 
.A(n_14021),
.Y(n_14651)
);

OAI21xp5_ASAP7_75t_L g14652 ( 
.A1(n_14268),
.A2(n_2268),
.B(n_2270),
.Y(n_14652)
);

O2A1O1Ixp33_ASAP7_75t_L g14653 ( 
.A1(n_14176),
.A2(n_2271),
.B(n_2268),
.C(n_2270),
.Y(n_14653)
);

AND2x4_ASAP7_75t_L g14654 ( 
.A(n_14109),
.B(n_2271),
.Y(n_14654)
);

A2O1A1Ixp33_ASAP7_75t_L g14655 ( 
.A1(n_14257),
.A2(n_2275),
.B(n_2272),
.C(n_2274),
.Y(n_14655)
);

INVx1_ASAP7_75t_L g14656 ( 
.A(n_14148),
.Y(n_14656)
);

AOI21xp5_ASAP7_75t_L g14657 ( 
.A1(n_14038),
.A2(n_2272),
.B(n_2274),
.Y(n_14657)
);

INVx4_ASAP7_75t_L g14658 ( 
.A(n_14273),
.Y(n_14658)
);

AOI21xp5_ASAP7_75t_SL g14659 ( 
.A1(n_14156),
.A2(n_2275),
.B(n_2276),
.Y(n_14659)
);

A2O1A1Ixp33_ASAP7_75t_L g14660 ( 
.A1(n_14149),
.A2(n_2279),
.B(n_2277),
.C(n_2278),
.Y(n_14660)
);

AOI21xp5_ASAP7_75t_L g14661 ( 
.A1(n_14183),
.A2(n_2277),
.B(n_2278),
.Y(n_14661)
);

OA21x2_ASAP7_75t_L g14662 ( 
.A1(n_14233),
.A2(n_2280),
.B(n_2281),
.Y(n_14662)
);

AOI221x1_ASAP7_75t_L g14663 ( 
.A1(n_14200),
.A2(n_2283),
.B1(n_2280),
.B2(n_2282),
.C(n_2284),
.Y(n_14663)
);

INVx1_ASAP7_75t_L g14664 ( 
.A(n_14493),
.Y(n_14664)
);

INVx2_ASAP7_75t_L g14665 ( 
.A(n_14375),
.Y(n_14665)
);

INVx1_ASAP7_75t_L g14666 ( 
.A(n_14501),
.Y(n_14666)
);

AND2x2_ASAP7_75t_L g14667 ( 
.A(n_14431),
.B(n_14237),
.Y(n_14667)
);

AND2x2_ASAP7_75t_L g14668 ( 
.A(n_14283),
.B(n_14154),
.Y(n_14668)
);

OR2x2_ASAP7_75t_L g14669 ( 
.A(n_14280),
.B(n_14557),
.Y(n_14669)
);

INVx1_ASAP7_75t_L g14670 ( 
.A(n_14510),
.Y(n_14670)
);

AND2x2_ASAP7_75t_L g14671 ( 
.A(n_14333),
.B(n_14130),
.Y(n_14671)
);

HB1xp67_ASAP7_75t_L g14672 ( 
.A(n_14309),
.Y(n_14672)
);

INVx1_ASAP7_75t_L g14673 ( 
.A(n_14540),
.Y(n_14673)
);

INVx2_ASAP7_75t_L g14674 ( 
.A(n_14442),
.Y(n_14674)
);

NAND2xp5_ASAP7_75t_L g14675 ( 
.A(n_14535),
.B(n_14213),
.Y(n_14675)
);

OAI21x1_ASAP7_75t_L g14676 ( 
.A1(n_14363),
.A2(n_14037),
.B(n_14034),
.Y(n_14676)
);

INVx2_ASAP7_75t_L g14677 ( 
.A(n_14442),
.Y(n_14677)
);

INVx1_ASAP7_75t_L g14678 ( 
.A(n_14558),
.Y(n_14678)
);

INVx3_ASAP7_75t_L g14679 ( 
.A(n_14322),
.Y(n_14679)
);

INVx3_ASAP7_75t_L g14680 ( 
.A(n_14322),
.Y(n_14680)
);

INVx1_ASAP7_75t_L g14681 ( 
.A(n_14561),
.Y(n_14681)
);

NAND2xp5_ASAP7_75t_L g14682 ( 
.A(n_14286),
.B(n_14223),
.Y(n_14682)
);

INVx2_ASAP7_75t_L g14683 ( 
.A(n_14462),
.Y(n_14683)
);

HB1xp67_ASAP7_75t_L g14684 ( 
.A(n_14315),
.Y(n_14684)
);

INVx1_ASAP7_75t_L g14685 ( 
.A(n_14281),
.Y(n_14685)
);

OR2x6_ASAP7_75t_L g14686 ( 
.A(n_14438),
.B(n_14077),
.Y(n_14686)
);

OAI22xp5_ASAP7_75t_L g14687 ( 
.A1(n_14337),
.A2(n_14152),
.B1(n_13946),
.B2(n_14242),
.Y(n_14687)
);

INVx2_ASAP7_75t_SL g14688 ( 
.A(n_14352),
.Y(n_14688)
);

INVx2_ASAP7_75t_L g14689 ( 
.A(n_14520),
.Y(n_14689)
);

INVxp67_ASAP7_75t_L g14690 ( 
.A(n_14511),
.Y(n_14690)
);

INVx3_ASAP7_75t_L g14691 ( 
.A(n_14352),
.Y(n_14691)
);

INVx3_ASAP7_75t_L g14692 ( 
.A(n_14592),
.Y(n_14692)
);

NOR2xp33_ASAP7_75t_L g14693 ( 
.A(n_14386),
.B(n_14083),
.Y(n_14693)
);

INVx3_ASAP7_75t_L g14694 ( 
.A(n_14412),
.Y(n_14694)
);

INVx2_ASAP7_75t_L g14695 ( 
.A(n_14385),
.Y(n_14695)
);

INVx2_ASAP7_75t_L g14696 ( 
.A(n_14311),
.Y(n_14696)
);

CKINVDCx5p33_ASAP7_75t_R g14697 ( 
.A(n_14543),
.Y(n_14697)
);

OA21x2_ASAP7_75t_L g14698 ( 
.A1(n_14343),
.A2(n_14095),
.B(n_14086),
.Y(n_14698)
);

BUFx6f_ASAP7_75t_L g14699 ( 
.A(n_14412),
.Y(n_14699)
);

INVx1_ASAP7_75t_L g14700 ( 
.A(n_14307),
.Y(n_14700)
);

INVx2_ASAP7_75t_L g14701 ( 
.A(n_14441),
.Y(n_14701)
);

INVx2_ASAP7_75t_L g14702 ( 
.A(n_14454),
.Y(n_14702)
);

INVx1_ASAP7_75t_L g14703 ( 
.A(n_14312),
.Y(n_14703)
);

HB1xp67_ASAP7_75t_L g14704 ( 
.A(n_14321),
.Y(n_14704)
);

INVx1_ASAP7_75t_L g14705 ( 
.A(n_14320),
.Y(n_14705)
);

INVxp67_ASAP7_75t_SL g14706 ( 
.A(n_14399),
.Y(n_14706)
);

INVx2_ASAP7_75t_L g14707 ( 
.A(n_14552),
.Y(n_14707)
);

INVx3_ASAP7_75t_L g14708 ( 
.A(n_14388),
.Y(n_14708)
);

AO31x2_ASAP7_75t_L g14709 ( 
.A1(n_14622),
.A2(n_14152),
.A3(n_14234),
.B(n_14242),
.Y(n_14709)
);

OAI21x1_ASAP7_75t_L g14710 ( 
.A1(n_14306),
.A2(n_14069),
.B(n_14127),
.Y(n_14710)
);

INVx1_ASAP7_75t_L g14711 ( 
.A(n_14329),
.Y(n_14711)
);

INVx2_ASAP7_75t_L g14712 ( 
.A(n_14367),
.Y(n_14712)
);

INVx1_ASAP7_75t_L g14713 ( 
.A(n_14339),
.Y(n_14713)
);

INVx2_ASAP7_75t_L g14714 ( 
.A(n_14567),
.Y(n_14714)
);

INVx1_ASAP7_75t_L g14715 ( 
.A(n_14348),
.Y(n_14715)
);

INVx2_ASAP7_75t_L g14716 ( 
.A(n_14523),
.Y(n_14716)
);

BUFx2_ASAP7_75t_L g14717 ( 
.A(n_14587),
.Y(n_14717)
);

INVx1_ASAP7_75t_L g14718 ( 
.A(n_14349),
.Y(n_14718)
);

INVx4_ASAP7_75t_SL g14719 ( 
.A(n_14464),
.Y(n_14719)
);

INVx1_ASAP7_75t_L g14720 ( 
.A(n_14353),
.Y(n_14720)
);

NAND2x1p5_ASAP7_75t_L g14721 ( 
.A(n_14294),
.B(n_13946),
.Y(n_14721)
);

OR2x2_ASAP7_75t_L g14722 ( 
.A(n_14549),
.B(n_14258),
.Y(n_14722)
);

INVx1_ASAP7_75t_L g14723 ( 
.A(n_14354),
.Y(n_14723)
);

INVx1_ASAP7_75t_L g14724 ( 
.A(n_14360),
.Y(n_14724)
);

OA21x2_ASAP7_75t_L g14725 ( 
.A1(n_14356),
.A2(n_14234),
.B(n_14258),
.Y(n_14725)
);

OAI21xp5_ASAP7_75t_L g14726 ( 
.A1(n_14376),
.A2(n_14282),
.B(n_14279),
.Y(n_14726)
);

INVx1_ASAP7_75t_L g14727 ( 
.A(n_14372),
.Y(n_14727)
);

NAND4xp25_ASAP7_75t_L g14728 ( 
.A(n_14323),
.B(n_14262),
.C(n_2284),
.D(n_2282),
.Y(n_14728)
);

BUFx3_ASAP7_75t_L g14729 ( 
.A(n_14475),
.Y(n_14729)
);

INVx2_ASAP7_75t_L g14730 ( 
.A(n_14523),
.Y(n_14730)
);

INVx1_ASAP7_75t_L g14731 ( 
.A(n_14384),
.Y(n_14731)
);

INVx1_ASAP7_75t_L g14732 ( 
.A(n_14401),
.Y(n_14732)
);

INVx2_ASAP7_75t_L g14733 ( 
.A(n_14608),
.Y(n_14733)
);

BUFx2_ASAP7_75t_SL g14734 ( 
.A(n_14374),
.Y(n_14734)
);

OAI21xp33_ASAP7_75t_SL g14735 ( 
.A1(n_14426),
.A2(n_14262),
.B(n_2283),
.Y(n_14735)
);

AOI22xp33_ASAP7_75t_SL g14736 ( 
.A1(n_14490),
.A2(n_2287),
.B1(n_2285),
.B2(n_2286),
.Y(n_14736)
);

AOI22xp33_ASAP7_75t_SL g14737 ( 
.A1(n_14284),
.A2(n_2289),
.B1(n_2287),
.B2(n_2288),
.Y(n_14737)
);

BUFx3_ASAP7_75t_L g14738 ( 
.A(n_14584),
.Y(n_14738)
);

INVx1_ASAP7_75t_L g14739 ( 
.A(n_14407),
.Y(n_14739)
);

INVx2_ASAP7_75t_L g14740 ( 
.A(n_14608),
.Y(n_14740)
);

OAI21x1_ASAP7_75t_L g14741 ( 
.A1(n_14551),
.A2(n_2288),
.B(n_2289),
.Y(n_14741)
);

INVx1_ASAP7_75t_L g14742 ( 
.A(n_14409),
.Y(n_14742)
);

INVx1_ASAP7_75t_L g14743 ( 
.A(n_14410),
.Y(n_14743)
);

OR2x6_ASAP7_75t_L g14744 ( 
.A(n_14341),
.B(n_2290),
.Y(n_14744)
);

INVx1_ASAP7_75t_L g14745 ( 
.A(n_14411),
.Y(n_14745)
);

CKINVDCx11_ASAP7_75t_R g14746 ( 
.A(n_14300),
.Y(n_14746)
);

AOI22xp33_ASAP7_75t_L g14747 ( 
.A1(n_14299),
.A2(n_2292),
.B1(n_2290),
.B2(n_2291),
.Y(n_14747)
);

AO21x2_ASAP7_75t_L g14748 ( 
.A1(n_14572),
.A2(n_2291),
.B(n_2293),
.Y(n_14748)
);

HB1xp67_ASAP7_75t_L g14749 ( 
.A(n_14457),
.Y(n_14749)
);

INVx1_ASAP7_75t_L g14750 ( 
.A(n_14419),
.Y(n_14750)
);

HB1xp67_ASAP7_75t_L g14751 ( 
.A(n_14440),
.Y(n_14751)
);

INVxp67_ASAP7_75t_L g14752 ( 
.A(n_14291),
.Y(n_14752)
);

AND2x2_ASAP7_75t_L g14753 ( 
.A(n_14336),
.B(n_2293),
.Y(n_14753)
);

AND2x6_ASAP7_75t_L g14754 ( 
.A(n_14515),
.B(n_2294),
.Y(n_14754)
);

NOR2x1_ASAP7_75t_SL g14755 ( 
.A(n_14617),
.B(n_2294),
.Y(n_14755)
);

AND2x2_ASAP7_75t_L g14756 ( 
.A(n_14537),
.B(n_2295),
.Y(n_14756)
);

OAI21xp5_ASAP7_75t_L g14757 ( 
.A1(n_14327),
.A2(n_2295),
.B(n_2296),
.Y(n_14757)
);

BUFx2_ASAP7_75t_L g14758 ( 
.A(n_14613),
.Y(n_14758)
);

INVx2_ASAP7_75t_L g14759 ( 
.A(n_14516),
.Y(n_14759)
);

OAI22xp5_ASAP7_75t_L g14760 ( 
.A1(n_14332),
.A2(n_2298),
.B1(n_2296),
.B2(n_2297),
.Y(n_14760)
);

INVx3_ASAP7_75t_L g14761 ( 
.A(n_14473),
.Y(n_14761)
);

INVx2_ASAP7_75t_L g14762 ( 
.A(n_14544),
.Y(n_14762)
);

NAND2xp5_ASAP7_75t_L g14763 ( 
.A(n_14460),
.B(n_2297),
.Y(n_14763)
);

INVx1_ASAP7_75t_L g14764 ( 
.A(n_14430),
.Y(n_14764)
);

INVx2_ASAP7_75t_L g14765 ( 
.A(n_14324),
.Y(n_14765)
);

INVx1_ASAP7_75t_L g14766 ( 
.A(n_14456),
.Y(n_14766)
);

INVx3_ASAP7_75t_L g14767 ( 
.A(n_14601),
.Y(n_14767)
);

OR2x2_ASAP7_75t_L g14768 ( 
.A(n_14287),
.B(n_2298),
.Y(n_14768)
);

NAND2xp5_ASAP7_75t_SL g14769 ( 
.A(n_14633),
.B(n_2299),
.Y(n_14769)
);

INVx2_ASAP7_75t_L g14770 ( 
.A(n_14278),
.Y(n_14770)
);

INVx2_ASAP7_75t_L g14771 ( 
.A(n_14623),
.Y(n_14771)
);

HB1xp67_ASAP7_75t_L g14772 ( 
.A(n_14292),
.Y(n_14772)
);

INVx4_ASAP7_75t_L g14773 ( 
.A(n_14453),
.Y(n_14773)
);

INVx1_ASAP7_75t_L g14774 ( 
.A(n_14471),
.Y(n_14774)
);

INVx1_ASAP7_75t_L g14775 ( 
.A(n_14560),
.Y(n_14775)
);

INVx1_ASAP7_75t_L g14776 ( 
.A(n_14525),
.Y(n_14776)
);

INVx2_ASAP7_75t_SL g14777 ( 
.A(n_14585),
.Y(n_14777)
);

INVx1_ASAP7_75t_L g14778 ( 
.A(n_14448),
.Y(n_14778)
);

NAND2x1p5_ASAP7_75t_L g14779 ( 
.A(n_14290),
.B(n_2300),
.Y(n_14779)
);

A2O1A1Ixp33_ASAP7_75t_SL g14780 ( 
.A1(n_14536),
.A2(n_2302),
.B(n_2300),
.C(n_2301),
.Y(n_14780)
);

AO21x2_ASAP7_75t_L g14781 ( 
.A1(n_14416),
.A2(n_2301),
.B(n_2302),
.Y(n_14781)
);

INVx1_ASAP7_75t_L g14782 ( 
.A(n_14392),
.Y(n_14782)
);

INVx1_ASAP7_75t_L g14783 ( 
.A(n_14398),
.Y(n_14783)
);

HB1xp67_ASAP7_75t_L g14784 ( 
.A(n_14477),
.Y(n_14784)
);

INVx1_ASAP7_75t_L g14785 ( 
.A(n_14521),
.Y(n_14785)
);

NAND2xp5_ASAP7_75t_L g14786 ( 
.A(n_14647),
.B(n_2303),
.Y(n_14786)
);

AO32x2_ASAP7_75t_L g14787 ( 
.A1(n_14570),
.A2(n_2305),
.A3(n_2303),
.B1(n_2304),
.B2(n_2306),
.Y(n_14787)
);

AND2x4_ASAP7_75t_L g14788 ( 
.A(n_14615),
.B(n_2305),
.Y(n_14788)
);

INVx1_ASAP7_75t_L g14789 ( 
.A(n_14577),
.Y(n_14789)
);

INVx2_ASAP7_75t_L g14790 ( 
.A(n_14623),
.Y(n_14790)
);

HB1xp67_ASAP7_75t_L g14791 ( 
.A(n_14338),
.Y(n_14791)
);

INVx1_ASAP7_75t_L g14792 ( 
.A(n_14463),
.Y(n_14792)
);

INVx1_ASAP7_75t_L g14793 ( 
.A(n_14468),
.Y(n_14793)
);

INVx2_ASAP7_75t_L g14794 ( 
.A(n_14326),
.Y(n_14794)
);

OAI21x1_ASAP7_75t_L g14795 ( 
.A1(n_14325),
.A2(n_14277),
.B(n_14503),
.Y(n_14795)
);

INVx1_ASAP7_75t_L g14796 ( 
.A(n_14470),
.Y(n_14796)
);

OAI21xp5_ASAP7_75t_L g14797 ( 
.A1(n_14357),
.A2(n_2306),
.B(n_2307),
.Y(n_14797)
);

INVx1_ASAP7_75t_L g14798 ( 
.A(n_14361),
.Y(n_14798)
);

AND2x2_ASAP7_75t_L g14799 ( 
.A(n_14295),
.B(n_2307),
.Y(n_14799)
);

INVx1_ASAP7_75t_L g14800 ( 
.A(n_14368),
.Y(n_14800)
);

INVx2_ASAP7_75t_L g14801 ( 
.A(n_14276),
.Y(n_14801)
);

INVx2_ASAP7_75t_L g14802 ( 
.A(n_14371),
.Y(n_14802)
);

INVx1_ASAP7_75t_L g14803 ( 
.A(n_14379),
.Y(n_14803)
);

INVx1_ASAP7_75t_L g14804 ( 
.A(n_14387),
.Y(n_14804)
);

NAND2xp5_ASAP7_75t_L g14805 ( 
.A(n_14641),
.B(n_2308),
.Y(n_14805)
);

INVx1_ASAP7_75t_L g14806 ( 
.A(n_14437),
.Y(n_14806)
);

INVx1_ASAP7_75t_L g14807 ( 
.A(n_14447),
.Y(n_14807)
);

INVx1_ASAP7_75t_L g14808 ( 
.A(n_14451),
.Y(n_14808)
);

INVx2_ASAP7_75t_L g14809 ( 
.A(n_14579),
.Y(n_14809)
);

INVx1_ASAP7_75t_L g14810 ( 
.A(n_14604),
.Y(n_14810)
);

INVx1_ASAP7_75t_L g14811 ( 
.A(n_14366),
.Y(n_14811)
);

INVx2_ASAP7_75t_L g14812 ( 
.A(n_14585),
.Y(n_14812)
);

INVx1_ASAP7_75t_L g14813 ( 
.A(n_14482),
.Y(n_14813)
);

AND2x4_ASAP7_75t_L g14814 ( 
.A(n_14583),
.B(n_2308),
.Y(n_14814)
);

INVx1_ASAP7_75t_L g14815 ( 
.A(n_14380),
.Y(n_14815)
);

INVx2_ASAP7_75t_L g14816 ( 
.A(n_14331),
.Y(n_14816)
);

BUFx3_ASAP7_75t_L g14817 ( 
.A(n_14390),
.Y(n_14817)
);

OR2x6_ASAP7_75t_L g14818 ( 
.A(n_14395),
.B(n_14408),
.Y(n_14818)
);

INVx1_ASAP7_75t_L g14819 ( 
.A(n_14445),
.Y(n_14819)
);

NAND2xp5_ASAP7_75t_L g14820 ( 
.A(n_14370),
.B(n_14624),
.Y(n_14820)
);

AOI211xp5_ASAP7_75t_L g14821 ( 
.A1(n_14342),
.A2(n_2311),
.B(n_2309),
.C(n_2310),
.Y(n_14821)
);

INVx2_ASAP7_75t_L g14822 ( 
.A(n_14573),
.Y(n_14822)
);

INVx1_ASAP7_75t_L g14823 ( 
.A(n_14637),
.Y(n_14823)
);

OAI22xp5_ASAP7_75t_L g14824 ( 
.A1(n_14359),
.A2(n_2312),
.B1(n_2310),
.B2(n_2311),
.Y(n_14824)
);

INVx1_ASAP7_75t_L g14825 ( 
.A(n_14345),
.Y(n_14825)
);

INVx1_ASAP7_75t_L g14826 ( 
.A(n_14346),
.Y(n_14826)
);

OAI21x1_ASAP7_75t_L g14827 ( 
.A1(n_14505),
.A2(n_2312),
.B(n_2313),
.Y(n_14827)
);

INVx2_ASAP7_75t_L g14828 ( 
.A(n_14563),
.Y(n_14828)
);

OR2x2_ASAP7_75t_L g14829 ( 
.A(n_14304),
.B(n_2313),
.Y(n_14829)
);

HB1xp67_ASAP7_75t_L g14830 ( 
.A(n_14512),
.Y(n_14830)
);

INVx1_ASAP7_75t_L g14831 ( 
.A(n_14494),
.Y(n_14831)
);

INVx1_ASAP7_75t_L g14832 ( 
.A(n_14506),
.Y(n_14832)
);

INVx3_ASAP7_75t_L g14833 ( 
.A(n_14486),
.Y(n_14833)
);

OAI21x1_ASAP7_75t_L g14834 ( 
.A1(n_14458),
.A2(n_2314),
.B(n_2315),
.Y(n_14834)
);

INVx1_ASAP7_75t_L g14835 ( 
.A(n_14507),
.Y(n_14835)
);

AND2x2_ASAP7_75t_L g14836 ( 
.A(n_14308),
.B(n_2314),
.Y(n_14836)
);

INVx1_ASAP7_75t_L g14837 ( 
.A(n_14519),
.Y(n_14837)
);

AOI21x1_ASAP7_75t_L g14838 ( 
.A1(n_14397),
.A2(n_2315),
.B(n_2316),
.Y(n_14838)
);

CKINVDCx20_ASAP7_75t_R g14839 ( 
.A(n_14598),
.Y(n_14839)
);

OAI21x1_ASAP7_75t_L g14840 ( 
.A1(n_14330),
.A2(n_2317),
.B(n_2318),
.Y(n_14840)
);

INVx1_ASAP7_75t_L g14841 ( 
.A(n_14545),
.Y(n_14841)
);

INVx1_ASAP7_75t_L g14842 ( 
.A(n_14547),
.Y(n_14842)
);

INVx2_ASAP7_75t_L g14843 ( 
.A(n_14651),
.Y(n_14843)
);

AND2x2_ASAP7_75t_L g14844 ( 
.A(n_14582),
.B(n_2318),
.Y(n_14844)
);

INVx2_ASAP7_75t_L g14845 ( 
.A(n_14658),
.Y(n_14845)
);

INVx2_ASAP7_75t_L g14846 ( 
.A(n_14518),
.Y(n_14846)
);

OAI21x1_ASAP7_75t_L g14847 ( 
.A1(n_14335),
.A2(n_2319),
.B(n_2320),
.Y(n_14847)
);

AO21x2_ASAP7_75t_L g14848 ( 
.A1(n_14293),
.A2(n_2319),
.B(n_2320),
.Y(n_14848)
);

INVx1_ASAP7_75t_L g14849 ( 
.A(n_14564),
.Y(n_14849)
);

INVx2_ASAP7_75t_L g14850 ( 
.A(n_14633),
.Y(n_14850)
);

INVx1_ASAP7_75t_L g14851 ( 
.A(n_14509),
.Y(n_14851)
);

INVx2_ASAP7_75t_L g14852 ( 
.A(n_14497),
.Y(n_14852)
);

INVx2_ASAP7_75t_L g14853 ( 
.A(n_14553),
.Y(n_14853)
);

OAI21x1_ASAP7_75t_L g14854 ( 
.A1(n_14302),
.A2(n_2321),
.B(n_2322),
.Y(n_14854)
);

INVx2_ASAP7_75t_L g14855 ( 
.A(n_14648),
.Y(n_14855)
);

INVx1_ASAP7_75t_L g14856 ( 
.A(n_14393),
.Y(n_14856)
);

AO21x2_ASAP7_75t_L g14857 ( 
.A1(n_14593),
.A2(n_2322),
.B(n_2323),
.Y(n_14857)
);

INVx1_ASAP7_75t_L g14858 ( 
.A(n_14344),
.Y(n_14858)
);

A2O1A1Ixp33_ASAP7_75t_SL g14859 ( 
.A1(n_14602),
.A2(n_2325),
.B(n_2323),
.C(n_2324),
.Y(n_14859)
);

INVx2_ASAP7_75t_L g14860 ( 
.A(n_14650),
.Y(n_14860)
);

OR2x2_ASAP7_75t_L g14861 ( 
.A(n_14391),
.B(n_14586),
.Y(n_14861)
);

INVx2_ASAP7_75t_L g14862 ( 
.A(n_14656),
.Y(n_14862)
);

AND2x2_ASAP7_75t_L g14863 ( 
.A(n_14305),
.B(n_2324),
.Y(n_14863)
);

INVx3_ASAP7_75t_L g14864 ( 
.A(n_14491),
.Y(n_14864)
);

INVx2_ASAP7_75t_L g14865 ( 
.A(n_14303),
.Y(n_14865)
);

INVx1_ASAP7_75t_L g14866 ( 
.A(n_14662),
.Y(n_14866)
);

INVx2_ASAP7_75t_SL g14867 ( 
.A(n_14405),
.Y(n_14867)
);

OAI21x1_ASAP7_75t_L g14868 ( 
.A1(n_14358),
.A2(n_2326),
.B(n_2327),
.Y(n_14868)
);

INVx2_ASAP7_75t_SL g14869 ( 
.A(n_14513),
.Y(n_14869)
);

HB1xp67_ASAP7_75t_L g14870 ( 
.A(n_14508),
.Y(n_14870)
);

INVx1_ASAP7_75t_L g14871 ( 
.A(n_14377),
.Y(n_14871)
);

INVx1_ASAP7_75t_L g14872 ( 
.A(n_14403),
.Y(n_14872)
);

INVx2_ASAP7_75t_L g14873 ( 
.A(n_14638),
.Y(n_14873)
);

AND2x2_ASAP7_75t_L g14874 ( 
.A(n_14310),
.B(n_2326),
.Y(n_14874)
);

INVx2_ASAP7_75t_SL g14875 ( 
.A(n_14435),
.Y(n_14875)
);

AND2x4_ASAP7_75t_L g14876 ( 
.A(n_14383),
.B(n_2328),
.Y(n_14876)
);

OAI21x1_ASAP7_75t_L g14877 ( 
.A1(n_14297),
.A2(n_2328),
.B(n_2329),
.Y(n_14877)
);

INVx4_ASAP7_75t_L g14878 ( 
.A(n_14480),
.Y(n_14878)
);

INVx1_ASAP7_75t_L g14879 ( 
.A(n_14424),
.Y(n_14879)
);

INVx1_ASAP7_75t_L g14880 ( 
.A(n_14611),
.Y(n_14880)
);

INVx2_ASAP7_75t_L g14881 ( 
.A(n_14301),
.Y(n_14881)
);

INVx1_ASAP7_75t_L g14882 ( 
.A(n_14568),
.Y(n_14882)
);

INVxp67_ASAP7_75t_SL g14883 ( 
.A(n_14428),
.Y(n_14883)
);

INVx1_ASAP7_75t_L g14884 ( 
.A(n_14531),
.Y(n_14884)
);

OAI21x1_ASAP7_75t_L g14885 ( 
.A1(n_14319),
.A2(n_2329),
.B(n_2330),
.Y(n_14885)
);

OAI22xp5_ASAP7_75t_L g14886 ( 
.A1(n_14485),
.A2(n_2332),
.B1(n_2330),
.B2(n_2331),
.Y(n_14886)
);

AO21x2_ASAP7_75t_L g14887 ( 
.A1(n_14596),
.A2(n_2331),
.B(n_2332),
.Y(n_14887)
);

AND2x2_ASAP7_75t_L g14888 ( 
.A(n_14562),
.B(n_2333),
.Y(n_14888)
);

OA21x2_ASAP7_75t_L g14889 ( 
.A1(n_14461),
.A2(n_2333),
.B(n_2334),
.Y(n_14889)
);

OAI221xp5_ASAP7_75t_L g14890 ( 
.A1(n_14355),
.A2(n_2336),
.B1(n_2334),
.B2(n_2335),
.C(n_2337),
.Y(n_14890)
);

BUFx3_ASAP7_75t_L g14891 ( 
.A(n_14429),
.Y(n_14891)
);

INVx1_ASAP7_75t_L g14892 ( 
.A(n_14541),
.Y(n_14892)
);

INVx1_ASAP7_75t_L g14893 ( 
.A(n_14542),
.Y(n_14893)
);

INVx1_ASAP7_75t_L g14894 ( 
.A(n_14496),
.Y(n_14894)
);

OA21x2_ASAP7_75t_L g14895 ( 
.A1(n_14350),
.A2(n_2335),
.B(n_2336),
.Y(n_14895)
);

BUFx6f_ASAP7_75t_L g14896 ( 
.A(n_14548),
.Y(n_14896)
);

INVx1_ASAP7_75t_L g14897 ( 
.A(n_14459),
.Y(n_14897)
);

BUFx3_ASAP7_75t_L g14898 ( 
.A(n_14479),
.Y(n_14898)
);

OR2x2_ASAP7_75t_L g14899 ( 
.A(n_14421),
.B(n_2337),
.Y(n_14899)
);

INVx1_ASAP7_75t_L g14900 ( 
.A(n_14414),
.Y(n_14900)
);

INVx2_ASAP7_75t_L g14901 ( 
.A(n_14472),
.Y(n_14901)
);

NAND2x1_ASAP7_75t_L g14902 ( 
.A(n_14550),
.B(n_2338),
.Y(n_14902)
);

HB1xp67_ASAP7_75t_L g14903 ( 
.A(n_14340),
.Y(n_14903)
);

AND2x2_ASAP7_75t_L g14904 ( 
.A(n_14415),
.B(n_2339),
.Y(n_14904)
);

INVx1_ASAP7_75t_L g14905 ( 
.A(n_14439),
.Y(n_14905)
);

INVx1_ASAP7_75t_SL g14906 ( 
.A(n_14476),
.Y(n_14906)
);

AND2x2_ASAP7_75t_L g14907 ( 
.A(n_14396),
.B(n_2340),
.Y(n_14907)
);

INVx2_ASAP7_75t_L g14908 ( 
.A(n_14483),
.Y(n_14908)
);

BUFx2_ASAP7_75t_L g14909 ( 
.A(n_14594),
.Y(n_14909)
);

INVx1_ASAP7_75t_L g14910 ( 
.A(n_14605),
.Y(n_14910)
);

INVx2_ASAP7_75t_L g14911 ( 
.A(n_14418),
.Y(n_14911)
);

HB1xp67_ASAP7_75t_L g14912 ( 
.A(n_14627),
.Y(n_14912)
);

BUFx6f_ASAP7_75t_SL g14913 ( 
.A(n_14594),
.Y(n_14913)
);

INVx3_ASAP7_75t_L g14914 ( 
.A(n_14635),
.Y(n_14914)
);

BUFx2_ASAP7_75t_L g14915 ( 
.A(n_14449),
.Y(n_14915)
);

BUFx3_ASAP7_75t_L g14916 ( 
.A(n_14554),
.Y(n_14916)
);

INVx1_ASAP7_75t_L g14917 ( 
.A(n_14606),
.Y(n_14917)
);

OR2x2_ASAP7_75t_L g14918 ( 
.A(n_14373),
.B(n_2340),
.Y(n_14918)
);

OA21x2_ASAP7_75t_L g14919 ( 
.A1(n_14402),
.A2(n_2341),
.B(n_2342),
.Y(n_14919)
);

OA21x2_ASAP7_75t_L g14920 ( 
.A1(n_14444),
.A2(n_14614),
.B(n_14328),
.Y(n_14920)
);

OA21x2_ASAP7_75t_L g14921 ( 
.A1(n_14404),
.A2(n_2341),
.B(n_2342),
.Y(n_14921)
);

INVx2_ASAP7_75t_L g14922 ( 
.A(n_14382),
.Y(n_14922)
);

INVx2_ASAP7_75t_L g14923 ( 
.A(n_14502),
.Y(n_14923)
);

INVx2_ASAP7_75t_L g14924 ( 
.A(n_14481),
.Y(n_14924)
);

INVx3_ASAP7_75t_L g14925 ( 
.A(n_14555),
.Y(n_14925)
);

BUFx2_ASAP7_75t_L g14926 ( 
.A(n_14649),
.Y(n_14926)
);

INVx2_ASAP7_75t_L g14927 ( 
.A(n_14484),
.Y(n_14927)
);

NAND2xp5_ASAP7_75t_L g14928 ( 
.A(n_14625),
.B(n_2343),
.Y(n_14928)
);

BUFx3_ASAP7_75t_L g14929 ( 
.A(n_14556),
.Y(n_14929)
);

AND2x2_ASAP7_75t_L g14930 ( 
.A(n_14420),
.B(n_2343),
.Y(n_14930)
);

BUFx2_ASAP7_75t_L g14931 ( 
.A(n_14654),
.Y(n_14931)
);

CKINVDCx20_ASAP7_75t_R g14932 ( 
.A(n_14626),
.Y(n_14932)
);

INVx2_ASAP7_75t_L g14933 ( 
.A(n_14489),
.Y(n_14933)
);

INVx2_ASAP7_75t_SL g14934 ( 
.A(n_14526),
.Y(n_14934)
);

INVx1_ASAP7_75t_L g14935 ( 
.A(n_14492),
.Y(n_14935)
);

INVx1_ASAP7_75t_L g14936 ( 
.A(n_14469),
.Y(n_14936)
);

AOI22xp33_ASAP7_75t_L g14937 ( 
.A1(n_14369),
.A2(n_2346),
.B1(n_2344),
.B2(n_2345),
.Y(n_14937)
);

NAND2x1p5_ASAP7_75t_L g14938 ( 
.A(n_14446),
.B(n_2344),
.Y(n_14938)
);

INVx1_ASAP7_75t_L g14939 ( 
.A(n_14609),
.Y(n_14939)
);

OAI21x1_ASAP7_75t_L g14940 ( 
.A1(n_14285),
.A2(n_2345),
.B(n_2346),
.Y(n_14940)
);

HB1xp67_ASAP7_75t_L g14941 ( 
.A(n_14289),
.Y(n_14941)
);

INVx1_ASAP7_75t_L g14942 ( 
.A(n_14436),
.Y(n_14942)
);

INVx1_ASAP7_75t_L g14943 ( 
.A(n_14400),
.Y(n_14943)
);

INVx2_ASAP7_75t_L g14944 ( 
.A(n_14532),
.Y(n_14944)
);

INVx1_ASAP7_75t_L g14945 ( 
.A(n_14631),
.Y(n_14945)
);

INVx1_ASAP7_75t_L g14946 ( 
.A(n_14632),
.Y(n_14946)
);

INVx2_ASAP7_75t_L g14947 ( 
.A(n_14645),
.Y(n_14947)
);

INVx3_ASAP7_75t_L g14948 ( 
.A(n_14569),
.Y(n_14948)
);

INVx4_ASAP7_75t_L g14949 ( 
.A(n_14559),
.Y(n_14949)
);

AO21x1_ASAP7_75t_L g14950 ( 
.A1(n_14425),
.A2(n_2347),
.B(n_2348),
.Y(n_14950)
);

INVx2_ASAP7_75t_SL g14951 ( 
.A(n_14610),
.Y(n_14951)
);

INVx1_ASAP7_75t_L g14952 ( 
.A(n_14465),
.Y(n_14952)
);

BUFx3_ASAP7_75t_L g14953 ( 
.A(n_14618),
.Y(n_14953)
);

INVx3_ASAP7_75t_L g14954 ( 
.A(n_14566),
.Y(n_14954)
);

INVx1_ASAP7_75t_L g14955 ( 
.A(n_14466),
.Y(n_14955)
);

INVx1_ASAP7_75t_L g14956 ( 
.A(n_14534),
.Y(n_14956)
);

INVx3_ASAP7_75t_L g14957 ( 
.A(n_14629),
.Y(n_14957)
);

BUFx3_ASAP7_75t_L g14958 ( 
.A(n_14580),
.Y(n_14958)
);

INVx1_ASAP7_75t_L g14959 ( 
.A(n_14517),
.Y(n_14959)
);

AO21x2_ASAP7_75t_L g14960 ( 
.A1(n_14621),
.A2(n_2347),
.B(n_2348),
.Y(n_14960)
);

AND2x2_ASAP7_75t_L g14961 ( 
.A(n_14314),
.B(n_2349),
.Y(n_14961)
);

BUFx6f_ASAP7_75t_L g14962 ( 
.A(n_14581),
.Y(n_14962)
);

OA21x2_ASAP7_75t_L g14963 ( 
.A1(n_14318),
.A2(n_2349),
.B(n_2350),
.Y(n_14963)
);

INVx1_ASAP7_75t_L g14964 ( 
.A(n_14527),
.Y(n_14964)
);

INVx2_ASAP7_75t_L g14965 ( 
.A(n_14565),
.Y(n_14965)
);

INVx1_ASAP7_75t_L g14966 ( 
.A(n_14612),
.Y(n_14966)
);

INVx1_ASAP7_75t_L g14967 ( 
.A(n_14642),
.Y(n_14967)
);

OAI21xp5_ASAP7_75t_L g14968 ( 
.A1(n_14539),
.A2(n_2350),
.B(n_2351),
.Y(n_14968)
);

AND2x2_ASAP7_75t_L g14969 ( 
.A(n_14576),
.B(n_2351),
.Y(n_14969)
);

AO21x2_ASAP7_75t_L g14970 ( 
.A1(n_14538),
.A2(n_2352),
.B(n_2353),
.Y(n_14970)
);

INVx1_ASAP7_75t_L g14971 ( 
.A(n_14630),
.Y(n_14971)
);

INVx2_ASAP7_75t_L g14972 ( 
.A(n_14591),
.Y(n_14972)
);

INVx1_ASAP7_75t_L g14973 ( 
.A(n_14652),
.Y(n_14973)
);

HB1xp67_ASAP7_75t_L g14974 ( 
.A(n_14616),
.Y(n_14974)
);

INVx3_ASAP7_75t_L g14975 ( 
.A(n_14578),
.Y(n_14975)
);

NAND2xp5_ASAP7_75t_L g14976 ( 
.A(n_14433),
.B(n_2354),
.Y(n_14976)
);

INVx1_ASAP7_75t_SL g14977 ( 
.A(n_14646),
.Y(n_14977)
);

BUFx2_ASAP7_75t_L g14978 ( 
.A(n_14607),
.Y(n_14978)
);

BUFx3_ASAP7_75t_L g14979 ( 
.A(n_14417),
.Y(n_14979)
);

AOI21xp5_ASAP7_75t_L g14980 ( 
.A1(n_14288),
.A2(n_2354),
.B(n_2355),
.Y(n_14980)
);

NAND2xp5_ASAP7_75t_L g14981 ( 
.A(n_14661),
.B(n_2356),
.Y(n_14981)
);

INVx1_ASAP7_75t_L g14982 ( 
.A(n_14406),
.Y(n_14982)
);

CKINVDCx5p33_ASAP7_75t_R g14983 ( 
.A(n_14636),
.Y(n_14983)
);

INVx1_ASAP7_75t_L g14984 ( 
.A(n_14589),
.Y(n_14984)
);

INVx1_ASAP7_75t_L g14985 ( 
.A(n_14660),
.Y(n_14985)
);

INVx2_ASAP7_75t_L g14986 ( 
.A(n_14603),
.Y(n_14986)
);

INVx2_ASAP7_75t_L g14987 ( 
.A(n_14659),
.Y(n_14987)
);

INVx3_ASAP7_75t_L g14988 ( 
.A(n_14474),
.Y(n_14988)
);

CKINVDCx11_ASAP7_75t_R g14989 ( 
.A(n_14487),
.Y(n_14989)
);

INVx1_ASAP7_75t_L g14990 ( 
.A(n_14546),
.Y(n_14990)
);

HB1xp67_ASAP7_75t_L g14991 ( 
.A(n_14634),
.Y(n_14991)
);

INVx2_ASAP7_75t_L g14992 ( 
.A(n_14528),
.Y(n_14992)
);

INVx3_ASAP7_75t_L g14993 ( 
.A(n_14620),
.Y(n_14993)
);

INVx2_ASAP7_75t_L g14994 ( 
.A(n_14533),
.Y(n_14994)
);

INVx2_ASAP7_75t_L g14995 ( 
.A(n_14389),
.Y(n_14995)
);

OAI21xp5_ASAP7_75t_L g14996 ( 
.A1(n_14571),
.A2(n_14450),
.B(n_14529),
.Y(n_14996)
);

AND2x4_ASAP7_75t_L g14997 ( 
.A(n_14364),
.B(n_2357),
.Y(n_14997)
);

INVx1_ASAP7_75t_L g14998 ( 
.A(n_14495),
.Y(n_14998)
);

AND2x2_ASAP7_75t_L g14999 ( 
.A(n_14639),
.B(n_2357),
.Y(n_14999)
);

OAI21x1_ASAP7_75t_L g15000 ( 
.A1(n_14334),
.A2(n_2358),
.B(n_2359),
.Y(n_15000)
);

OAI21xp5_ASAP7_75t_L g15001 ( 
.A1(n_14296),
.A2(n_2358),
.B(n_2359),
.Y(n_15001)
);

INVx1_ASAP7_75t_L g15002 ( 
.A(n_14500),
.Y(n_15002)
);

INVx2_ASAP7_75t_L g15003 ( 
.A(n_14597),
.Y(n_15003)
);

INVx1_ASAP7_75t_L g15004 ( 
.A(n_14504),
.Y(n_15004)
);

INVx2_ASAP7_75t_SL g15005 ( 
.A(n_14595),
.Y(n_15005)
);

HB1xp67_ASAP7_75t_L g15006 ( 
.A(n_14588),
.Y(n_15006)
);

INVx1_ASAP7_75t_L g15007 ( 
.A(n_14514),
.Y(n_15007)
);

INVx2_ASAP7_75t_L g15008 ( 
.A(n_14394),
.Y(n_15008)
);

HB1xp67_ASAP7_75t_L g15009 ( 
.A(n_14643),
.Y(n_15009)
);

INVx2_ASAP7_75t_L g15010 ( 
.A(n_14498),
.Y(n_15010)
);

HB1xp67_ASAP7_75t_L g15011 ( 
.A(n_14351),
.Y(n_15011)
);

HB1xp67_ASAP7_75t_L g15012 ( 
.A(n_14365),
.Y(n_15012)
);

INVx1_ASAP7_75t_L g15013 ( 
.A(n_14653),
.Y(n_15013)
);

HB1xp67_ASAP7_75t_L g15014 ( 
.A(n_14452),
.Y(n_15014)
);

HB1xp67_ASAP7_75t_L g15015 ( 
.A(n_14655),
.Y(n_15015)
);

AND2x2_ASAP7_75t_L g15016 ( 
.A(n_14640),
.B(n_2360),
.Y(n_15016)
);

BUFx3_ASAP7_75t_L g15017 ( 
.A(n_14644),
.Y(n_15017)
);

AO21x2_ASAP7_75t_L g15018 ( 
.A1(n_14619),
.A2(n_2361),
.B(n_2362),
.Y(n_15018)
);

INVx1_ASAP7_75t_L g15019 ( 
.A(n_14663),
.Y(n_15019)
);

INVx3_ASAP7_75t_L g15020 ( 
.A(n_14347),
.Y(n_15020)
);

INVx2_ASAP7_75t_SL g15021 ( 
.A(n_14574),
.Y(n_15021)
);

INVx3_ASAP7_75t_L g15022 ( 
.A(n_14317),
.Y(n_15022)
);

AO21x2_ASAP7_75t_L g15023 ( 
.A1(n_14423),
.A2(n_2362),
.B(n_2363),
.Y(n_15023)
);

INVx2_ASAP7_75t_L g15024 ( 
.A(n_14427),
.Y(n_15024)
);

NOR3xp33_ASAP7_75t_SL g15025 ( 
.A(n_14890),
.B(n_14599),
.C(n_14522),
.Y(n_15025)
);

INVx2_ASAP7_75t_L g15026 ( 
.A(n_14679),
.Y(n_15026)
);

NAND2xp5_ASAP7_75t_L g15027 ( 
.A(n_14828),
.B(n_15012),
.Y(n_15027)
);

INVx8_ASAP7_75t_L g15028 ( 
.A(n_14754),
.Y(n_15028)
);

INVx1_ASAP7_75t_L g15029 ( 
.A(n_14704),
.Y(n_15029)
);

INVx3_ASAP7_75t_L g15030 ( 
.A(n_14680),
.Y(n_15030)
);

CKINVDCx20_ASAP7_75t_R g15031 ( 
.A(n_14746),
.Y(n_15031)
);

INVx2_ASAP7_75t_L g15032 ( 
.A(n_14691),
.Y(n_15032)
);

NAND2xp5_ASAP7_75t_L g15033 ( 
.A(n_15019),
.B(n_14657),
.Y(n_15033)
);

INVx1_ASAP7_75t_L g15034 ( 
.A(n_14749),
.Y(n_15034)
);

OR2x6_ASAP7_75t_L g15035 ( 
.A(n_14744),
.B(n_14381),
.Y(n_15035)
);

NOR2xp33_ASAP7_75t_L g15036 ( 
.A(n_14717),
.B(n_14316),
.Y(n_15036)
);

AND2x2_ASAP7_75t_L g15037 ( 
.A(n_14761),
.B(n_14524),
.Y(n_15037)
);

AND2x2_ASAP7_75t_L g15038 ( 
.A(n_14758),
.B(n_14362),
.Y(n_15038)
);

INVx1_ASAP7_75t_L g15039 ( 
.A(n_14672),
.Y(n_15039)
);

HB1xp67_ASAP7_75t_L g15040 ( 
.A(n_14751),
.Y(n_15040)
);

HB1xp67_ASAP7_75t_L g15041 ( 
.A(n_14830),
.Y(n_15041)
);

NAND2xp5_ASAP7_75t_SL g15042 ( 
.A(n_15022),
.B(n_14378),
.Y(n_15042)
);

CKINVDCx5p33_ASAP7_75t_R g15043 ( 
.A(n_14697),
.Y(n_15043)
);

INVx2_ASAP7_75t_L g15044 ( 
.A(n_14692),
.Y(n_15044)
);

CKINVDCx16_ASAP7_75t_R g15045 ( 
.A(n_14839),
.Y(n_15045)
);

HB1xp67_ASAP7_75t_L g15046 ( 
.A(n_14684),
.Y(n_15046)
);

OR2x2_ASAP7_75t_L g15047 ( 
.A(n_14669),
.B(n_14298),
.Y(n_15047)
);

OR2x6_ASAP7_75t_L g15048 ( 
.A(n_14744),
.B(n_14478),
.Y(n_15048)
);

CKINVDCx5p33_ASAP7_75t_R g15049 ( 
.A(n_14983),
.Y(n_15049)
);

INVx2_ASAP7_75t_L g15050 ( 
.A(n_14688),
.Y(n_15050)
);

HB1xp67_ASAP7_75t_L g15051 ( 
.A(n_14978),
.Y(n_15051)
);

INVx1_ASAP7_75t_L g15052 ( 
.A(n_14810),
.Y(n_15052)
);

NOR2xp33_ASAP7_75t_R g15053 ( 
.A(n_14932),
.B(n_2363),
.Y(n_15053)
);

INVx2_ASAP7_75t_L g15054 ( 
.A(n_14708),
.Y(n_15054)
);

AO32x2_ASAP7_75t_L g15055 ( 
.A1(n_14687),
.A2(n_14499),
.A3(n_14313),
.B1(n_14443),
.B2(n_14467),
.Y(n_15055)
);

OR2x6_ASAP7_75t_L g15056 ( 
.A(n_14734),
.B(n_14818),
.Y(n_15056)
);

CKINVDCx16_ASAP7_75t_R g15057 ( 
.A(n_14913),
.Y(n_15057)
);

BUFx3_ASAP7_75t_L g15058 ( 
.A(n_14898),
.Y(n_15058)
);

NAND2xp5_ASAP7_75t_L g15059 ( 
.A(n_14706),
.B(n_14422),
.Y(n_15059)
);

CKINVDCx5p33_ASAP7_75t_R g15060 ( 
.A(n_14729),
.Y(n_15060)
);

INVx1_ASAP7_75t_L g15061 ( 
.A(n_14664),
.Y(n_15061)
);

INVx1_ASAP7_75t_L g15062 ( 
.A(n_14666),
.Y(n_15062)
);

NOR3xp33_ASAP7_75t_SL g15063 ( 
.A(n_14820),
.B(n_14488),
.C(n_14432),
.Y(n_15063)
);

INVx1_ASAP7_75t_L g15064 ( 
.A(n_14670),
.Y(n_15064)
);

OR2x6_ASAP7_75t_L g15065 ( 
.A(n_14818),
.B(n_14434),
.Y(n_15065)
);

NAND2xp33_ASAP7_75t_R g15066 ( 
.A(n_14920),
.B(n_14575),
.Y(n_15066)
);

NOR3xp33_ASAP7_75t_SL g15067 ( 
.A(n_14726),
.B(n_14628),
.C(n_14413),
.Y(n_15067)
);

AND2x2_ASAP7_75t_L g15068 ( 
.A(n_14941),
.B(n_14590),
.Y(n_15068)
);

INVx2_ASAP7_75t_L g15069 ( 
.A(n_14674),
.Y(n_15069)
);

AND2x2_ASAP7_75t_L g15070 ( 
.A(n_14738),
.B(n_14600),
.Y(n_15070)
);

AOI22xp33_ASAP7_75t_SL g15071 ( 
.A1(n_15009),
.A2(n_14455),
.B1(n_14530),
.B2(n_2366),
.Y(n_15071)
);

HB1xp67_ASAP7_75t_L g15072 ( 
.A(n_14909),
.Y(n_15072)
);

INVx1_ASAP7_75t_L g15073 ( 
.A(n_14673),
.Y(n_15073)
);

NOR2xp33_ASAP7_75t_L g15074 ( 
.A(n_14914),
.B(n_2364),
.Y(n_15074)
);

INVx1_ASAP7_75t_L g15075 ( 
.A(n_14678),
.Y(n_15075)
);

INVx4_ASAP7_75t_L g15076 ( 
.A(n_14699),
.Y(n_15076)
);

INVx1_ASAP7_75t_L g15077 ( 
.A(n_14681),
.Y(n_15077)
);

INVx1_ASAP7_75t_L g15078 ( 
.A(n_14813),
.Y(n_15078)
);

AND2x2_ASAP7_75t_L g15079 ( 
.A(n_14677),
.B(n_2364),
.Y(n_15079)
);

INVx3_ASAP7_75t_L g15080 ( 
.A(n_14773),
.Y(n_15080)
);

BUFx6f_ASAP7_75t_L g15081 ( 
.A(n_14699),
.Y(n_15081)
);

INVx2_ASAP7_75t_L g15082 ( 
.A(n_14719),
.Y(n_15082)
);

AND2x2_ASAP7_75t_L g15083 ( 
.A(n_14695),
.B(n_2365),
.Y(n_15083)
);

INVx3_ASAP7_75t_L g15084 ( 
.A(n_14817),
.Y(n_15084)
);

HB1xp67_ASAP7_75t_L g15085 ( 
.A(n_14883),
.Y(n_15085)
);

AND2x4_ASAP7_75t_L g15086 ( 
.A(n_14716),
.B(n_2365),
.Y(n_15086)
);

AND2x2_ASAP7_75t_L g15087 ( 
.A(n_14665),
.B(n_2366),
.Y(n_15087)
);

AOI22xp33_ASAP7_75t_L g15088 ( 
.A1(n_15015),
.A2(n_2369),
.B1(n_2367),
.B2(n_2368),
.Y(n_15088)
);

AND2x2_ASAP7_75t_L g15089 ( 
.A(n_14730),
.B(n_2367),
.Y(n_15089)
);

AND2x4_ASAP7_75t_L g15090 ( 
.A(n_14733),
.B(n_2368),
.Y(n_15090)
);

BUFx6f_ASAP7_75t_L g15091 ( 
.A(n_14740),
.Y(n_15091)
);

AND2x2_ASAP7_75t_L g15092 ( 
.A(n_14767),
.B(n_2369),
.Y(n_15092)
);

BUFx6f_ASAP7_75t_L g15093 ( 
.A(n_14814),
.Y(n_15093)
);

AO31x2_ASAP7_75t_L g15094 ( 
.A1(n_14915),
.A2(n_2372),
.A3(n_2370),
.B(n_2371),
.Y(n_15094)
);

AND2x2_ASAP7_75t_L g15095 ( 
.A(n_14701),
.B(n_14949),
.Y(n_15095)
);

CKINVDCx16_ASAP7_75t_R g15096 ( 
.A(n_14977),
.Y(n_15096)
);

INVx3_ASAP7_75t_L g15097 ( 
.A(n_14891),
.Y(n_15097)
);

INVx2_ASAP7_75t_L g15098 ( 
.A(n_14719),
.Y(n_15098)
);

NOR2x1p5_ASAP7_75t_L g15099 ( 
.A(n_14902),
.B(n_2372),
.Y(n_15099)
);

OA21x2_ASAP7_75t_L g15100 ( 
.A1(n_14903),
.A2(n_2373),
.B(n_2374),
.Y(n_15100)
);

INVx1_ASAP7_75t_L g15101 ( 
.A(n_14939),
.Y(n_15101)
);

NAND2xp33_ASAP7_75t_SL g15102 ( 
.A(n_14747),
.B(n_2373),
.Y(n_15102)
);

AND2x2_ASAP7_75t_L g15103 ( 
.A(n_14702),
.B(n_2374),
.Y(n_15103)
);

INVx1_ASAP7_75t_L g15104 ( 
.A(n_14772),
.Y(n_15104)
);

INVx1_ASAP7_75t_L g15105 ( 
.A(n_14776),
.Y(n_15105)
);

BUFx6f_ASAP7_75t_L g15106 ( 
.A(n_14754),
.Y(n_15106)
);

INVx1_ASAP7_75t_L g15107 ( 
.A(n_14685),
.Y(n_15107)
);

HB1xp67_ASAP7_75t_L g15108 ( 
.A(n_14870),
.Y(n_15108)
);

INVx2_ASAP7_75t_L g15109 ( 
.A(n_14896),
.Y(n_15109)
);

OR2x6_ASAP7_75t_L g15110 ( 
.A(n_14980),
.B(n_2375),
.Y(n_15110)
);

BUFx3_ASAP7_75t_L g15111 ( 
.A(n_14938),
.Y(n_15111)
);

NAND2xp5_ASAP7_75t_L g15112 ( 
.A(n_15014),
.B(n_2375),
.Y(n_15112)
);

NAND2xp33_ASAP7_75t_SL g15113 ( 
.A(n_15006),
.B(n_2376),
.Y(n_15113)
);

NAND2x1p5_ASAP7_75t_L g15114 ( 
.A(n_14906),
.B(n_2377),
.Y(n_15114)
);

INVx2_ASAP7_75t_L g15115 ( 
.A(n_14896),
.Y(n_15115)
);

NAND2xp33_ASAP7_75t_R g15116 ( 
.A(n_14919),
.B(n_2377),
.Y(n_15116)
);

AO31x2_ASAP7_75t_L g15117 ( 
.A1(n_14760),
.A2(n_2380),
.A3(n_2378),
.B(n_2379),
.Y(n_15117)
);

NAND2xp5_ASAP7_75t_L g15118 ( 
.A(n_14982),
.B(n_2378),
.Y(n_15118)
);

AOI22xp33_ASAP7_75t_L g15119 ( 
.A1(n_14989),
.A2(n_2382),
.B1(n_2379),
.B2(n_2381),
.Y(n_15119)
);

OAI22xp5_ASAP7_75t_L g15120 ( 
.A1(n_14821),
.A2(n_2384),
.B1(n_2381),
.B2(n_2383),
.Y(n_15120)
);

OAI21xp5_ASAP7_75t_L g15121 ( 
.A1(n_14757),
.A2(n_2383),
.B(n_2384),
.Y(n_15121)
);

INVx2_ASAP7_75t_L g15122 ( 
.A(n_14694),
.Y(n_15122)
);

NAND2xp33_ASAP7_75t_R g15123 ( 
.A(n_14963),
.B(n_2385),
.Y(n_15123)
);

AND2x4_ASAP7_75t_L g15124 ( 
.A(n_14777),
.B(n_2386),
.Y(n_15124)
);

INVx2_ASAP7_75t_L g15125 ( 
.A(n_14962),
.Y(n_15125)
);

NOR2x1_ASAP7_75t_L g15126 ( 
.A(n_14781),
.B(n_2386),
.Y(n_15126)
);

NAND3xp33_ASAP7_75t_SL g15127 ( 
.A(n_14996),
.B(n_2387),
.C(n_2388),
.Y(n_15127)
);

INVxp33_ASAP7_75t_SL g15128 ( 
.A(n_14991),
.Y(n_15128)
);

OR2x2_ASAP7_75t_L g15129 ( 
.A(n_14957),
.B(n_2387),
.Y(n_15129)
);

INVx1_ASAP7_75t_L g15130 ( 
.A(n_14700),
.Y(n_15130)
);

INVx1_ASAP7_75t_L g15131 ( 
.A(n_14703),
.Y(n_15131)
);

AND2x4_ASAP7_75t_L g15132 ( 
.A(n_14916),
.B(n_2388),
.Y(n_15132)
);

NAND2xp33_ASAP7_75t_SL g15133 ( 
.A(n_15023),
.B(n_2389),
.Y(n_15133)
);

AO31x2_ASAP7_75t_L g15134 ( 
.A1(n_14785),
.A2(n_2392),
.A3(n_2390),
.B(n_2391),
.Y(n_15134)
);

INVx1_ASAP7_75t_L g15135 ( 
.A(n_14705),
.Y(n_15135)
);

AND2x2_ASAP7_75t_L g15136 ( 
.A(n_14926),
.B(n_2391),
.Y(n_15136)
);

HB1xp67_ASAP7_75t_L g15137 ( 
.A(n_14931),
.Y(n_15137)
);

INVx3_ASAP7_75t_L g15138 ( 
.A(n_14878),
.Y(n_15138)
);

INVx1_ASAP7_75t_L g15139 ( 
.A(n_14711),
.Y(n_15139)
);

OAI22xp5_ASAP7_75t_L g15140 ( 
.A1(n_14686),
.A2(n_14690),
.B1(n_14937),
.B2(n_14721),
.Y(n_15140)
);

INVx1_ASAP7_75t_L g15141 ( 
.A(n_14713),
.Y(n_15141)
);

AND2x2_ASAP7_75t_L g15142 ( 
.A(n_14954),
.B(n_2392),
.Y(n_15142)
);

AND2x2_ASAP7_75t_L g15143 ( 
.A(n_14683),
.B(n_2394),
.Y(n_15143)
);

BUFx3_ASAP7_75t_L g15144 ( 
.A(n_14754),
.Y(n_15144)
);

OR2x6_ASAP7_75t_L g15145 ( 
.A(n_15001),
.B(n_2394),
.Y(n_15145)
);

INVx2_ASAP7_75t_L g15146 ( 
.A(n_14962),
.Y(n_15146)
);

NAND2xp5_ASAP7_75t_L g15147 ( 
.A(n_14990),
.B(n_2395),
.Y(n_15147)
);

NOR2xp33_ASAP7_75t_R g15148 ( 
.A(n_14988),
.B(n_2395),
.Y(n_15148)
);

NAND2xp5_ASAP7_75t_L g15149 ( 
.A(n_14985),
.B(n_2396),
.Y(n_15149)
);

NAND2xp5_ASAP7_75t_L g15150 ( 
.A(n_14998),
.B(n_2396),
.Y(n_15150)
);

BUFx2_ASAP7_75t_L g15151 ( 
.A(n_14929),
.Y(n_15151)
);

INVx3_ASAP7_75t_L g15152 ( 
.A(n_14833),
.Y(n_15152)
);

OR2x2_ASAP7_75t_L g15153 ( 
.A(n_14752),
.B(n_2397),
.Y(n_15153)
);

INVx1_ASAP7_75t_L g15154 ( 
.A(n_14715),
.Y(n_15154)
);

AND2x4_ASAP7_75t_L g15155 ( 
.A(n_14812),
.B(n_2397),
.Y(n_15155)
);

NAND2xp33_ASAP7_75t_SL g15156 ( 
.A(n_14966),
.B(n_2398),
.Y(n_15156)
);

INVx2_ASAP7_75t_L g15157 ( 
.A(n_14953),
.Y(n_15157)
);

INVx1_ASAP7_75t_L g15158 ( 
.A(n_14718),
.Y(n_15158)
);

HB1xp67_ASAP7_75t_L g15159 ( 
.A(n_14948),
.Y(n_15159)
);

NAND2xp5_ASAP7_75t_L g15160 ( 
.A(n_15002),
.B(n_2398),
.Y(n_15160)
);

NAND2xp5_ASAP7_75t_L g15161 ( 
.A(n_15004),
.B(n_2399),
.Y(n_15161)
);

INVx2_ASAP7_75t_L g15162 ( 
.A(n_14864),
.Y(n_15162)
);

NAND2xp5_ASAP7_75t_L g15163 ( 
.A(n_15007),
.B(n_2400),
.Y(n_15163)
);

CKINVDCx5p33_ASAP7_75t_R g15164 ( 
.A(n_14979),
.Y(n_15164)
);

INVx2_ASAP7_75t_L g15165 ( 
.A(n_14958),
.Y(n_15165)
);

INVxp67_ASAP7_75t_L g15166 ( 
.A(n_14912),
.Y(n_15166)
);

NAND2xp5_ASAP7_75t_L g15167 ( 
.A(n_15011),
.B(n_2400),
.Y(n_15167)
);

INVx1_ASAP7_75t_L g15168 ( 
.A(n_14720),
.Y(n_15168)
);

AND2x4_ASAP7_75t_L g15169 ( 
.A(n_14845),
.B(n_2401),
.Y(n_15169)
);

INVx1_ASAP7_75t_L g15170 ( 
.A(n_14723),
.Y(n_15170)
);

NAND2xp33_ASAP7_75t_R g15171 ( 
.A(n_14921),
.B(n_2401),
.Y(n_15171)
);

INVx1_ASAP7_75t_L g15172 ( 
.A(n_14724),
.Y(n_15172)
);

NAND2xp5_ASAP7_75t_L g15173 ( 
.A(n_14967),
.B(n_2402),
.Y(n_15173)
);

INVx2_ASAP7_75t_L g15174 ( 
.A(n_14869),
.Y(n_15174)
);

CKINVDCx5p33_ASAP7_75t_R g15175 ( 
.A(n_14876),
.Y(n_15175)
);

HB1xp67_ASAP7_75t_L g15176 ( 
.A(n_14846),
.Y(n_15176)
);

INVx2_ASAP7_75t_L g15177 ( 
.A(n_14925),
.Y(n_15177)
);

AND2x4_ASAP7_75t_L g15178 ( 
.A(n_14707),
.B(n_2402),
.Y(n_15178)
);

AND2x2_ASAP7_75t_L g15179 ( 
.A(n_14689),
.B(n_2403),
.Y(n_15179)
);

INVxp67_ASAP7_75t_L g15180 ( 
.A(n_14686),
.Y(n_15180)
);

NAND2xp5_ASAP7_75t_L g15181 ( 
.A(n_15013),
.B(n_2403),
.Y(n_15181)
);

NAND2xp33_ASAP7_75t_R g15182 ( 
.A(n_14889),
.B(n_2404),
.Y(n_15182)
);

CKINVDCx5p33_ASAP7_75t_R g15183 ( 
.A(n_14961),
.Y(n_15183)
);

AND2x2_ASAP7_75t_L g15184 ( 
.A(n_14975),
.B(n_2404),
.Y(n_15184)
);

BUFx10_ASAP7_75t_L g15185 ( 
.A(n_14788),
.Y(n_15185)
);

CKINVDCx11_ASAP7_75t_R g15186 ( 
.A(n_14995),
.Y(n_15186)
);

AOI22xp33_ASAP7_75t_L g15187 ( 
.A1(n_15020),
.A2(n_2407),
.B1(n_2405),
.B2(n_2406),
.Y(n_15187)
);

NAND3xp33_ASAP7_75t_L g15188 ( 
.A(n_14784),
.B(n_2405),
.C(n_2406),
.Y(n_15188)
);

OAI21xp5_ASAP7_75t_L g15189 ( 
.A1(n_14797),
.A2(n_2407),
.B(n_2408),
.Y(n_15189)
);

OR2x2_ASAP7_75t_L g15190 ( 
.A(n_14861),
.B(n_2408),
.Y(n_15190)
);

INVx1_ASAP7_75t_L g15191 ( 
.A(n_14727),
.Y(n_15191)
);

CKINVDCx16_ASAP7_75t_R g15192 ( 
.A(n_15017),
.Y(n_15192)
);

AND2x4_ASAP7_75t_L g15193 ( 
.A(n_14762),
.B(n_2409),
.Y(n_15193)
);

INVx1_ASAP7_75t_L g15194 ( 
.A(n_14731),
.Y(n_15194)
);

AND2x2_ASAP7_75t_L g15195 ( 
.A(n_14671),
.B(n_2409),
.Y(n_15195)
);

INVx3_ASAP7_75t_L g15196 ( 
.A(n_14801),
.Y(n_15196)
);

CKINVDCx5p33_ASAP7_75t_R g15197 ( 
.A(n_15016),
.Y(n_15197)
);

BUFx3_ASAP7_75t_L g15198 ( 
.A(n_14993),
.Y(n_15198)
);

NOR2xp33_ASAP7_75t_R g15199 ( 
.A(n_14838),
.B(n_2410),
.Y(n_15199)
);

CKINVDCx5p33_ASAP7_75t_R g15200 ( 
.A(n_15010),
.Y(n_15200)
);

NOR3xp33_ASAP7_75t_SL g15201 ( 
.A(n_14728),
.B(n_2410),
.C(n_2411),
.Y(n_15201)
);

NAND2xp5_ASAP7_75t_L g15202 ( 
.A(n_14943),
.B(n_2411),
.Y(n_15202)
);

NAND2xp33_ASAP7_75t_R g15203 ( 
.A(n_14895),
.B(n_2412),
.Y(n_15203)
);

AND2x4_ASAP7_75t_SL g15204 ( 
.A(n_14927),
.B(n_2412),
.Y(n_15204)
);

HB1xp67_ASAP7_75t_L g15205 ( 
.A(n_14791),
.Y(n_15205)
);

CKINVDCx16_ASAP7_75t_R g15206 ( 
.A(n_14997),
.Y(n_15206)
);

AND2x2_ASAP7_75t_L g15207 ( 
.A(n_14986),
.B(n_2413),
.Y(n_15207)
);

INVx1_ASAP7_75t_L g15208 ( 
.A(n_14732),
.Y(n_15208)
);

OAI21xp5_ASAP7_75t_L g15209 ( 
.A1(n_14735),
.A2(n_2413),
.B(n_2414),
.Y(n_15209)
);

NAND3xp33_ASAP7_75t_L g15210 ( 
.A(n_14736),
.B(n_2414),
.C(n_2415),
.Y(n_15210)
);

OAI22xp5_ASAP7_75t_L g15211 ( 
.A1(n_14973),
.A2(n_14974),
.B1(n_14779),
.B2(n_15005),
.Y(n_15211)
);

AO21x2_ASAP7_75t_L g15212 ( 
.A1(n_14866),
.A2(n_2415),
.B(n_2416),
.Y(n_15212)
);

BUFx8_ASAP7_75t_SL g15213 ( 
.A(n_14888),
.Y(n_15213)
);

INVx4_ASAP7_75t_L g15214 ( 
.A(n_14904),
.Y(n_15214)
);

AND2x2_ASAP7_75t_L g15215 ( 
.A(n_14668),
.B(n_14922),
.Y(n_15215)
);

BUFx3_ASAP7_75t_L g15216 ( 
.A(n_14944),
.Y(n_15216)
);

AND2x2_ASAP7_75t_L g15217 ( 
.A(n_14901),
.B(n_2416),
.Y(n_15217)
);

BUFx3_ASAP7_75t_L g15218 ( 
.A(n_14875),
.Y(n_15218)
);

NOR2x1_ASAP7_75t_R g15219 ( 
.A(n_14769),
.B(n_2417),
.Y(n_15219)
);

NAND2xp5_ASAP7_75t_L g15220 ( 
.A(n_15003),
.B(n_2417),
.Y(n_15220)
);

OR2x2_ASAP7_75t_L g15221 ( 
.A(n_14831),
.B(n_2418),
.Y(n_15221)
);

INVx1_ASAP7_75t_L g15222 ( 
.A(n_14739),
.Y(n_15222)
);

NAND2xp33_ASAP7_75t_R g15223 ( 
.A(n_14698),
.B(n_2418),
.Y(n_15223)
);

HB1xp67_ASAP7_75t_L g15224 ( 
.A(n_14887),
.Y(n_15224)
);

INVx3_ASAP7_75t_L g15225 ( 
.A(n_14770),
.Y(n_15225)
);

OR2x6_ASAP7_75t_L g15226 ( 
.A(n_14987),
.B(n_2419),
.Y(n_15226)
);

NOR2xp33_ASAP7_75t_L g15227 ( 
.A(n_14976),
.B(n_2419),
.Y(n_15227)
);

AOI22xp33_ASAP7_75t_L g15228 ( 
.A1(n_14682),
.A2(n_14956),
.B1(n_14955),
.B2(n_14952),
.Y(n_15228)
);

AOI22xp33_ASAP7_75t_L g15229 ( 
.A1(n_15021),
.A2(n_2422),
.B1(n_2420),
.B2(n_2421),
.Y(n_15229)
);

NAND2xp33_ASAP7_75t_R g15230 ( 
.A(n_14799),
.B(n_2420),
.Y(n_15230)
);

NOR2xp33_ASAP7_75t_L g15231 ( 
.A(n_14992),
.B(n_2421),
.Y(n_15231)
);

AOI22xp5_ASAP7_75t_L g15232 ( 
.A1(n_14950),
.A2(n_2424),
.B1(n_2422),
.B2(n_2423),
.Y(n_15232)
);

INVx1_ASAP7_75t_L g15233 ( 
.A(n_14742),
.Y(n_15233)
);

NAND2xp33_ASAP7_75t_SL g15234 ( 
.A(n_15018),
.B(n_2426),
.Y(n_15234)
);

INVx1_ASAP7_75t_L g15235 ( 
.A(n_14743),
.Y(n_15235)
);

NAND2xp33_ASAP7_75t_R g15236 ( 
.A(n_14753),
.B(n_2426),
.Y(n_15236)
);

INVx2_ASAP7_75t_L g15237 ( 
.A(n_14965),
.Y(n_15237)
);

INVx1_ASAP7_75t_L g15238 ( 
.A(n_14745),
.Y(n_15238)
);

OR2x6_ASAP7_75t_L g15239 ( 
.A(n_14756),
.B(n_2427),
.Y(n_15239)
);

OR2x2_ASAP7_75t_L g15240 ( 
.A(n_14832),
.B(n_2427),
.Y(n_15240)
);

CKINVDCx16_ASAP7_75t_R g15241 ( 
.A(n_14844),
.Y(n_15241)
);

INVx2_ASAP7_75t_SL g15242 ( 
.A(n_14816),
.Y(n_15242)
);

CKINVDCx5p33_ASAP7_75t_R g15243 ( 
.A(n_14994),
.Y(n_15243)
);

CKINVDCx5p33_ASAP7_75t_R g15244 ( 
.A(n_14737),
.Y(n_15244)
);

NOR2xp33_ASAP7_75t_L g15245 ( 
.A(n_14934),
.B(n_2428),
.Y(n_15245)
);

BUFx12f_ASAP7_75t_L g15246 ( 
.A(n_14918),
.Y(n_15246)
);

INVx1_ASAP7_75t_L g15247 ( 
.A(n_14750),
.Y(n_15247)
);

NOR2xp33_ASAP7_75t_R g15248 ( 
.A(n_14969),
.B(n_2428),
.Y(n_15248)
);

OR2x4_ASAP7_75t_L g15249 ( 
.A(n_14693),
.B(n_2429),
.Y(n_15249)
);

INVx1_ASAP7_75t_L g15250 ( 
.A(n_14764),
.Y(n_15250)
);

NAND2xp5_ASAP7_75t_L g15251 ( 
.A(n_15008),
.B(n_2429),
.Y(n_15251)
);

AOI22xp33_ASAP7_75t_L g15252 ( 
.A1(n_15024),
.A2(n_2432),
.B1(n_2430),
.B2(n_2431),
.Y(n_15252)
);

BUFx10_ASAP7_75t_L g15253 ( 
.A(n_14872),
.Y(n_15253)
);

AO31x2_ASAP7_75t_L g15254 ( 
.A1(n_14852),
.A2(n_2433),
.A3(n_2430),
.B(n_2432),
.Y(n_15254)
);

INVx1_ASAP7_75t_L g15255 ( 
.A(n_14766),
.Y(n_15255)
);

BUFx3_ASAP7_75t_L g15256 ( 
.A(n_14972),
.Y(n_15256)
);

CKINVDCx5p33_ASAP7_75t_R g15257 ( 
.A(n_14824),
.Y(n_15257)
);

INVx2_ASAP7_75t_L g15258 ( 
.A(n_14951),
.Y(n_15258)
);

INVx2_ASAP7_75t_L g15259 ( 
.A(n_14714),
.Y(n_15259)
);

INVx1_ASAP7_75t_L g15260 ( 
.A(n_14774),
.Y(n_15260)
);

AO31x2_ASAP7_75t_L g15261 ( 
.A1(n_14850),
.A2(n_2435),
.A3(n_2433),
.B(n_2434),
.Y(n_15261)
);

INVx2_ASAP7_75t_L g15262 ( 
.A(n_14933),
.Y(n_15262)
);

AOI22xp33_ASAP7_75t_SL g15263 ( 
.A1(n_14968),
.A2(n_2436),
.B1(n_2434),
.B2(n_2435),
.Y(n_15263)
);

AND2x2_ASAP7_75t_L g15264 ( 
.A(n_14911),
.B(n_2436),
.Y(n_15264)
);

INVx3_ASAP7_75t_L g15265 ( 
.A(n_14765),
.Y(n_15265)
);

AOI21x1_ASAP7_75t_L g15266 ( 
.A1(n_14836),
.A2(n_2437),
.B(n_2438),
.Y(n_15266)
);

INVx1_ASAP7_75t_L g15267 ( 
.A(n_14815),
.Y(n_15267)
);

INVx1_ASAP7_75t_L g15268 ( 
.A(n_14835),
.Y(n_15268)
);

INVx1_ASAP7_75t_L g15269 ( 
.A(n_14837),
.Y(n_15269)
);

NAND2xp5_ASAP7_75t_L g15270 ( 
.A(n_14874),
.B(n_2439),
.Y(n_15270)
);

INVx2_ASAP7_75t_L g15271 ( 
.A(n_14924),
.Y(n_15271)
);

AND2x4_ASAP7_75t_L g15272 ( 
.A(n_14867),
.B(n_2440),
.Y(n_15272)
);

BUFx6f_ASAP7_75t_L g15273 ( 
.A(n_14907),
.Y(n_15273)
);

NAND2xp33_ASAP7_75t_R g15274 ( 
.A(n_14725),
.B(n_2440),
.Y(n_15274)
);

NOR2xp33_ASAP7_75t_R g15275 ( 
.A(n_14899),
.B(n_14999),
.Y(n_15275)
);

INVx1_ASAP7_75t_L g15276 ( 
.A(n_14841),
.Y(n_15276)
);

INVx2_ASAP7_75t_L g15277 ( 
.A(n_14923),
.Y(n_15277)
);

NOR3xp33_ASAP7_75t_SL g15278 ( 
.A(n_14880),
.B(n_2441),
.C(n_2442),
.Y(n_15278)
);

INVx2_ASAP7_75t_L g15279 ( 
.A(n_14908),
.Y(n_15279)
);

BUFx2_ASAP7_75t_L g15280 ( 
.A(n_14853),
.Y(n_15280)
);

HB1xp67_ASAP7_75t_L g15281 ( 
.A(n_14709),
.Y(n_15281)
);

INVx6_ASAP7_75t_L g15282 ( 
.A(n_14930),
.Y(n_15282)
);

NAND2xp5_ASAP7_75t_L g15283 ( 
.A(n_14863),
.B(n_2441),
.Y(n_15283)
);

INVx2_ASAP7_75t_L g15284 ( 
.A(n_14794),
.Y(n_15284)
);

INVxp67_ASAP7_75t_L g15285 ( 
.A(n_14755),
.Y(n_15285)
);

INVx1_ASAP7_75t_L g15286 ( 
.A(n_14842),
.Y(n_15286)
);

AND2x4_ASAP7_75t_L g15287 ( 
.A(n_14942),
.B(n_2442),
.Y(n_15287)
);

INVx1_ASAP7_75t_L g15288 ( 
.A(n_14849),
.Y(n_15288)
);

AOI21xp5_ASAP7_75t_L g15289 ( 
.A1(n_14981),
.A2(n_2443),
.B(n_2444),
.Y(n_15289)
);

AND2x2_ASAP7_75t_L g15290 ( 
.A(n_15057),
.B(n_14947),
.Y(n_15290)
);

AND2x2_ASAP7_75t_L g15291 ( 
.A(n_15045),
.B(n_14696),
.Y(n_15291)
);

OR2x2_ASAP7_75t_L g15292 ( 
.A(n_15096),
.B(n_14712),
.Y(n_15292)
);

INVx1_ASAP7_75t_L g15293 ( 
.A(n_15046),
.Y(n_15293)
);

OAI21xp5_ASAP7_75t_L g15294 ( 
.A1(n_15067),
.A2(n_15140),
.B(n_15065),
.Y(n_15294)
);

O2A1O1Ixp33_ASAP7_75t_L g15295 ( 
.A1(n_15065),
.A2(n_14859),
.B(n_14780),
.C(n_14819),
.Y(n_15295)
);

AOI22xp33_ASAP7_75t_L g15296 ( 
.A1(n_15128),
.A2(n_14971),
.B1(n_14865),
.B2(n_14970),
.Y(n_15296)
);

BUFx3_ASAP7_75t_L g15297 ( 
.A(n_15031),
.Y(n_15297)
);

NAND2xp33_ASAP7_75t_R g15298 ( 
.A(n_15199),
.B(n_15201),
.Y(n_15298)
);

AND2x4_ASAP7_75t_L g15299 ( 
.A(n_15082),
.B(n_14984),
.Y(n_15299)
);

AND2x2_ASAP7_75t_L g15300 ( 
.A(n_15058),
.B(n_14945),
.Y(n_15300)
);

NOR2xp33_ASAP7_75t_L g15301 ( 
.A(n_15106),
.B(n_14871),
.Y(n_15301)
);

AND2x2_ASAP7_75t_L g15302 ( 
.A(n_15030),
.B(n_14946),
.Y(n_15302)
);

CKINVDCx5p33_ASAP7_75t_R g15303 ( 
.A(n_15043),
.Y(n_15303)
);

INVx1_ASAP7_75t_L g15304 ( 
.A(n_15051),
.Y(n_15304)
);

AO21x2_ASAP7_75t_L g15305 ( 
.A1(n_15281),
.A2(n_14857),
.B(n_14848),
.Y(n_15305)
);

A2O1A1Ixp33_ASAP7_75t_L g15306 ( 
.A1(n_15133),
.A2(n_15000),
.B(n_14834),
.C(n_14868),
.Y(n_15306)
);

AND2x2_ASAP7_75t_L g15307 ( 
.A(n_15098),
.B(n_14667),
.Y(n_15307)
);

OR2x2_ASAP7_75t_L g15308 ( 
.A(n_15072),
.B(n_14882),
.Y(n_15308)
);

INVx1_ASAP7_75t_L g15309 ( 
.A(n_15040),
.Y(n_15309)
);

AOI221xp5_ASAP7_75t_L g15310 ( 
.A1(n_15228),
.A2(n_14811),
.B1(n_14823),
.B2(n_14886),
.C(n_14778),
.Y(n_15310)
);

BUFx2_ASAP7_75t_L g15311 ( 
.A(n_15213),
.Y(n_15311)
);

AND2x4_ASAP7_75t_L g15312 ( 
.A(n_15198),
.B(n_14905),
.Y(n_15312)
);

AO32x2_ASAP7_75t_L g15313 ( 
.A1(n_15211),
.A2(n_14787),
.A3(n_14879),
.B1(n_14917),
.B2(n_14910),
.Y(n_15313)
);

O2A1O1Ixp33_ASAP7_75t_SL g15314 ( 
.A1(n_15285),
.A2(n_14763),
.B(n_14675),
.C(n_14768),
.Y(n_15314)
);

NOR3xp33_ASAP7_75t_L g15315 ( 
.A(n_15192),
.B(n_14900),
.C(n_14892),
.Y(n_15315)
);

AND2x2_ASAP7_75t_L g15316 ( 
.A(n_15241),
.B(n_14935),
.Y(n_15316)
);

INVx2_ASAP7_75t_L g15317 ( 
.A(n_15028),
.Y(n_15317)
);

BUFx4f_ASAP7_75t_SL g15318 ( 
.A(n_15076),
.Y(n_15318)
);

NOR2xp33_ASAP7_75t_L g15319 ( 
.A(n_15106),
.B(n_14884),
.Y(n_15319)
);

AND2x2_ASAP7_75t_L g15320 ( 
.A(n_15144),
.B(n_14936),
.Y(n_15320)
);

INVx2_ASAP7_75t_L g15321 ( 
.A(n_15028),
.Y(n_15321)
);

AOI221xp5_ASAP7_75t_L g15322 ( 
.A1(n_15166),
.A2(n_14894),
.B1(n_14897),
.B2(n_14893),
.C(n_14798),
.Y(n_15322)
);

AND2x2_ASAP7_75t_L g15323 ( 
.A(n_15080),
.B(n_14964),
.Y(n_15323)
);

AND2x2_ASAP7_75t_L g15324 ( 
.A(n_15056),
.B(n_14851),
.Y(n_15324)
);

AO21x2_ASAP7_75t_L g15325 ( 
.A1(n_15167),
.A2(n_14786),
.B(n_14759),
.Y(n_15325)
);

A2O1A1Ixp33_ASAP7_75t_L g15326 ( 
.A1(n_15234),
.A2(n_14877),
.B(n_14854),
.C(n_14710),
.Y(n_15326)
);

OR2x6_ASAP7_75t_L g15327 ( 
.A(n_15056),
.B(n_14928),
.Y(n_15327)
);

AND2x2_ASAP7_75t_L g15328 ( 
.A(n_15084),
.B(n_14959),
.Y(n_15328)
);

AND2x4_ASAP7_75t_L g15329 ( 
.A(n_15218),
.B(n_15050),
.Y(n_15329)
);

INVx3_ASAP7_75t_L g15330 ( 
.A(n_15185),
.Y(n_15330)
);

AND2x4_ASAP7_75t_L g15331 ( 
.A(n_15054),
.B(n_14771),
.Y(n_15331)
);

OR2x2_ASAP7_75t_L g15332 ( 
.A(n_15027),
.B(n_14829),
.Y(n_15332)
);

AO32x2_ASAP7_75t_L g15333 ( 
.A1(n_15242),
.A2(n_14787),
.A3(n_14709),
.B1(n_14856),
.B2(n_14858),
.Y(n_15333)
);

OAI21xp5_ASAP7_75t_L g15334 ( 
.A1(n_15071),
.A2(n_14676),
.B(n_14795),
.Y(n_15334)
);

A2O1A1Ixp33_ASAP7_75t_L g15335 ( 
.A1(n_15063),
.A2(n_14847),
.B(n_14827),
.C(n_14940),
.Y(n_15335)
);

INVx1_ASAP7_75t_L g15336 ( 
.A(n_15041),
.Y(n_15336)
);

AO21x2_ASAP7_75t_L g15337 ( 
.A1(n_15112),
.A2(n_14805),
.B(n_14790),
.Y(n_15337)
);

AND2x4_ASAP7_75t_L g15338 ( 
.A(n_15026),
.B(n_14782),
.Y(n_15338)
);

NAND2xp5_ASAP7_75t_L g15339 ( 
.A(n_15085),
.B(n_14960),
.Y(n_15339)
);

NAND2xp5_ASAP7_75t_L g15340 ( 
.A(n_15244),
.B(n_14748),
.Y(n_15340)
);

AND2x2_ASAP7_75t_L g15341 ( 
.A(n_15097),
.B(n_14873),
.Y(n_15341)
);

AND2x2_ASAP7_75t_L g15342 ( 
.A(n_15151),
.B(n_15032),
.Y(n_15342)
);

NOR2xp33_ASAP7_75t_L g15343 ( 
.A(n_15060),
.B(n_14789),
.Y(n_15343)
);

AOI21xp5_ASAP7_75t_L g15344 ( 
.A1(n_15042),
.A2(n_14722),
.B(n_14855),
.Y(n_15344)
);

NAND2x1_ASAP7_75t_L g15345 ( 
.A(n_15282),
.B(n_14775),
.Y(n_15345)
);

OAI21xp5_ASAP7_75t_L g15346 ( 
.A1(n_15126),
.A2(n_15209),
.B(n_15048),
.Y(n_15346)
);

OA21x2_ASAP7_75t_L g15347 ( 
.A1(n_15180),
.A2(n_14843),
.B(n_14822),
.Y(n_15347)
);

AND2x2_ASAP7_75t_L g15348 ( 
.A(n_15044),
.B(n_14802),
.Y(n_15348)
);

CKINVDCx6p67_ASAP7_75t_R g15349 ( 
.A(n_15186),
.Y(n_15349)
);

BUFx2_ASAP7_75t_L g15350 ( 
.A(n_15246),
.Y(n_15350)
);

INVx1_ASAP7_75t_L g15351 ( 
.A(n_15137),
.Y(n_15351)
);

INVx1_ASAP7_75t_SL g15352 ( 
.A(n_15053),
.Y(n_15352)
);

AND2x2_ASAP7_75t_L g15353 ( 
.A(n_15152),
.B(n_14825),
.Y(n_15353)
);

INVxp67_ASAP7_75t_L g15354 ( 
.A(n_15230),
.Y(n_15354)
);

NAND2xp5_ASAP7_75t_L g15355 ( 
.A(n_15038),
.B(n_14783),
.Y(n_15355)
);

A2O1A1Ixp33_ASAP7_75t_L g15356 ( 
.A1(n_15232),
.A2(n_14885),
.B(n_14840),
.C(n_14741),
.Y(n_15356)
);

AOI22xp33_ASAP7_75t_L g15357 ( 
.A1(n_15048),
.A2(n_14860),
.B1(n_14862),
.B2(n_14826),
.Y(n_15357)
);

A2O1A1Ixp33_ASAP7_75t_L g15358 ( 
.A1(n_15113),
.A2(n_14881),
.B(n_14793),
.C(n_14796),
.Y(n_15358)
);

OAI21xp5_ASAP7_75t_L g15359 ( 
.A1(n_15210),
.A2(n_15188),
.B(n_15025),
.Y(n_15359)
);

AOI22xp5_ASAP7_75t_L g15360 ( 
.A1(n_15066),
.A2(n_14800),
.B1(n_14803),
.B2(n_14792),
.Y(n_15360)
);

INVx3_ASAP7_75t_L g15361 ( 
.A(n_15093),
.Y(n_15361)
);

INVx2_ASAP7_75t_L g15362 ( 
.A(n_15081),
.Y(n_15362)
);

HB1xp67_ASAP7_75t_L g15363 ( 
.A(n_15226),
.Y(n_15363)
);

OR2x2_ASAP7_75t_L g15364 ( 
.A(n_15033),
.B(n_14804),
.Y(n_15364)
);

OA21x2_ASAP7_75t_L g15365 ( 
.A1(n_15224),
.A2(n_14809),
.B(n_14807),
.Y(n_15365)
);

OR2x2_ASAP7_75t_L g15366 ( 
.A(n_15104),
.B(n_15047),
.Y(n_15366)
);

AOI21xp5_ASAP7_75t_L g15367 ( 
.A1(n_15156),
.A2(n_14808),
.B(n_14806),
.Y(n_15367)
);

NAND2xp5_ASAP7_75t_L g15368 ( 
.A(n_15200),
.B(n_2443),
.Y(n_15368)
);

AND2x2_ASAP7_75t_L g15369 ( 
.A(n_15095),
.B(n_2444),
.Y(n_15369)
);

OAI211xp5_ASAP7_75t_L g15370 ( 
.A1(n_15121),
.A2(n_2447),
.B(n_2445),
.C(n_2446),
.Y(n_15370)
);

AO32x2_ASAP7_75t_L g15371 ( 
.A1(n_15214),
.A2(n_2447),
.A3(n_2445),
.B1(n_2446),
.B2(n_2448),
.Y(n_15371)
);

AND2x2_ASAP7_75t_L g15372 ( 
.A(n_15111),
.B(n_2448),
.Y(n_15372)
);

NAND2xp5_ASAP7_75t_L g15373 ( 
.A(n_15068),
.B(n_15206),
.Y(n_15373)
);

CKINVDCx5p33_ASAP7_75t_R g15374 ( 
.A(n_15049),
.Y(n_15374)
);

AO32x2_ASAP7_75t_L g15375 ( 
.A1(n_15120),
.A2(n_2451),
.A3(n_2449),
.B1(n_2450),
.B2(n_2452),
.Y(n_15375)
);

OAI21xp5_ASAP7_75t_L g15376 ( 
.A1(n_15127),
.A2(n_2450),
.B(n_2451),
.Y(n_15376)
);

INVx3_ASAP7_75t_L g15377 ( 
.A(n_15093),
.Y(n_15377)
);

INVx1_ASAP7_75t_L g15378 ( 
.A(n_15108),
.Y(n_15378)
);

AND2x2_ASAP7_75t_L g15379 ( 
.A(n_15081),
.B(n_2452),
.Y(n_15379)
);

OR2x2_ASAP7_75t_L g15380 ( 
.A(n_15159),
.B(n_2453),
.Y(n_15380)
);

BUFx3_ASAP7_75t_L g15381 ( 
.A(n_15091),
.Y(n_15381)
);

OR2x2_ASAP7_75t_L g15382 ( 
.A(n_15029),
.B(n_2454),
.Y(n_15382)
);

AOI22xp33_ASAP7_75t_L g15383 ( 
.A1(n_15036),
.A2(n_2456),
.B1(n_2454),
.B2(n_2455),
.Y(n_15383)
);

HB1xp67_ASAP7_75t_L g15384 ( 
.A(n_15226),
.Y(n_15384)
);

INVx5_ASAP7_75t_SL g15385 ( 
.A(n_15132),
.Y(n_15385)
);

O2A1O1Ixp33_ASAP7_75t_L g15386 ( 
.A1(n_15035),
.A2(n_2458),
.B(n_2456),
.C(n_2457),
.Y(n_15386)
);

AOI22xp33_ASAP7_75t_L g15387 ( 
.A1(n_15145),
.A2(n_2460),
.B1(n_2457),
.B2(n_2459),
.Y(n_15387)
);

AND2x2_ASAP7_75t_L g15388 ( 
.A(n_15174),
.B(n_15125),
.Y(n_15388)
);

OR2x2_ASAP7_75t_L g15389 ( 
.A(n_15034),
.B(n_15039),
.Y(n_15389)
);

AOI21xp5_ASAP7_75t_L g15390 ( 
.A1(n_15289),
.A2(n_2459),
.B(n_2460),
.Y(n_15390)
);

CKINVDCx11_ASAP7_75t_R g15391 ( 
.A(n_15091),
.Y(n_15391)
);

OAI22xp5_ASAP7_75t_L g15392 ( 
.A1(n_15145),
.A2(n_2463),
.B1(n_2461),
.B2(n_2462),
.Y(n_15392)
);

NOR2xp33_ASAP7_75t_L g15393 ( 
.A(n_15183),
.B(n_15164),
.Y(n_15393)
);

AND2x2_ASAP7_75t_L g15394 ( 
.A(n_15146),
.B(n_2461),
.Y(n_15394)
);

OR2x2_ASAP7_75t_L g15395 ( 
.A(n_15069),
.B(n_15059),
.Y(n_15395)
);

AND2x4_ASAP7_75t_L g15396 ( 
.A(n_15122),
.B(n_2462),
.Y(n_15396)
);

AOI21xp5_ASAP7_75t_L g15397 ( 
.A1(n_15035),
.A2(n_2464),
.B(n_2465),
.Y(n_15397)
);

NOR2x1_ASAP7_75t_SL g15398 ( 
.A(n_15212),
.B(n_2465),
.Y(n_15398)
);

BUFx12f_ASAP7_75t_L g15399 ( 
.A(n_15243),
.Y(n_15399)
);

OR2x2_ASAP7_75t_L g15400 ( 
.A(n_15190),
.B(n_2466),
.Y(n_15400)
);

OA21x2_ASAP7_75t_L g15401 ( 
.A1(n_15173),
.A2(n_2466),
.B(n_2467),
.Y(n_15401)
);

INVx1_ASAP7_75t_L g15402 ( 
.A(n_15176),
.Y(n_15402)
);

INVx1_ASAP7_75t_L g15403 ( 
.A(n_15205),
.Y(n_15403)
);

AND2x2_ASAP7_75t_L g15404 ( 
.A(n_15109),
.B(n_2467),
.Y(n_15404)
);

CKINVDCx5p33_ASAP7_75t_R g15405 ( 
.A(n_15236),
.Y(n_15405)
);

BUFx3_ASAP7_75t_L g15406 ( 
.A(n_15124),
.Y(n_15406)
);

CKINVDCx14_ASAP7_75t_R g15407 ( 
.A(n_15148),
.Y(n_15407)
);

AND2x4_ASAP7_75t_L g15408 ( 
.A(n_15115),
.B(n_2468),
.Y(n_15408)
);

INVx1_ASAP7_75t_L g15409 ( 
.A(n_15052),
.Y(n_15409)
);

OR2x2_ASAP7_75t_L g15410 ( 
.A(n_15256),
.B(n_2468),
.Y(n_15410)
);

AOI21xp5_ASAP7_75t_L g15411 ( 
.A1(n_15202),
.A2(n_2469),
.B(n_2470),
.Y(n_15411)
);

INVx1_ASAP7_75t_L g15412 ( 
.A(n_15253),
.Y(n_15412)
);

AO32x2_ASAP7_75t_L g15413 ( 
.A1(n_15274),
.A2(n_15223),
.A3(n_15055),
.B1(n_15249),
.B2(n_15182),
.Y(n_15413)
);

INVx1_ASAP7_75t_L g15414 ( 
.A(n_15221),
.Y(n_15414)
);

HB1xp67_ASAP7_75t_L g15415 ( 
.A(n_15197),
.Y(n_15415)
);

O2A1O1Ixp33_ASAP7_75t_SL g15416 ( 
.A1(n_15189),
.A2(n_2472),
.B(n_2469),
.C(n_2471),
.Y(n_15416)
);

INVx2_ASAP7_75t_L g15417 ( 
.A(n_15273),
.Y(n_15417)
);

A2O1A1Ixp33_ASAP7_75t_L g15418 ( 
.A1(n_15102),
.A2(n_2474),
.B(n_2471),
.C(n_2473),
.Y(n_15418)
);

INVx2_ASAP7_75t_L g15419 ( 
.A(n_15273),
.Y(n_15419)
);

AOI21xp33_ASAP7_75t_SL g15420 ( 
.A1(n_15116),
.A2(n_2474),
.B(n_2475),
.Y(n_15420)
);

AO21x2_ASAP7_75t_L g15421 ( 
.A1(n_15181),
.A2(n_2475),
.B(n_2476),
.Y(n_15421)
);

AND2x4_ASAP7_75t_L g15422 ( 
.A(n_15162),
.B(n_2476),
.Y(n_15422)
);

NOR2x1_ASAP7_75t_SL g15423 ( 
.A(n_15110),
.B(n_2477),
.Y(n_15423)
);

AND2x4_ASAP7_75t_L g15424 ( 
.A(n_15157),
.B(n_2478),
.Y(n_15424)
);

OAI22xp5_ASAP7_75t_L g15425 ( 
.A1(n_15257),
.A2(n_2481),
.B1(n_2479),
.B2(n_2480),
.Y(n_15425)
);

AO21x2_ASAP7_75t_L g15426 ( 
.A1(n_15118),
.A2(n_2479),
.B(n_2480),
.Y(n_15426)
);

OR2x6_ASAP7_75t_L g15427 ( 
.A(n_15114),
.B(n_15138),
.Y(n_15427)
);

NAND2x1_ASAP7_75t_L g15428 ( 
.A(n_15280),
.B(n_2481),
.Y(n_15428)
);

AND2x2_ASAP7_75t_L g15429 ( 
.A(n_15215),
.B(n_2482),
.Y(n_15429)
);

NOR2x1_ASAP7_75t_SL g15430 ( 
.A(n_15110),
.B(n_2482),
.Y(n_15430)
);

AND2x4_ASAP7_75t_SL g15431 ( 
.A(n_15239),
.B(n_15092),
.Y(n_15431)
);

INVx1_ASAP7_75t_L g15432 ( 
.A(n_15240),
.Y(n_15432)
);

CKINVDCx10_ASAP7_75t_R g15433 ( 
.A(n_15239),
.Y(n_15433)
);

AND2x2_ASAP7_75t_L g15434 ( 
.A(n_15165),
.B(n_2483),
.Y(n_15434)
);

BUFx5_ASAP7_75t_L g15435 ( 
.A(n_15089),
.Y(n_15435)
);

AOI21xp5_ASAP7_75t_L g15436 ( 
.A1(n_15227),
.A2(n_2484),
.B(n_2485),
.Y(n_15436)
);

HB1xp67_ASAP7_75t_L g15437 ( 
.A(n_15275),
.Y(n_15437)
);

AND2x2_ASAP7_75t_L g15438 ( 
.A(n_15177),
.B(n_2484),
.Y(n_15438)
);

INVx1_ASAP7_75t_L g15439 ( 
.A(n_15153),
.Y(n_15439)
);

OAI211xp5_ASAP7_75t_L g15440 ( 
.A1(n_15263),
.A2(n_2487),
.B(n_2485),
.C(n_2486),
.Y(n_15440)
);

AND2x4_ASAP7_75t_SL g15441 ( 
.A(n_15272),
.B(n_2486),
.Y(n_15441)
);

AOI22xp5_ASAP7_75t_L g15442 ( 
.A1(n_15203),
.A2(n_15171),
.B1(n_15123),
.B2(n_15037),
.Y(n_15442)
);

AND2x2_ASAP7_75t_L g15443 ( 
.A(n_15196),
.B(n_2487),
.Y(n_15443)
);

AND2x2_ASAP7_75t_L g15444 ( 
.A(n_15225),
.B(n_2488),
.Y(n_15444)
);

INVx1_ASAP7_75t_L g15445 ( 
.A(n_15129),
.Y(n_15445)
);

OAI21xp5_ASAP7_75t_SL g15446 ( 
.A1(n_15119),
.A2(n_2488),
.B(n_2489),
.Y(n_15446)
);

NOR2x1_ASAP7_75t_SL g15447 ( 
.A(n_15195),
.B(n_2489),
.Y(n_15447)
);

INVx2_ASAP7_75t_L g15448 ( 
.A(n_15175),
.Y(n_15448)
);

A2O1A1Ixp33_ASAP7_75t_L g15449 ( 
.A1(n_15278),
.A2(n_2492),
.B(n_2490),
.C(n_2491),
.Y(n_15449)
);

INVxp67_ASAP7_75t_L g15450 ( 
.A(n_15219),
.Y(n_15450)
);

AND2x2_ASAP7_75t_L g15451 ( 
.A(n_15265),
.B(n_2490),
.Y(n_15451)
);

AND2x2_ASAP7_75t_L g15452 ( 
.A(n_15216),
.B(n_2491),
.Y(n_15452)
);

INVx1_ASAP7_75t_L g15453 ( 
.A(n_15207),
.Y(n_15453)
);

INVx1_ASAP7_75t_L g15454 ( 
.A(n_15061),
.Y(n_15454)
);

NOR2x1_ASAP7_75t_SL g15455 ( 
.A(n_15266),
.B(n_2492),
.Y(n_15455)
);

AND2x2_ASAP7_75t_L g15456 ( 
.A(n_15258),
.B(n_2493),
.Y(n_15456)
);

AND2x2_ASAP7_75t_L g15457 ( 
.A(n_15070),
.B(n_2494),
.Y(n_15457)
);

BUFx2_ASAP7_75t_L g15458 ( 
.A(n_15248),
.Y(n_15458)
);

AND2x4_ASAP7_75t_L g15459 ( 
.A(n_15099),
.B(n_2494),
.Y(n_15459)
);

OAI21xp5_ASAP7_75t_L g15460 ( 
.A1(n_15088),
.A2(n_2495),
.B(n_2496),
.Y(n_15460)
);

A2O1A1Ixp33_ASAP7_75t_L g15461 ( 
.A1(n_15055),
.A2(n_2498),
.B(n_2496),
.C(n_2497),
.Y(n_15461)
);

BUFx3_ASAP7_75t_L g15462 ( 
.A(n_15204),
.Y(n_15462)
);

AND2x2_ASAP7_75t_L g15463 ( 
.A(n_15259),
.B(n_2497),
.Y(n_15463)
);

BUFx2_ASAP7_75t_L g15464 ( 
.A(n_15100),
.Y(n_15464)
);

INVx2_ASAP7_75t_L g15465 ( 
.A(n_15079),
.Y(n_15465)
);

AND2x4_ASAP7_75t_L g15466 ( 
.A(n_15179),
.B(n_2498),
.Y(n_15466)
);

AND2x2_ASAP7_75t_L g15467 ( 
.A(n_15136),
.B(n_2499),
.Y(n_15467)
);

AND2x2_ASAP7_75t_L g15468 ( 
.A(n_15284),
.B(n_2500),
.Y(n_15468)
);

OAI22xp5_ASAP7_75t_L g15469 ( 
.A1(n_15229),
.A2(n_2503),
.B1(n_2501),
.B2(n_2502),
.Y(n_15469)
);

NAND2xp5_ASAP7_75t_L g15470 ( 
.A(n_15117),
.B(n_2501),
.Y(n_15470)
);

NAND2xp33_ASAP7_75t_R g15471 ( 
.A(n_15086),
.B(n_2502),
.Y(n_15471)
);

A2O1A1Ixp33_ASAP7_75t_L g15472 ( 
.A1(n_15187),
.A2(n_15252),
.B(n_15147),
.C(n_15150),
.Y(n_15472)
);

AND2x4_ASAP7_75t_L g15473 ( 
.A(n_15271),
.B(n_2503),
.Y(n_15473)
);

INVx1_ASAP7_75t_L g15474 ( 
.A(n_15062),
.Y(n_15474)
);

NOR2x1_ASAP7_75t_SL g15475 ( 
.A(n_15142),
.B(n_2504),
.Y(n_15475)
);

INVx2_ASAP7_75t_L g15476 ( 
.A(n_15087),
.Y(n_15476)
);

NAND2xp5_ASAP7_75t_L g15477 ( 
.A(n_15117),
.B(n_2505),
.Y(n_15477)
);

NOR2xp33_ASAP7_75t_L g15478 ( 
.A(n_15220),
.B(n_2505),
.Y(n_15478)
);

INVx1_ASAP7_75t_L g15479 ( 
.A(n_15064),
.Y(n_15479)
);

INVx1_ASAP7_75t_L g15480 ( 
.A(n_15073),
.Y(n_15480)
);

OR2x2_ASAP7_75t_L g15481 ( 
.A(n_15279),
.B(n_2506),
.Y(n_15481)
);

AND2x4_ASAP7_75t_L g15482 ( 
.A(n_15262),
.B(n_2506),
.Y(n_15482)
);

INVx5_ASAP7_75t_L g15483 ( 
.A(n_15090),
.Y(n_15483)
);

OAI21xp5_ASAP7_75t_L g15484 ( 
.A1(n_15149),
.A2(n_2507),
.B(n_2508),
.Y(n_15484)
);

INVx2_ASAP7_75t_L g15485 ( 
.A(n_15143),
.Y(n_15485)
);

NAND2xp5_ASAP7_75t_L g15486 ( 
.A(n_15277),
.B(n_15237),
.Y(n_15486)
);

AND2x2_ASAP7_75t_L g15487 ( 
.A(n_15103),
.B(n_2507),
.Y(n_15487)
);

AND2x2_ASAP7_75t_L g15488 ( 
.A(n_15083),
.B(n_2508),
.Y(n_15488)
);

A2O1A1Ixp33_ASAP7_75t_L g15489 ( 
.A1(n_15160),
.A2(n_2511),
.B(n_2509),
.C(n_2510),
.Y(n_15489)
);

O2A1O1Ixp33_ASAP7_75t_L g15490 ( 
.A1(n_15161),
.A2(n_2512),
.B(n_2509),
.C(n_2510),
.Y(n_15490)
);

INVxp67_ASAP7_75t_L g15491 ( 
.A(n_15231),
.Y(n_15491)
);

BUFx12f_ASAP7_75t_L g15492 ( 
.A(n_15169),
.Y(n_15492)
);

AND2x2_ASAP7_75t_L g15493 ( 
.A(n_15184),
.B(n_2512),
.Y(n_15493)
);

AO32x2_ASAP7_75t_L g15494 ( 
.A1(n_15078),
.A2(n_2515),
.A3(n_2513),
.B1(n_2514),
.B2(n_2516),
.Y(n_15494)
);

AOI21xp5_ASAP7_75t_L g15495 ( 
.A1(n_15295),
.A2(n_15163),
.B(n_15251),
.Y(n_15495)
);

AND2x2_ASAP7_75t_L g15496 ( 
.A(n_15349),
.B(n_15267),
.Y(n_15496)
);

AND2x2_ASAP7_75t_L g15497 ( 
.A(n_15311),
.B(n_15268),
.Y(n_15497)
);

AND2x2_ASAP7_75t_L g15498 ( 
.A(n_15297),
.B(n_15269),
.Y(n_15498)
);

INVx2_ASAP7_75t_L g15499 ( 
.A(n_15483),
.Y(n_15499)
);

INVx2_ASAP7_75t_L g15500 ( 
.A(n_15483),
.Y(n_15500)
);

INVx1_ASAP7_75t_L g15501 ( 
.A(n_15309),
.Y(n_15501)
);

INVx1_ASAP7_75t_L g15502 ( 
.A(n_15336),
.Y(n_15502)
);

INVx1_ASAP7_75t_L g15503 ( 
.A(n_15351),
.Y(n_15503)
);

AND2x4_ASAP7_75t_L g15504 ( 
.A(n_15462),
.B(n_15193),
.Y(n_15504)
);

INVx2_ASAP7_75t_L g15505 ( 
.A(n_15391),
.Y(n_15505)
);

HB1xp67_ASAP7_75t_L g15506 ( 
.A(n_15407),
.Y(n_15506)
);

INVx1_ASAP7_75t_SL g15507 ( 
.A(n_15433),
.Y(n_15507)
);

AOI22xp33_ASAP7_75t_L g15508 ( 
.A1(n_15315),
.A2(n_15276),
.B1(n_15288),
.B2(n_15286),
.Y(n_15508)
);

INVx1_ASAP7_75t_L g15509 ( 
.A(n_15403),
.Y(n_15509)
);

BUFx2_ASAP7_75t_L g15510 ( 
.A(n_15399),
.Y(n_15510)
);

INVx1_ASAP7_75t_L g15511 ( 
.A(n_15304),
.Y(n_15511)
);

AND2x2_ASAP7_75t_L g15512 ( 
.A(n_15350),
.B(n_15101),
.Y(n_15512)
);

OR2x2_ASAP7_75t_L g15513 ( 
.A(n_15354),
.B(n_15105),
.Y(n_15513)
);

AOI33xp33_ASAP7_75t_L g15514 ( 
.A1(n_15357),
.A2(n_15296),
.A3(n_15442),
.B1(n_15360),
.B2(n_15314),
.B3(n_15412),
.Y(n_15514)
);

OA21x2_ASAP7_75t_L g15515 ( 
.A1(n_15464),
.A2(n_15077),
.B(n_15075),
.Y(n_15515)
);

INVx2_ASAP7_75t_L g15516 ( 
.A(n_15435),
.Y(n_15516)
);

AND2x2_ASAP7_75t_L g15517 ( 
.A(n_15290),
.B(n_15458),
.Y(n_15517)
);

INVx1_ASAP7_75t_L g15518 ( 
.A(n_15380),
.Y(n_15518)
);

AND2x2_ASAP7_75t_L g15519 ( 
.A(n_15352),
.B(n_15074),
.Y(n_15519)
);

INVx2_ASAP7_75t_L g15520 ( 
.A(n_15435),
.Y(n_15520)
);

INVx2_ASAP7_75t_SL g15521 ( 
.A(n_15345),
.Y(n_15521)
);

OR2x2_ASAP7_75t_L g15522 ( 
.A(n_15373),
.B(n_15107),
.Y(n_15522)
);

INVx1_ASAP7_75t_L g15523 ( 
.A(n_15293),
.Y(n_15523)
);

OR2x2_ASAP7_75t_L g15524 ( 
.A(n_15363),
.B(n_15130),
.Y(n_15524)
);

AOI221xp5_ASAP7_75t_L g15525 ( 
.A1(n_15461),
.A2(n_15135),
.B1(n_15141),
.B2(n_15139),
.C(n_15131),
.Y(n_15525)
);

OR2x2_ASAP7_75t_L g15526 ( 
.A(n_15384),
.B(n_15154),
.Y(n_15526)
);

OR2x2_ASAP7_75t_L g15527 ( 
.A(n_15437),
.B(n_15158),
.Y(n_15527)
);

AND2x4_ASAP7_75t_L g15528 ( 
.A(n_15406),
.B(n_15178),
.Y(n_15528)
);

OR2x2_ASAP7_75t_L g15529 ( 
.A(n_15308),
.B(n_15292),
.Y(n_15529)
);

INVx1_ASAP7_75t_L g15530 ( 
.A(n_15378),
.Y(n_15530)
);

AND2x2_ASAP7_75t_L g15531 ( 
.A(n_15316),
.B(n_15217),
.Y(n_15531)
);

INVx3_ASAP7_75t_L g15532 ( 
.A(n_15492),
.Y(n_15532)
);

INVx1_ASAP7_75t_L g15533 ( 
.A(n_15389),
.Y(n_15533)
);

INVx1_ASAP7_75t_L g15534 ( 
.A(n_15402),
.Y(n_15534)
);

INVx2_ASAP7_75t_L g15535 ( 
.A(n_15435),
.Y(n_15535)
);

INVx1_ASAP7_75t_L g15536 ( 
.A(n_15481),
.Y(n_15536)
);

INVx2_ASAP7_75t_L g15537 ( 
.A(n_15330),
.Y(n_15537)
);

NAND2xp5_ASAP7_75t_L g15538 ( 
.A(n_15405),
.B(n_15264),
.Y(n_15538)
);

OAI21x1_ASAP7_75t_L g15539 ( 
.A1(n_15344),
.A2(n_15367),
.B(n_15365),
.Y(n_15539)
);

AND2x2_ASAP7_75t_L g15540 ( 
.A(n_15291),
.B(n_15155),
.Y(n_15540)
);

INVx2_ASAP7_75t_L g15541 ( 
.A(n_15318),
.Y(n_15541)
);

AOI21xp33_ASAP7_75t_L g15542 ( 
.A1(n_15334),
.A2(n_15170),
.B(n_15168),
.Y(n_15542)
);

INVx2_ASAP7_75t_L g15543 ( 
.A(n_15381),
.Y(n_15543)
);

INVxp67_ASAP7_75t_SL g15544 ( 
.A(n_15423),
.Y(n_15544)
);

INVx1_ASAP7_75t_L g15545 ( 
.A(n_15400),
.Y(n_15545)
);

OR2x2_ASAP7_75t_L g15546 ( 
.A(n_15366),
.B(n_15172),
.Y(n_15546)
);

INVx1_ASAP7_75t_L g15547 ( 
.A(n_15382),
.Y(n_15547)
);

AND2x2_ASAP7_75t_L g15548 ( 
.A(n_15385),
.B(n_15287),
.Y(n_15548)
);

AND2x4_ASAP7_75t_SL g15549 ( 
.A(n_15329),
.B(n_15245),
.Y(n_15549)
);

OAI22xp5_ASAP7_75t_L g15550 ( 
.A1(n_15335),
.A2(n_15270),
.B1(n_15283),
.B2(n_15191),
.Y(n_15550)
);

INVx2_ASAP7_75t_L g15551 ( 
.A(n_15361),
.Y(n_15551)
);

NAND2xp5_ASAP7_75t_L g15552 ( 
.A(n_15420),
.B(n_15094),
.Y(n_15552)
);

OR2x2_ASAP7_75t_L g15553 ( 
.A(n_15465),
.B(n_15194),
.Y(n_15553)
);

NOR2x1_ASAP7_75t_L g15554 ( 
.A(n_15305),
.B(n_15208),
.Y(n_15554)
);

AND2x2_ASAP7_75t_L g15555 ( 
.A(n_15427),
.B(n_15222),
.Y(n_15555)
);

OR2x2_ASAP7_75t_L g15556 ( 
.A(n_15332),
.B(n_15233),
.Y(n_15556)
);

HB1xp67_ASAP7_75t_L g15557 ( 
.A(n_15428),
.Y(n_15557)
);

NOR2x1_ASAP7_75t_L g15558 ( 
.A(n_15427),
.B(n_15235),
.Y(n_15558)
);

NAND2x1p5_ASAP7_75t_L g15559 ( 
.A(n_15459),
.B(n_15238),
.Y(n_15559)
);

INVx1_ASAP7_75t_L g15560 ( 
.A(n_15463),
.Y(n_15560)
);

INVx1_ASAP7_75t_L g15561 ( 
.A(n_15468),
.Y(n_15561)
);

INVx2_ASAP7_75t_L g15562 ( 
.A(n_15377),
.Y(n_15562)
);

INVx1_ASAP7_75t_L g15563 ( 
.A(n_15410),
.Y(n_15563)
);

AND2x4_ASAP7_75t_L g15564 ( 
.A(n_15317),
.B(n_15247),
.Y(n_15564)
);

INVx1_ASAP7_75t_L g15565 ( 
.A(n_15414),
.Y(n_15565)
);

AND2x2_ASAP7_75t_L g15566 ( 
.A(n_15300),
.B(n_15250),
.Y(n_15566)
);

INVx2_ASAP7_75t_L g15567 ( 
.A(n_15431),
.Y(n_15567)
);

INVx2_ASAP7_75t_L g15568 ( 
.A(n_15321),
.Y(n_15568)
);

INVx2_ASAP7_75t_L g15569 ( 
.A(n_15475),
.Y(n_15569)
);

INVx2_ASAP7_75t_L g15570 ( 
.A(n_15430),
.Y(n_15570)
);

NAND2xp5_ASAP7_75t_L g15571 ( 
.A(n_15450),
.B(n_15094),
.Y(n_15571)
);

BUFx2_ASAP7_75t_L g15572 ( 
.A(n_15327),
.Y(n_15572)
);

AND2x2_ASAP7_75t_L g15573 ( 
.A(n_15342),
.B(n_15255),
.Y(n_15573)
);

INVx2_ASAP7_75t_L g15574 ( 
.A(n_15447),
.Y(n_15574)
);

AND2x2_ASAP7_75t_L g15575 ( 
.A(n_15448),
.B(n_15260),
.Y(n_15575)
);

INVx2_ASAP7_75t_L g15576 ( 
.A(n_15362),
.Y(n_15576)
);

AND2x2_ASAP7_75t_L g15577 ( 
.A(n_15302),
.B(n_15134),
.Y(n_15577)
);

INVx1_ASAP7_75t_L g15578 ( 
.A(n_15432),
.Y(n_15578)
);

INVx3_ASAP7_75t_L g15579 ( 
.A(n_15299),
.Y(n_15579)
);

INVx1_ASAP7_75t_L g15580 ( 
.A(n_15453),
.Y(n_15580)
);

INVx1_ASAP7_75t_L g15581 ( 
.A(n_15320),
.Y(n_15581)
);

HB1xp67_ASAP7_75t_L g15582 ( 
.A(n_15415),
.Y(n_15582)
);

OA21x2_ASAP7_75t_L g15583 ( 
.A1(n_15346),
.A2(n_15134),
.B(n_15254),
.Y(n_15583)
);

HB1xp67_ASAP7_75t_L g15584 ( 
.A(n_15471),
.Y(n_15584)
);

AND2x4_ASAP7_75t_L g15585 ( 
.A(n_15417),
.B(n_15261),
.Y(n_15585)
);

INVx3_ASAP7_75t_L g15586 ( 
.A(n_15312),
.Y(n_15586)
);

INVx2_ASAP7_75t_L g15587 ( 
.A(n_15419),
.Y(n_15587)
);

INVx2_ASAP7_75t_SL g15588 ( 
.A(n_15441),
.Y(n_15588)
);

AND2x4_ASAP7_75t_L g15589 ( 
.A(n_15388),
.B(n_15261),
.Y(n_15589)
);

HB1xp67_ASAP7_75t_L g15590 ( 
.A(n_15347),
.Y(n_15590)
);

INVx2_ASAP7_75t_L g15591 ( 
.A(n_15341),
.Y(n_15591)
);

INVx2_ASAP7_75t_L g15592 ( 
.A(n_15324),
.Y(n_15592)
);

AND2x2_ASAP7_75t_L g15593 ( 
.A(n_15307),
.B(n_15254),
.Y(n_15593)
);

INVx1_ASAP7_75t_L g15594 ( 
.A(n_15439),
.Y(n_15594)
);

AND2x2_ASAP7_75t_L g15595 ( 
.A(n_15327),
.B(n_2513),
.Y(n_15595)
);

NOR2x1_ASAP7_75t_L g15596 ( 
.A(n_15426),
.B(n_2514),
.Y(n_15596)
);

NAND2xp5_ASAP7_75t_L g15597 ( 
.A(n_15398),
.B(n_15457),
.Y(n_15597)
);

INVx3_ASAP7_75t_L g15598 ( 
.A(n_15331),
.Y(n_15598)
);

OA21x2_ASAP7_75t_L g15599 ( 
.A1(n_15294),
.A2(n_15359),
.B(n_15340),
.Y(n_15599)
);

INVx2_ASAP7_75t_L g15600 ( 
.A(n_15452),
.Y(n_15600)
);

INVx2_ASAP7_75t_L g15601 ( 
.A(n_15372),
.Y(n_15601)
);

AND2x4_ASAP7_75t_L g15602 ( 
.A(n_15369),
.B(n_15323),
.Y(n_15602)
);

OAI221xp5_ASAP7_75t_L g15603 ( 
.A1(n_15326),
.A2(n_2517),
.B1(n_2515),
.B2(n_2516),
.C(n_2518),
.Y(n_15603)
);

AOI22xp33_ASAP7_75t_L g15604 ( 
.A1(n_15310),
.A2(n_15476),
.B1(n_15485),
.B2(n_15301),
.Y(n_15604)
);

INVx1_ASAP7_75t_L g15605 ( 
.A(n_15445),
.Y(n_15605)
);

INVx2_ASAP7_75t_L g15606 ( 
.A(n_15422),
.Y(n_15606)
);

AND2x2_ASAP7_75t_L g15607 ( 
.A(n_15393),
.B(n_15353),
.Y(n_15607)
);

INVx1_ASAP7_75t_L g15608 ( 
.A(n_15456),
.Y(n_15608)
);

INVx2_ASAP7_75t_L g15609 ( 
.A(n_15396),
.Y(n_15609)
);

AND2x2_ASAP7_75t_L g15610 ( 
.A(n_15328),
.B(n_15348),
.Y(n_15610)
);

AND2x2_ASAP7_75t_L g15611 ( 
.A(n_15429),
.B(n_2518),
.Y(n_15611)
);

INVx2_ASAP7_75t_L g15612 ( 
.A(n_15408),
.Y(n_15612)
);

OR2x2_ASAP7_75t_L g15613 ( 
.A(n_15395),
.B(n_2519),
.Y(n_15613)
);

HB1xp67_ASAP7_75t_L g15614 ( 
.A(n_15298),
.Y(n_15614)
);

INVx1_ASAP7_75t_L g15615 ( 
.A(n_15443),
.Y(n_15615)
);

AOI22xp5_ASAP7_75t_L g15616 ( 
.A1(n_15343),
.A2(n_2522),
.B1(n_2520),
.B2(n_2521),
.Y(n_15616)
);

AND2x2_ASAP7_75t_L g15617 ( 
.A(n_15319),
.B(n_15303),
.Y(n_15617)
);

AND2x2_ASAP7_75t_L g15618 ( 
.A(n_15374),
.B(n_2521),
.Y(n_15618)
);

OR2x2_ASAP7_75t_L g15619 ( 
.A(n_15339),
.B(n_2522),
.Y(n_15619)
);

OR2x2_ASAP7_75t_L g15620 ( 
.A(n_15355),
.B(n_2524),
.Y(n_15620)
);

OR2x2_ASAP7_75t_L g15621 ( 
.A(n_15486),
.B(n_2524),
.Y(n_15621)
);

AND2x2_ASAP7_75t_L g15622 ( 
.A(n_15491),
.B(n_2525),
.Y(n_15622)
);

NAND2xp5_ASAP7_75t_L g15623 ( 
.A(n_15455),
.B(n_15397),
.Y(n_15623)
);

INVxp67_ASAP7_75t_L g15624 ( 
.A(n_15421),
.Y(n_15624)
);

INVx1_ASAP7_75t_L g15625 ( 
.A(n_15444),
.Y(n_15625)
);

INVx3_ASAP7_75t_L g15626 ( 
.A(n_15338),
.Y(n_15626)
);

NAND2xp5_ASAP7_75t_L g15627 ( 
.A(n_15306),
.B(n_2525),
.Y(n_15627)
);

INVx1_ASAP7_75t_L g15628 ( 
.A(n_15451),
.Y(n_15628)
);

INVx1_ASAP7_75t_L g15629 ( 
.A(n_15438),
.Y(n_15629)
);

NAND2xp5_ASAP7_75t_L g15630 ( 
.A(n_15390),
.B(n_2526),
.Y(n_15630)
);

NAND2xp5_ASAP7_75t_L g15631 ( 
.A(n_15411),
.B(n_2526),
.Y(n_15631)
);

OAI21xp33_ASAP7_75t_L g15632 ( 
.A1(n_15358),
.A2(n_2527),
.B(n_2528),
.Y(n_15632)
);

INVx2_ASAP7_75t_L g15633 ( 
.A(n_15473),
.Y(n_15633)
);

INVx1_ASAP7_75t_L g15634 ( 
.A(n_15394),
.Y(n_15634)
);

BUFx6f_ASAP7_75t_L g15635 ( 
.A(n_15424),
.Y(n_15635)
);

BUFx3_ASAP7_75t_L g15636 ( 
.A(n_15379),
.Y(n_15636)
);

AND2x2_ASAP7_75t_L g15637 ( 
.A(n_15413),
.B(n_2527),
.Y(n_15637)
);

INVx4_ASAP7_75t_R g15638 ( 
.A(n_15467),
.Y(n_15638)
);

INVx1_ASAP7_75t_L g15639 ( 
.A(n_15404),
.Y(n_15639)
);

HB1xp67_ASAP7_75t_L g15640 ( 
.A(n_15401),
.Y(n_15640)
);

INVx1_ASAP7_75t_L g15641 ( 
.A(n_15364),
.Y(n_15641)
);

NAND2xp5_ASAP7_75t_L g15642 ( 
.A(n_15436),
.B(n_2528),
.Y(n_15642)
);

AOI22xp33_ASAP7_75t_L g15643 ( 
.A1(n_15325),
.A2(n_2531),
.B1(n_2529),
.B2(n_2530),
.Y(n_15643)
);

NAND2xp5_ASAP7_75t_L g15644 ( 
.A(n_15356),
.B(n_2529),
.Y(n_15644)
);

OR2x2_ASAP7_75t_L g15645 ( 
.A(n_15337),
.B(n_2530),
.Y(n_15645)
);

INVx2_ASAP7_75t_L g15646 ( 
.A(n_15482),
.Y(n_15646)
);

AND2x2_ASAP7_75t_L g15647 ( 
.A(n_15413),
.B(n_2531),
.Y(n_15647)
);

INVx1_ASAP7_75t_L g15648 ( 
.A(n_15434),
.Y(n_15648)
);

NAND2xp5_ASAP7_75t_L g15649 ( 
.A(n_15472),
.B(n_15386),
.Y(n_15649)
);

INVx1_ASAP7_75t_L g15650 ( 
.A(n_15371),
.Y(n_15650)
);

INVx1_ASAP7_75t_L g15651 ( 
.A(n_15371),
.Y(n_15651)
);

OAI221xp5_ASAP7_75t_SL g15652 ( 
.A1(n_15514),
.A2(n_15446),
.B1(n_15387),
.B2(n_15370),
.C(n_15440),
.Y(n_15652)
);

NAND2xp5_ASAP7_75t_L g15653 ( 
.A(n_15506),
.B(n_15489),
.Y(n_15653)
);

AOI21xp5_ASAP7_75t_SL g15654 ( 
.A1(n_15637),
.A2(n_15490),
.B(n_15418),
.Y(n_15654)
);

AND2x2_ASAP7_75t_L g15655 ( 
.A(n_15507),
.B(n_15487),
.Y(n_15655)
);

NAND2xp5_ASAP7_75t_SL g15656 ( 
.A(n_15635),
.B(n_15322),
.Y(n_15656)
);

AND2x2_ASAP7_75t_L g15657 ( 
.A(n_15517),
.B(n_15488),
.Y(n_15657)
);

AND2x2_ASAP7_75t_L g15658 ( 
.A(n_15505),
.B(n_15333),
.Y(n_15658)
);

NAND2xp5_ASAP7_75t_L g15659 ( 
.A(n_15584),
.B(n_15478),
.Y(n_15659)
);

AND2x2_ASAP7_75t_SL g15660 ( 
.A(n_15647),
.B(n_15466),
.Y(n_15660)
);

AOI22xp33_ASAP7_75t_L g15661 ( 
.A1(n_15599),
.A2(n_15376),
.B1(n_15454),
.B2(n_15409),
.Y(n_15661)
);

NAND2xp5_ASAP7_75t_L g15662 ( 
.A(n_15544),
.B(n_15470),
.Y(n_15662)
);

NAND2xp5_ASAP7_75t_L g15663 ( 
.A(n_15499),
.B(n_15477),
.Y(n_15663)
);

AOI22xp33_ASAP7_75t_L g15664 ( 
.A1(n_15649),
.A2(n_15474),
.B1(n_15480),
.B2(n_15479),
.Y(n_15664)
);

OAI21xp33_ASAP7_75t_L g15665 ( 
.A1(n_15604),
.A2(n_15383),
.B(n_15449),
.Y(n_15665)
);

AND2x2_ASAP7_75t_L g15666 ( 
.A(n_15510),
.B(n_15548),
.Y(n_15666)
);

AND2x2_ASAP7_75t_L g15667 ( 
.A(n_15532),
.B(n_15333),
.Y(n_15667)
);

AND2x2_ASAP7_75t_L g15668 ( 
.A(n_15572),
.B(n_15493),
.Y(n_15668)
);

NAND2xp5_ASAP7_75t_L g15669 ( 
.A(n_15500),
.B(n_15579),
.Y(n_15669)
);

NAND2xp5_ASAP7_75t_L g15670 ( 
.A(n_15650),
.B(n_15484),
.Y(n_15670)
);

NAND2xp5_ASAP7_75t_L g15671 ( 
.A(n_15651),
.B(n_15368),
.Y(n_15671)
);

AOI22xp33_ASAP7_75t_SL g15672 ( 
.A1(n_15640),
.A2(n_15392),
.B1(n_15469),
.B2(n_15460),
.Y(n_15672)
);

NAND3xp33_ASAP7_75t_L g15673 ( 
.A(n_15554),
.B(n_15416),
.C(n_15425),
.Y(n_15673)
);

AND2x2_ASAP7_75t_L g15674 ( 
.A(n_15540),
.B(n_15313),
.Y(n_15674)
);

AOI22xp5_ASAP7_75t_L g15675 ( 
.A1(n_15496),
.A2(n_15313),
.B1(n_15375),
.B2(n_15494),
.Y(n_15675)
);

NAND2xp5_ASAP7_75t_L g15676 ( 
.A(n_15570),
.B(n_15375),
.Y(n_15676)
);

NOR3xp33_ASAP7_75t_SL g15677 ( 
.A(n_15603),
.B(n_15495),
.C(n_15571),
.Y(n_15677)
);

NAND2xp5_ASAP7_75t_L g15678 ( 
.A(n_15557),
.B(n_15494),
.Y(n_15678)
);

NOR2xp33_ASAP7_75t_L g15679 ( 
.A(n_15574),
.B(n_2532),
.Y(n_15679)
);

AND2x2_ASAP7_75t_SL g15680 ( 
.A(n_15549),
.B(n_2532),
.Y(n_15680)
);

OAI21xp5_ASAP7_75t_SL g15681 ( 
.A1(n_15542),
.A2(n_2533),
.B(n_2534),
.Y(n_15681)
);

NAND3xp33_ASAP7_75t_L g15682 ( 
.A(n_15558),
.B(n_2533),
.C(n_2534),
.Y(n_15682)
);

NAND2xp5_ASAP7_75t_SL g15683 ( 
.A(n_15635),
.B(n_2535),
.Y(n_15683)
);

NAND3xp33_ASAP7_75t_L g15684 ( 
.A(n_15590),
.B(n_15644),
.C(n_15627),
.Y(n_15684)
);

OAI21xp5_ASAP7_75t_SL g15685 ( 
.A1(n_15643),
.A2(n_2535),
.B(n_2536),
.Y(n_15685)
);

NAND2xp5_ASAP7_75t_L g15686 ( 
.A(n_15588),
.B(n_2536),
.Y(n_15686)
);

AND2x2_ASAP7_75t_L g15687 ( 
.A(n_15586),
.B(n_2537),
.Y(n_15687)
);

NAND4xp25_ASAP7_75t_SL g15688 ( 
.A(n_15552),
.B(n_2539),
.C(n_2537),
.D(n_2538),
.Y(n_15688)
);

NAND2xp5_ASAP7_75t_L g15689 ( 
.A(n_15598),
.B(n_2538),
.Y(n_15689)
);

AND2x2_ASAP7_75t_L g15690 ( 
.A(n_15531),
.B(n_2539),
.Y(n_15690)
);

AND2x2_ASAP7_75t_L g15691 ( 
.A(n_15541),
.B(n_2540),
.Y(n_15691)
);

NAND2xp5_ASAP7_75t_L g15692 ( 
.A(n_15569),
.B(n_2540),
.Y(n_15692)
);

AND2x2_ASAP7_75t_L g15693 ( 
.A(n_15567),
.B(n_2541),
.Y(n_15693)
);

NAND2xp33_ASAP7_75t_R g15694 ( 
.A(n_15515),
.B(n_2541),
.Y(n_15694)
);

NAND2xp5_ASAP7_75t_L g15695 ( 
.A(n_15614),
.B(n_2542),
.Y(n_15695)
);

INVx1_ASAP7_75t_L g15696 ( 
.A(n_15582),
.Y(n_15696)
);

OAI22xp5_ASAP7_75t_L g15697 ( 
.A1(n_15624),
.A2(n_2546),
.B1(n_2543),
.B2(n_2545),
.Y(n_15697)
);

NAND4xp25_ASAP7_75t_L g15698 ( 
.A(n_15508),
.B(n_2546),
.C(n_2543),
.D(n_2545),
.Y(n_15698)
);

AND2x2_ASAP7_75t_L g15699 ( 
.A(n_15504),
.B(n_2547),
.Y(n_15699)
);

AND2x2_ASAP7_75t_L g15700 ( 
.A(n_15519),
.B(n_2548),
.Y(n_15700)
);

AND2x2_ASAP7_75t_L g15701 ( 
.A(n_15497),
.B(n_2548),
.Y(n_15701)
);

AND2x2_ASAP7_75t_L g15702 ( 
.A(n_15610),
.B(n_2549),
.Y(n_15702)
);

AND2x2_ASAP7_75t_L g15703 ( 
.A(n_15592),
.B(n_2550),
.Y(n_15703)
);

NAND2xp5_ASAP7_75t_L g15704 ( 
.A(n_15528),
.B(n_2550),
.Y(n_15704)
);

OAI21xp5_ASAP7_75t_SL g15705 ( 
.A1(n_15596),
.A2(n_2551),
.B(n_2552),
.Y(n_15705)
);

NAND2xp5_ASAP7_75t_L g15706 ( 
.A(n_15626),
.B(n_2551),
.Y(n_15706)
);

AND2x2_ASAP7_75t_L g15707 ( 
.A(n_15537),
.B(n_2552),
.Y(n_15707)
);

AND2x2_ASAP7_75t_L g15708 ( 
.A(n_15512),
.B(n_2553),
.Y(n_15708)
);

OAI22xp5_ASAP7_75t_L g15709 ( 
.A1(n_15521),
.A2(n_2555),
.B1(n_2553),
.B2(n_2554),
.Y(n_15709)
);

AND2x2_ASAP7_75t_L g15710 ( 
.A(n_15607),
.B(n_2554),
.Y(n_15710)
);

NAND3xp33_ASAP7_75t_L g15711 ( 
.A(n_15583),
.B(n_2555),
.C(n_2556),
.Y(n_15711)
);

AND2x2_ASAP7_75t_SL g15712 ( 
.A(n_15529),
.B(n_2556),
.Y(n_15712)
);

NAND2xp5_ASAP7_75t_L g15713 ( 
.A(n_15577),
.B(n_2557),
.Y(n_15713)
);

NAND2xp5_ASAP7_75t_L g15714 ( 
.A(n_15581),
.B(n_2557),
.Y(n_15714)
);

OAI21xp33_ASAP7_75t_L g15715 ( 
.A1(n_15538),
.A2(n_2558),
.B(n_2559),
.Y(n_15715)
);

NAND3xp33_ASAP7_75t_L g15716 ( 
.A(n_15525),
.B(n_2558),
.C(n_2559),
.Y(n_15716)
);

AND2x2_ASAP7_75t_L g15717 ( 
.A(n_15498),
.B(n_2560),
.Y(n_15717)
);

AOI221xp5_ASAP7_75t_L g15718 ( 
.A1(n_15550),
.A2(n_15632),
.B1(n_15533),
.B2(n_15509),
.C(n_15523),
.Y(n_15718)
);

NAND2xp5_ASAP7_75t_L g15719 ( 
.A(n_15595),
.B(n_2560),
.Y(n_15719)
);

AND2x2_ASAP7_75t_L g15720 ( 
.A(n_15602),
.B(n_2561),
.Y(n_15720)
);

AND2x2_ASAP7_75t_L g15721 ( 
.A(n_15591),
.B(n_2561),
.Y(n_15721)
);

OAI22xp5_ASAP7_75t_L g15722 ( 
.A1(n_15597),
.A2(n_2564),
.B1(n_2562),
.B2(n_2563),
.Y(n_15722)
);

NAND3xp33_ASAP7_75t_L g15723 ( 
.A(n_15645),
.B(n_2562),
.C(n_2563),
.Y(n_15723)
);

AOI211xp5_ASAP7_75t_L g15724 ( 
.A1(n_15539),
.A2(n_2566),
.B(n_2564),
.C(n_2565),
.Y(n_15724)
);

NAND2xp5_ASAP7_75t_L g15725 ( 
.A(n_15593),
.B(n_2565),
.Y(n_15725)
);

NAND2xp5_ASAP7_75t_L g15726 ( 
.A(n_15551),
.B(n_2566),
.Y(n_15726)
);

NAND2xp5_ASAP7_75t_L g15727 ( 
.A(n_15562),
.B(n_2567),
.Y(n_15727)
);

NAND2xp5_ASAP7_75t_L g15728 ( 
.A(n_15612),
.B(n_2567),
.Y(n_15728)
);

OAI21xp5_ASAP7_75t_SL g15729 ( 
.A1(n_15623),
.A2(n_2568),
.B(n_2570),
.Y(n_15729)
);

AOI22xp33_ASAP7_75t_L g15730 ( 
.A1(n_15568),
.A2(n_2571),
.B1(n_2568),
.B2(n_2570),
.Y(n_15730)
);

OAI21xp5_ASAP7_75t_L g15731 ( 
.A1(n_15559),
.A2(n_15631),
.B(n_15630),
.Y(n_15731)
);

NAND2xp5_ASAP7_75t_L g15732 ( 
.A(n_15601),
.B(n_2571),
.Y(n_15732)
);

NAND4xp25_ASAP7_75t_L g15733 ( 
.A(n_15617),
.B(n_2574),
.C(n_2572),
.D(n_2573),
.Y(n_15733)
);

NAND2xp5_ASAP7_75t_SL g15734 ( 
.A(n_15606),
.B(n_2572),
.Y(n_15734)
);

NAND3xp33_ASAP7_75t_L g15735 ( 
.A(n_15555),
.B(n_2574),
.C(n_2575),
.Y(n_15735)
);

INVx3_ASAP7_75t_L g15736 ( 
.A(n_15636),
.Y(n_15736)
);

NAND2xp5_ASAP7_75t_SL g15737 ( 
.A(n_15609),
.B(n_2576),
.Y(n_15737)
);

AND2x2_ASAP7_75t_L g15738 ( 
.A(n_15543),
.B(n_2576),
.Y(n_15738)
);

AND2x2_ASAP7_75t_L g15739 ( 
.A(n_15633),
.B(n_2577),
.Y(n_15739)
);

AOI211xp5_ASAP7_75t_SL g15740 ( 
.A1(n_15503),
.A2(n_2580),
.B(n_2577),
.C(n_2578),
.Y(n_15740)
);

AND2x2_ASAP7_75t_L g15741 ( 
.A(n_15646),
.B(n_2580),
.Y(n_15741)
);

AND2x2_ASAP7_75t_L g15742 ( 
.A(n_15600),
.B(n_2581),
.Y(n_15742)
);

AND2x2_ASAP7_75t_L g15743 ( 
.A(n_15573),
.B(n_15566),
.Y(n_15743)
);

NAND3xp33_ASAP7_75t_L g15744 ( 
.A(n_15511),
.B(n_2581),
.C(n_2582),
.Y(n_15744)
);

AND2x2_ASAP7_75t_L g15745 ( 
.A(n_15576),
.B(n_2583),
.Y(n_15745)
);

NAND2xp5_ASAP7_75t_L g15746 ( 
.A(n_15634),
.B(n_2584),
.Y(n_15746)
);

OAI21xp33_ASAP7_75t_L g15747 ( 
.A1(n_15648),
.A2(n_2584),
.B(n_2585),
.Y(n_15747)
);

NAND2xp5_ASAP7_75t_SL g15748 ( 
.A(n_15589),
.B(n_2585),
.Y(n_15748)
);

AND2x2_ASAP7_75t_L g15749 ( 
.A(n_15587),
.B(n_2586),
.Y(n_15749)
);

AND2x2_ASAP7_75t_L g15750 ( 
.A(n_15639),
.B(n_2587),
.Y(n_15750)
);

NAND2xp5_ASAP7_75t_L g15751 ( 
.A(n_15629),
.B(n_2588),
.Y(n_15751)
);

AND2x2_ASAP7_75t_SL g15752 ( 
.A(n_15527),
.B(n_2588),
.Y(n_15752)
);

INVx1_ASAP7_75t_L g15753 ( 
.A(n_15524),
.Y(n_15753)
);

NAND3xp33_ASAP7_75t_L g15754 ( 
.A(n_15501),
.B(n_15530),
.C(n_15502),
.Y(n_15754)
);

NAND2xp5_ASAP7_75t_L g15755 ( 
.A(n_15608),
.B(n_2589),
.Y(n_15755)
);

AND2x2_ASAP7_75t_L g15756 ( 
.A(n_15615),
.B(n_2590),
.Y(n_15756)
);

AND2x2_ASAP7_75t_L g15757 ( 
.A(n_15625),
.B(n_2590),
.Y(n_15757)
);

AND2x2_ASAP7_75t_L g15758 ( 
.A(n_15628),
.B(n_2591),
.Y(n_15758)
);

OAI22xp33_ASAP7_75t_SL g15759 ( 
.A1(n_15516),
.A2(n_2594),
.B1(n_2592),
.B2(n_2593),
.Y(n_15759)
);

AOI22xp33_ASAP7_75t_SL g15760 ( 
.A1(n_15518),
.A2(n_2594),
.B1(n_2592),
.B2(n_2593),
.Y(n_15760)
);

NAND4xp25_ASAP7_75t_L g15761 ( 
.A(n_15522),
.B(n_2597),
.C(n_2595),
.D(n_2596),
.Y(n_15761)
);

OAI21xp5_ASAP7_75t_L g15762 ( 
.A1(n_15642),
.A2(n_2595),
.B(n_2596),
.Y(n_15762)
);

OAI211xp5_ASAP7_75t_L g15763 ( 
.A1(n_15534),
.A2(n_2599),
.B(n_2597),
.C(n_2598),
.Y(n_15763)
);

OAI22xp5_ASAP7_75t_L g15764 ( 
.A1(n_15616),
.A2(n_2600),
.B1(n_2598),
.B2(n_2599),
.Y(n_15764)
);

AOI21xp33_ASAP7_75t_SL g15765 ( 
.A1(n_15526),
.A2(n_2600),
.B(n_2601),
.Y(n_15765)
);

NAND3xp33_ASAP7_75t_L g15766 ( 
.A(n_15520),
.B(n_2601),
.C(n_2602),
.Y(n_15766)
);

OAI22xp5_ASAP7_75t_L g15767 ( 
.A1(n_15560),
.A2(n_2604),
.B1(n_2602),
.B2(n_2603),
.Y(n_15767)
);

NOR3xp33_ASAP7_75t_L g15768 ( 
.A(n_15545),
.B(n_2603),
.C(n_2604),
.Y(n_15768)
);

OAI221xp5_ASAP7_75t_SL g15769 ( 
.A1(n_15513),
.A2(n_2607),
.B1(n_2605),
.B2(n_2606),
.C(n_2608),
.Y(n_15769)
);

OAI221xp5_ASAP7_75t_SL g15770 ( 
.A1(n_15546),
.A2(n_2609),
.B1(n_2605),
.B2(n_2607),
.C(n_2610),
.Y(n_15770)
);

NOR3xp33_ASAP7_75t_L g15771 ( 
.A(n_15563),
.B(n_2609),
.C(n_2610),
.Y(n_15771)
);

AND2x2_ASAP7_75t_L g15772 ( 
.A(n_15575),
.B(n_2611),
.Y(n_15772)
);

OAI21xp5_ASAP7_75t_SL g15773 ( 
.A1(n_15561),
.A2(n_2611),
.B(n_2612),
.Y(n_15773)
);

NAND2xp33_ASAP7_75t_SL g15774 ( 
.A(n_15556),
.B(n_2612),
.Y(n_15774)
);

OAI22xp5_ASAP7_75t_L g15775 ( 
.A1(n_15641),
.A2(n_2615),
.B1(n_2613),
.B2(n_2614),
.Y(n_15775)
);

NAND2xp5_ASAP7_75t_L g15776 ( 
.A(n_15564),
.B(n_2615),
.Y(n_15776)
);

NAND2xp5_ASAP7_75t_L g15777 ( 
.A(n_15622),
.B(n_2616),
.Y(n_15777)
);

NAND3xp33_ASAP7_75t_L g15778 ( 
.A(n_15535),
.B(n_2616),
.C(n_2617),
.Y(n_15778)
);

OAI221xp5_ASAP7_75t_SL g15779 ( 
.A1(n_15553),
.A2(n_15605),
.B1(n_15580),
.B2(n_15565),
.C(n_15578),
.Y(n_15779)
);

OAI21xp5_ASAP7_75t_SL g15780 ( 
.A1(n_15547),
.A2(n_15594),
.B(n_15536),
.Y(n_15780)
);

NAND3xp33_ASAP7_75t_L g15781 ( 
.A(n_15619),
.B(n_2617),
.C(n_2618),
.Y(n_15781)
);

NAND2xp5_ASAP7_75t_L g15782 ( 
.A(n_15611),
.B(n_2618),
.Y(n_15782)
);

NAND2xp5_ASAP7_75t_L g15783 ( 
.A(n_15585),
.B(n_2619),
.Y(n_15783)
);

AND2x2_ASAP7_75t_L g15784 ( 
.A(n_15618),
.B(n_2619),
.Y(n_15784)
);

HB1xp67_ASAP7_75t_L g15785 ( 
.A(n_15680),
.Y(n_15785)
);

AND2x2_ASAP7_75t_L g15786 ( 
.A(n_15660),
.B(n_15620),
.Y(n_15786)
);

OAI21x1_ASAP7_75t_L g15787 ( 
.A1(n_15678),
.A2(n_15613),
.B(n_15621),
.Y(n_15787)
);

OAI21xp5_ASAP7_75t_L g15788 ( 
.A1(n_15673),
.A2(n_15638),
.B(n_2620),
.Y(n_15788)
);

HB1xp67_ASAP7_75t_L g15789 ( 
.A(n_15743),
.Y(n_15789)
);

INVx1_ASAP7_75t_L g15790 ( 
.A(n_15690),
.Y(n_15790)
);

NOR2xp33_ASAP7_75t_L g15791 ( 
.A(n_15666),
.B(n_2620),
.Y(n_15791)
);

INVx2_ASAP7_75t_L g15792 ( 
.A(n_15655),
.Y(n_15792)
);

INVx1_ASAP7_75t_L g15793 ( 
.A(n_15668),
.Y(n_15793)
);

OR2x2_ASAP7_75t_L g15794 ( 
.A(n_15676),
.B(n_2621),
.Y(n_15794)
);

OAI21x1_ASAP7_75t_L g15795 ( 
.A1(n_15748),
.A2(n_2621),
.B(n_2622),
.Y(n_15795)
);

INVx2_ASAP7_75t_L g15796 ( 
.A(n_15657),
.Y(n_15796)
);

INVx3_ASAP7_75t_L g15797 ( 
.A(n_15736),
.Y(n_15797)
);

CKINVDCx5p33_ASAP7_75t_R g15798 ( 
.A(n_15712),
.Y(n_15798)
);

NAND2xp5_ASAP7_75t_L g15799 ( 
.A(n_15667),
.B(n_2622),
.Y(n_15799)
);

BUFx12f_ASAP7_75t_L g15800 ( 
.A(n_15691),
.Y(n_15800)
);

HB1xp67_ASAP7_75t_L g15801 ( 
.A(n_15694),
.Y(n_15801)
);

A2O1A1Ixp33_ASAP7_75t_L g15802 ( 
.A1(n_15675),
.A2(n_2625),
.B(n_2623),
.C(n_2624),
.Y(n_15802)
);

INVx1_ASAP7_75t_L g15803 ( 
.A(n_15708),
.Y(n_15803)
);

INVx2_ASAP7_75t_L g15804 ( 
.A(n_15687),
.Y(n_15804)
);

INVx1_ASAP7_75t_L g15805 ( 
.A(n_15700),
.Y(n_15805)
);

INVx1_ASAP7_75t_L g15806 ( 
.A(n_15702),
.Y(n_15806)
);

OR2x6_ASAP7_75t_L g15807 ( 
.A(n_15669),
.B(n_2623),
.Y(n_15807)
);

INVx1_ASAP7_75t_L g15808 ( 
.A(n_15701),
.Y(n_15808)
);

INVx1_ASAP7_75t_L g15809 ( 
.A(n_15686),
.Y(n_15809)
);

INVx1_ASAP7_75t_L g15810 ( 
.A(n_15692),
.Y(n_15810)
);

BUFx3_ASAP7_75t_L g15811 ( 
.A(n_15699),
.Y(n_15811)
);

OA21x2_ASAP7_75t_L g15812 ( 
.A1(n_15711),
.A2(n_2624),
.B(n_2625),
.Y(n_15812)
);

BUFx3_ASAP7_75t_L g15813 ( 
.A(n_15693),
.Y(n_15813)
);

INVx1_ASAP7_75t_L g15814 ( 
.A(n_15696),
.Y(n_15814)
);

NAND2xp5_ASAP7_75t_SL g15815 ( 
.A(n_15752),
.B(n_2626),
.Y(n_15815)
);

INVx2_ASAP7_75t_L g15816 ( 
.A(n_15710),
.Y(n_15816)
);

OR2x2_ASAP7_75t_L g15817 ( 
.A(n_15671),
.B(n_2627),
.Y(n_15817)
);

AOI22xp5_ASAP7_75t_L g15818 ( 
.A1(n_15665),
.A2(n_2630),
.B1(n_2627),
.B2(n_2629),
.Y(n_15818)
);

INVx5_ASAP7_75t_L g15819 ( 
.A(n_15707),
.Y(n_15819)
);

AO21x2_ASAP7_75t_L g15820 ( 
.A1(n_15713),
.A2(n_2630),
.B(n_2631),
.Y(n_15820)
);

INVx2_ASAP7_75t_SL g15821 ( 
.A(n_15720),
.Y(n_15821)
);

INVx1_ASAP7_75t_L g15822 ( 
.A(n_15739),
.Y(n_15822)
);

INVx2_ASAP7_75t_L g15823 ( 
.A(n_15717),
.Y(n_15823)
);

AND2x2_ASAP7_75t_L g15824 ( 
.A(n_15658),
.B(n_2631),
.Y(n_15824)
);

AND2x2_ASAP7_75t_L g15825 ( 
.A(n_15674),
.B(n_2632),
.Y(n_15825)
);

A2O1A1Ixp33_ASAP7_75t_L g15826 ( 
.A1(n_15652),
.A2(n_2635),
.B(n_2632),
.C(n_2634),
.Y(n_15826)
);

INVx2_ASAP7_75t_L g15827 ( 
.A(n_15784),
.Y(n_15827)
);

OA21x2_ASAP7_75t_L g15828 ( 
.A1(n_15661),
.A2(n_2634),
.B(n_2636),
.Y(n_15828)
);

INVx2_ASAP7_75t_SL g15829 ( 
.A(n_15738),
.Y(n_15829)
);

INVx1_ASAP7_75t_L g15830 ( 
.A(n_15741),
.Y(n_15830)
);

INVx2_ASAP7_75t_L g15831 ( 
.A(n_15772),
.Y(n_15831)
);

NOR2xp33_ASAP7_75t_R g15832 ( 
.A(n_15774),
.B(n_2636),
.Y(n_15832)
);

OAI21x1_ASAP7_75t_L g15833 ( 
.A1(n_15731),
.A2(n_2637),
.B(n_2638),
.Y(n_15833)
);

INVx2_ASAP7_75t_L g15834 ( 
.A(n_15703),
.Y(n_15834)
);

INVx1_ASAP7_75t_L g15835 ( 
.A(n_15753),
.Y(n_15835)
);

NAND2xp5_ASAP7_75t_L g15836 ( 
.A(n_15740),
.B(n_2637),
.Y(n_15836)
);

INVx2_ASAP7_75t_L g15837 ( 
.A(n_15756),
.Y(n_15837)
);

INVx2_ASAP7_75t_L g15838 ( 
.A(n_15757),
.Y(n_15838)
);

INVx2_ASAP7_75t_L g15839 ( 
.A(n_15758),
.Y(n_15839)
);

INVx6_ASAP7_75t_L g15840 ( 
.A(n_15745),
.Y(n_15840)
);

AND2x2_ASAP7_75t_L g15841 ( 
.A(n_15750),
.B(n_2638),
.Y(n_15841)
);

INVx2_ASAP7_75t_L g15842 ( 
.A(n_15742),
.Y(n_15842)
);

INVx1_ASAP7_75t_L g15843 ( 
.A(n_15704),
.Y(n_15843)
);

INVx2_ASAP7_75t_L g15844 ( 
.A(n_15749),
.Y(n_15844)
);

A2O1A1Ixp33_ASAP7_75t_L g15845 ( 
.A1(n_15682),
.A2(n_2641),
.B(n_2639),
.C(n_2640),
.Y(n_15845)
);

CKINVDCx5p33_ASAP7_75t_R g15846 ( 
.A(n_15759),
.Y(n_15846)
);

INVx1_ASAP7_75t_L g15847 ( 
.A(n_15663),
.Y(n_15847)
);

AND2x2_ASAP7_75t_L g15848 ( 
.A(n_15721),
.B(n_2639),
.Y(n_15848)
);

INVx1_ASAP7_75t_L g15849 ( 
.A(n_15776),
.Y(n_15849)
);

INVx1_ASAP7_75t_L g15850 ( 
.A(n_15782),
.Y(n_15850)
);

INVx2_ASAP7_75t_L g15851 ( 
.A(n_15689),
.Y(n_15851)
);

INVx2_ASAP7_75t_L g15852 ( 
.A(n_15706),
.Y(n_15852)
);

INVx2_ASAP7_75t_L g15853 ( 
.A(n_15719),
.Y(n_15853)
);

BUFx3_ASAP7_75t_L g15854 ( 
.A(n_15726),
.Y(n_15854)
);

INVx3_ASAP7_75t_L g15855 ( 
.A(n_15727),
.Y(n_15855)
);

AND2x2_ASAP7_75t_SL g15856 ( 
.A(n_15670),
.B(n_2640),
.Y(n_15856)
);

INVx1_ASAP7_75t_L g15857 ( 
.A(n_15783),
.Y(n_15857)
);

AOI21xp5_ASAP7_75t_L g15858 ( 
.A1(n_15654),
.A2(n_2641),
.B(n_2642),
.Y(n_15858)
);

AND2x2_ASAP7_75t_SL g15859 ( 
.A(n_15653),
.B(n_2642),
.Y(n_15859)
);

INVx1_ASAP7_75t_L g15860 ( 
.A(n_15695),
.Y(n_15860)
);

AND2x2_ASAP7_75t_L g15861 ( 
.A(n_15679),
.B(n_2643),
.Y(n_15861)
);

AND2x6_ASAP7_75t_L g15862 ( 
.A(n_15728),
.B(n_2643),
.Y(n_15862)
);

AOI21xp5_ASAP7_75t_L g15863 ( 
.A1(n_15656),
.A2(n_2644),
.B(n_2645),
.Y(n_15863)
);

HB1xp67_ASAP7_75t_L g15864 ( 
.A(n_15688),
.Y(n_15864)
);

INVxp67_ASAP7_75t_L g15865 ( 
.A(n_15683),
.Y(n_15865)
);

AND2x2_ASAP7_75t_L g15866 ( 
.A(n_15659),
.B(n_2644),
.Y(n_15866)
);

INVx1_ASAP7_75t_SL g15867 ( 
.A(n_15662),
.Y(n_15867)
);

INVx1_ASAP7_75t_L g15868 ( 
.A(n_15777),
.Y(n_15868)
);

OA21x2_ASAP7_75t_L g15869 ( 
.A1(n_15681),
.A2(n_2645),
.B(n_2647),
.Y(n_15869)
);

AND2x2_ASAP7_75t_L g15870 ( 
.A(n_15762),
.B(n_2647),
.Y(n_15870)
);

A2O1A1Ixp33_ASAP7_75t_L g15871 ( 
.A1(n_15724),
.A2(n_2650),
.B(n_2648),
.C(n_2649),
.Y(n_15871)
);

INVx1_ASAP7_75t_L g15872 ( 
.A(n_15732),
.Y(n_15872)
);

INVx2_ASAP7_75t_L g15873 ( 
.A(n_15746),
.Y(n_15873)
);

NAND2xp5_ASAP7_75t_L g15874 ( 
.A(n_15672),
.B(n_2648),
.Y(n_15874)
);

INVx1_ASAP7_75t_SL g15875 ( 
.A(n_15734),
.Y(n_15875)
);

INVx4_ASAP7_75t_L g15876 ( 
.A(n_15780),
.Y(n_15876)
);

O2A1O1Ixp5_ASAP7_75t_L g15877 ( 
.A1(n_15779),
.A2(n_2652),
.B(n_2649),
.C(n_2651),
.Y(n_15877)
);

INVxp67_ASAP7_75t_L g15878 ( 
.A(n_15725),
.Y(n_15878)
);

OA21x2_ASAP7_75t_L g15879 ( 
.A1(n_15705),
.A2(n_2651),
.B(n_2653),
.Y(n_15879)
);

HB1xp67_ASAP7_75t_L g15880 ( 
.A(n_15737),
.Y(n_15880)
);

INVx2_ASAP7_75t_L g15881 ( 
.A(n_15751),
.Y(n_15881)
);

NAND2xp5_ASAP7_75t_L g15882 ( 
.A(n_15765),
.B(n_2653),
.Y(n_15882)
);

BUFx2_ASAP7_75t_L g15883 ( 
.A(n_15714),
.Y(n_15883)
);

NAND4xp25_ASAP7_75t_L g15884 ( 
.A(n_15718),
.B(n_2656),
.C(n_2654),
.D(n_2655),
.Y(n_15884)
);

INVx2_ASAP7_75t_L g15885 ( 
.A(n_15755),
.Y(n_15885)
);

INVx1_ASAP7_75t_L g15886 ( 
.A(n_15754),
.Y(n_15886)
);

INVxp67_ASAP7_75t_L g15887 ( 
.A(n_15735),
.Y(n_15887)
);

NOR2xp33_ASAP7_75t_L g15888 ( 
.A(n_15729),
.B(n_2654),
.Y(n_15888)
);

NAND2xp5_ASAP7_75t_L g15889 ( 
.A(n_15773),
.B(n_2655),
.Y(n_15889)
);

INVx2_ASAP7_75t_SL g15890 ( 
.A(n_15709),
.Y(n_15890)
);

INVx2_ASAP7_75t_L g15891 ( 
.A(n_15766),
.Y(n_15891)
);

BUFx3_ASAP7_75t_L g15892 ( 
.A(n_15778),
.Y(n_15892)
);

AND2x2_ASAP7_75t_L g15893 ( 
.A(n_15677),
.B(n_2656),
.Y(n_15893)
);

BUFx3_ASAP7_75t_L g15894 ( 
.A(n_15781),
.Y(n_15894)
);

BUFx3_ASAP7_75t_L g15895 ( 
.A(n_15723),
.Y(n_15895)
);

INVx1_ASAP7_75t_L g15896 ( 
.A(n_15697),
.Y(n_15896)
);

INVxp67_ASAP7_75t_L g15897 ( 
.A(n_15716),
.Y(n_15897)
);

AND4x1_ASAP7_75t_L g15898 ( 
.A(n_15684),
.B(n_2659),
.C(n_2657),
.D(n_2658),
.Y(n_15898)
);

A2O1A1Ixp33_ASAP7_75t_L g15899 ( 
.A1(n_15685),
.A2(n_2659),
.B(n_2657),
.C(n_2658),
.Y(n_15899)
);

NAND2xp5_ASAP7_75t_SL g15900 ( 
.A(n_15760),
.B(n_2660),
.Y(n_15900)
);

AOI22xp33_ASAP7_75t_L g15901 ( 
.A1(n_15876),
.A2(n_15664),
.B1(n_15698),
.B2(n_15768),
.Y(n_15901)
);

NAND3xp33_ASAP7_75t_L g15902 ( 
.A(n_15877),
.B(n_15771),
.C(n_15763),
.Y(n_15902)
);

INVx1_ASAP7_75t_L g15903 ( 
.A(n_15789),
.Y(n_15903)
);

AO22x1_ASAP7_75t_L g15904 ( 
.A1(n_15798),
.A2(n_15722),
.B1(n_15764),
.B2(n_15775),
.Y(n_15904)
);

AND2x2_ASAP7_75t_L g15905 ( 
.A(n_15785),
.B(n_15715),
.Y(n_15905)
);

NAND3xp33_ASAP7_75t_L g15906 ( 
.A(n_15802),
.B(n_15744),
.C(n_15770),
.Y(n_15906)
);

AND2x2_ASAP7_75t_SL g15907 ( 
.A(n_15801),
.B(n_15730),
.Y(n_15907)
);

NOR3xp33_ASAP7_75t_SL g15908 ( 
.A(n_15846),
.B(n_15761),
.C(n_15733),
.Y(n_15908)
);

INVxp67_ASAP7_75t_SL g15909 ( 
.A(n_15815),
.Y(n_15909)
);

XNOR2xp5_ASAP7_75t_L g15910 ( 
.A(n_15898),
.B(n_15864),
.Y(n_15910)
);

AND2x2_ASAP7_75t_L g15911 ( 
.A(n_15792),
.B(n_15747),
.Y(n_15911)
);

AND2x2_ASAP7_75t_L g15912 ( 
.A(n_15793),
.B(n_15767),
.Y(n_15912)
);

AND2x2_ASAP7_75t_L g15913 ( 
.A(n_15786),
.B(n_15769),
.Y(n_15913)
);

INVx1_ASAP7_75t_L g15914 ( 
.A(n_15796),
.Y(n_15914)
);

AOI22xp5_ASAP7_75t_L g15915 ( 
.A1(n_15886),
.A2(n_15890),
.B1(n_15797),
.B2(n_15825),
.Y(n_15915)
);

INVx2_ASAP7_75t_L g15916 ( 
.A(n_15819),
.Y(n_15916)
);

AND2x2_ASAP7_75t_L g15917 ( 
.A(n_15811),
.B(n_2661),
.Y(n_15917)
);

NOR3xp33_ASAP7_75t_L g15918 ( 
.A(n_15788),
.B(n_2661),
.C(n_2662),
.Y(n_15918)
);

AND2x4_ASAP7_75t_L g15919 ( 
.A(n_15819),
.B(n_2662),
.Y(n_15919)
);

NAND4xp75_ASAP7_75t_L g15920 ( 
.A(n_15828),
.B(n_2665),
.C(n_2663),
.D(n_2664),
.Y(n_15920)
);

NAND2xp5_ASAP7_75t_L g15921 ( 
.A(n_15862),
.B(n_2664),
.Y(n_15921)
);

NAND3xp33_ASAP7_75t_L g15922 ( 
.A(n_15858),
.B(n_2665),
.C(n_2666),
.Y(n_15922)
);

INVx1_ASAP7_75t_L g15923 ( 
.A(n_15807),
.Y(n_15923)
);

NAND3xp33_ASAP7_75t_L g15924 ( 
.A(n_15826),
.B(n_2666),
.C(n_2667),
.Y(n_15924)
);

NAND2xp5_ASAP7_75t_L g15925 ( 
.A(n_15862),
.B(n_2667),
.Y(n_15925)
);

OAI211xp5_ASAP7_75t_L g15926 ( 
.A1(n_15874),
.A2(n_2670),
.B(n_2668),
.C(n_2669),
.Y(n_15926)
);

NAND2xp5_ASAP7_75t_L g15927 ( 
.A(n_15862),
.B(n_2668),
.Y(n_15927)
);

AND2x2_ASAP7_75t_L g15928 ( 
.A(n_15813),
.B(n_15816),
.Y(n_15928)
);

AOI22xp5_ASAP7_75t_L g15929 ( 
.A1(n_15875),
.A2(n_2671),
.B1(n_2669),
.B2(n_2670),
.Y(n_15929)
);

NAND2xp5_ASAP7_75t_L g15930 ( 
.A(n_15824),
.B(n_2672),
.Y(n_15930)
);

OR2x2_ASAP7_75t_L g15931 ( 
.A(n_15799),
.B(n_2672),
.Y(n_15931)
);

OR2x2_ASAP7_75t_L g15932 ( 
.A(n_15884),
.B(n_2673),
.Y(n_15932)
);

OAI211xp5_ASAP7_75t_SL g15933 ( 
.A1(n_15867),
.A2(n_2675),
.B(n_2673),
.C(n_2674),
.Y(n_15933)
);

NAND2xp5_ASAP7_75t_L g15934 ( 
.A(n_15856),
.B(n_2675),
.Y(n_15934)
);

NAND3xp33_ASAP7_75t_L g15935 ( 
.A(n_15893),
.B(n_2676),
.C(n_2677),
.Y(n_15935)
);

OAI211xp5_ASAP7_75t_SL g15936 ( 
.A1(n_15878),
.A2(n_2679),
.B(n_2676),
.C(n_2678),
.Y(n_15936)
);

AOI22xp33_ASAP7_75t_L g15937 ( 
.A1(n_15800),
.A2(n_2680),
.B1(n_2678),
.B2(n_2679),
.Y(n_15937)
);

AND2x2_ASAP7_75t_L g15938 ( 
.A(n_15823),
.B(n_2680),
.Y(n_15938)
);

AND2x2_ASAP7_75t_L g15939 ( 
.A(n_15827),
.B(n_2682),
.Y(n_15939)
);

OR2x2_ASAP7_75t_L g15940 ( 
.A(n_15794),
.B(n_2682),
.Y(n_15940)
);

INVx2_ASAP7_75t_L g15941 ( 
.A(n_15840),
.Y(n_15941)
);

INVxp67_ASAP7_75t_SL g15942 ( 
.A(n_15880),
.Y(n_15942)
);

NAND2xp5_ASAP7_75t_L g15943 ( 
.A(n_15859),
.B(n_2683),
.Y(n_15943)
);

AO21x2_ASAP7_75t_L g15944 ( 
.A1(n_15832),
.A2(n_15863),
.B(n_15820),
.Y(n_15944)
);

NAND3xp33_ASAP7_75t_L g15945 ( 
.A(n_15865),
.B(n_2683),
.C(n_2684),
.Y(n_15945)
);

OR2x2_ASAP7_75t_L g15946 ( 
.A(n_15821),
.B(n_2685),
.Y(n_15946)
);

INVx2_ASAP7_75t_L g15947 ( 
.A(n_15807),
.Y(n_15947)
);

OR2x2_ASAP7_75t_L g15948 ( 
.A(n_15879),
.B(n_2685),
.Y(n_15948)
);

NAND3xp33_ASAP7_75t_L g15949 ( 
.A(n_15897),
.B(n_2686),
.C(n_2688),
.Y(n_15949)
);

NOR3xp33_ASAP7_75t_SL g15950 ( 
.A(n_15896),
.B(n_2686),
.C(n_2688),
.Y(n_15950)
);

AOI22xp5_ASAP7_75t_L g15951 ( 
.A1(n_15887),
.A2(n_2691),
.B1(n_2689),
.B2(n_2690),
.Y(n_15951)
);

NAND3xp33_ASAP7_75t_L g15952 ( 
.A(n_15814),
.B(n_15835),
.C(n_15812),
.Y(n_15952)
);

NAND4xp75_ASAP7_75t_L g15953 ( 
.A(n_15829),
.B(n_2691),
.C(n_2689),
.D(n_2690),
.Y(n_15953)
);

AOI211x1_ASAP7_75t_L g15954 ( 
.A1(n_15900),
.A2(n_2694),
.B(n_2692),
.C(n_2693),
.Y(n_15954)
);

INVx1_ASAP7_75t_L g15955 ( 
.A(n_15841),
.Y(n_15955)
);

NAND3xp33_ASAP7_75t_L g15956 ( 
.A(n_15891),
.B(n_2692),
.C(n_2693),
.Y(n_15956)
);

INVx1_ASAP7_75t_L g15957 ( 
.A(n_15848),
.Y(n_15957)
);

NAND3xp33_ASAP7_75t_L g15958 ( 
.A(n_15803),
.B(n_2694),
.C(n_2695),
.Y(n_15958)
);

NOR3xp33_ASAP7_75t_L g15959 ( 
.A(n_15847),
.B(n_2695),
.C(n_2696),
.Y(n_15959)
);

AND2x2_ASAP7_75t_L g15960 ( 
.A(n_15804),
.B(n_2696),
.Y(n_15960)
);

AND2x2_ASAP7_75t_L g15961 ( 
.A(n_15831),
.B(n_15808),
.Y(n_15961)
);

NAND3xp33_ASAP7_75t_L g15962 ( 
.A(n_15806),
.B(n_2697),
.C(n_2698),
.Y(n_15962)
);

NOR2x1_ASAP7_75t_SL g15963 ( 
.A(n_15805),
.B(n_2697),
.Y(n_15963)
);

AND2x2_ASAP7_75t_L g15964 ( 
.A(n_15790),
.B(n_2698),
.Y(n_15964)
);

NAND3xp33_ASAP7_75t_L g15965 ( 
.A(n_15817),
.B(n_2699),
.C(n_2700),
.Y(n_15965)
);

OR2x2_ASAP7_75t_L g15966 ( 
.A(n_15837),
.B(n_2699),
.Y(n_15966)
);

NOR2xp33_ASAP7_75t_L g15967 ( 
.A(n_15836),
.B(n_2701),
.Y(n_15967)
);

AO21x2_ASAP7_75t_L g15968 ( 
.A1(n_15866),
.A2(n_2701),
.B(n_2702),
.Y(n_15968)
);

NAND4xp75_ASAP7_75t_L g15969 ( 
.A(n_15822),
.B(n_2704),
.C(n_2702),
.D(n_2703),
.Y(n_15969)
);

AOI22xp5_ASAP7_75t_L g15970 ( 
.A1(n_15830),
.A2(n_2705),
.B1(n_2703),
.B2(n_2704),
.Y(n_15970)
);

NOR2xp33_ASAP7_75t_L g15971 ( 
.A(n_15838),
.B(n_2705),
.Y(n_15971)
);

INVx1_ASAP7_75t_L g15972 ( 
.A(n_15861),
.Y(n_15972)
);

NOR2xp33_ASAP7_75t_L g15973 ( 
.A(n_15839),
.B(n_2706),
.Y(n_15973)
);

INVx1_ASAP7_75t_L g15974 ( 
.A(n_15834),
.Y(n_15974)
);

NOR2xp33_ASAP7_75t_L g15975 ( 
.A(n_15882),
.B(n_2706),
.Y(n_15975)
);

INVx1_ASAP7_75t_L g15976 ( 
.A(n_15842),
.Y(n_15976)
);

INVx2_ASAP7_75t_L g15977 ( 
.A(n_15795),
.Y(n_15977)
);

AOI22xp33_ASAP7_75t_L g15978 ( 
.A1(n_15892),
.A2(n_2709),
.B1(n_2707),
.B2(n_2708),
.Y(n_15978)
);

NOR2xp33_ASAP7_75t_L g15979 ( 
.A(n_15844),
.B(n_2707),
.Y(n_15979)
);

NAND2xp33_ASAP7_75t_SL g15980 ( 
.A(n_15870),
.B(n_2708),
.Y(n_15980)
);

NAND4xp75_ASAP7_75t_L g15981 ( 
.A(n_15860),
.B(n_2711),
.C(n_2709),
.D(n_2710),
.Y(n_15981)
);

AND2x2_ASAP7_75t_L g15982 ( 
.A(n_15894),
.B(n_2710),
.Y(n_15982)
);

NOR3xp33_ASAP7_75t_L g15983 ( 
.A(n_15855),
.B(n_2711),
.C(n_2712),
.Y(n_15983)
);

NOR3xp33_ASAP7_75t_L g15984 ( 
.A(n_15787),
.B(n_2712),
.C(n_2713),
.Y(n_15984)
);

INVx1_ASAP7_75t_L g15985 ( 
.A(n_15791),
.Y(n_15985)
);

INVxp67_ASAP7_75t_SL g15986 ( 
.A(n_15888),
.Y(n_15986)
);

AOI221xp5_ASAP7_75t_L g15987 ( 
.A1(n_15895),
.A2(n_2715),
.B1(n_2713),
.B2(n_2714),
.C(n_2716),
.Y(n_15987)
);

NAND3xp33_ASAP7_75t_SL g15988 ( 
.A(n_15871),
.B(n_2715),
.C(n_2716),
.Y(n_15988)
);

OR2x2_ASAP7_75t_L g15989 ( 
.A(n_15869),
.B(n_2717),
.Y(n_15989)
);

OAI221xp5_ASAP7_75t_SL g15990 ( 
.A1(n_15818),
.A2(n_2719),
.B1(n_2717),
.B2(n_2718),
.C(n_2720),
.Y(n_15990)
);

HB1xp67_ASAP7_75t_L g15991 ( 
.A(n_15833),
.Y(n_15991)
);

INVx3_ASAP7_75t_L g15992 ( 
.A(n_15854),
.Y(n_15992)
);

NAND2xp5_ASAP7_75t_L g15993 ( 
.A(n_15845),
.B(n_2720),
.Y(n_15993)
);

NAND4xp75_ASAP7_75t_L g15994 ( 
.A(n_15857),
.B(n_2723),
.C(n_2721),
.D(n_2722),
.Y(n_15994)
);

AOI22xp33_ASAP7_75t_SL g15995 ( 
.A1(n_15883),
.A2(n_2723),
.B1(n_2721),
.B2(n_2722),
.Y(n_15995)
);

INVx1_ASAP7_75t_L g15996 ( 
.A(n_15853),
.Y(n_15996)
);

AND2x2_ASAP7_75t_L g15997 ( 
.A(n_15851),
.B(n_2724),
.Y(n_15997)
);

NAND2xp5_ASAP7_75t_L g15998 ( 
.A(n_15899),
.B(n_2724),
.Y(n_15998)
);

NAND2xp5_ASAP7_75t_L g15999 ( 
.A(n_15843),
.B(n_2725),
.Y(n_15999)
);

NAND2xp5_ASAP7_75t_SL g16000 ( 
.A(n_15889),
.B(n_2726),
.Y(n_16000)
);

INVx1_ASAP7_75t_L g16001 ( 
.A(n_15850),
.Y(n_16001)
);

NOR3xp33_ASAP7_75t_L g16002 ( 
.A(n_15809),
.B(n_2727),
.C(n_2728),
.Y(n_16002)
);

NAND3xp33_ASAP7_75t_L g16003 ( 
.A(n_15849),
.B(n_2727),
.C(n_2729),
.Y(n_16003)
);

OR2x2_ASAP7_75t_L g16004 ( 
.A(n_15852),
.B(n_2729),
.Y(n_16004)
);

HB1xp67_ASAP7_75t_L g16005 ( 
.A(n_15810),
.Y(n_16005)
);

NAND3xp33_ASAP7_75t_L g16006 ( 
.A(n_15872),
.B(n_2730),
.C(n_2731),
.Y(n_16006)
);

AND2x2_ASAP7_75t_L g16007 ( 
.A(n_15873),
.B(n_2730),
.Y(n_16007)
);

INVx1_ASAP7_75t_L g16008 ( 
.A(n_15868),
.Y(n_16008)
);

INVx2_ASAP7_75t_L g16009 ( 
.A(n_15881),
.Y(n_16009)
);

AND2x2_ASAP7_75t_L g16010 ( 
.A(n_15885),
.B(n_2731),
.Y(n_16010)
);

OR2x2_ASAP7_75t_L g16011 ( 
.A(n_15801),
.B(n_2732),
.Y(n_16011)
);

AND2x2_ASAP7_75t_L g16012 ( 
.A(n_15785),
.B(n_2732),
.Y(n_16012)
);

AOI22xp33_ASAP7_75t_L g16013 ( 
.A1(n_15876),
.A2(n_2735),
.B1(n_2733),
.B2(n_2734),
.Y(n_16013)
);

NOR3xp33_ASAP7_75t_L g16014 ( 
.A(n_15876),
.B(n_2733),
.C(n_2734),
.Y(n_16014)
);

INVx1_ASAP7_75t_L g16015 ( 
.A(n_15789),
.Y(n_16015)
);

INVx2_ASAP7_75t_SL g16016 ( 
.A(n_15819),
.Y(n_16016)
);

OR2x2_ASAP7_75t_L g16017 ( 
.A(n_15801),
.B(n_2735),
.Y(n_16017)
);

NAND3xp33_ASAP7_75t_L g16018 ( 
.A(n_15877),
.B(n_2736),
.C(n_2737),
.Y(n_16018)
);

INVx2_ASAP7_75t_L g16019 ( 
.A(n_15819),
.Y(n_16019)
);

AOI221xp5_ASAP7_75t_L g16020 ( 
.A1(n_15886),
.A2(n_2739),
.B1(n_2737),
.B2(n_2738),
.C(n_2740),
.Y(n_16020)
);

NAND2xp5_ASAP7_75t_L g16021 ( 
.A(n_15825),
.B(n_2739),
.Y(n_16021)
);

AOI211xp5_ASAP7_75t_L g16022 ( 
.A1(n_15886),
.A2(n_2743),
.B(n_2741),
.C(n_2742),
.Y(n_16022)
);

BUFx3_ASAP7_75t_L g16023 ( 
.A(n_15800),
.Y(n_16023)
);

NAND2xp5_ASAP7_75t_L g16024 ( 
.A(n_15825),
.B(n_2742),
.Y(n_16024)
);

NAND3xp33_ASAP7_75t_L g16025 ( 
.A(n_15877),
.B(n_2743),
.C(n_2744),
.Y(n_16025)
);

AND2x2_ASAP7_75t_L g16026 ( 
.A(n_15785),
.B(n_2744),
.Y(n_16026)
);

INVx2_ASAP7_75t_L g16027 ( 
.A(n_15963),
.Y(n_16027)
);

INVx1_ASAP7_75t_L g16028 ( 
.A(n_15919),
.Y(n_16028)
);

AND2x4_ASAP7_75t_L g16029 ( 
.A(n_16023),
.B(n_2745),
.Y(n_16029)
);

INVx2_ASAP7_75t_L g16030 ( 
.A(n_16016),
.Y(n_16030)
);

INVx1_ASAP7_75t_L g16031 ( 
.A(n_15919),
.Y(n_16031)
);

INVxp33_ASAP7_75t_L g16032 ( 
.A(n_15910),
.Y(n_16032)
);

INVx1_ASAP7_75t_L g16033 ( 
.A(n_16012),
.Y(n_16033)
);

INVx1_ASAP7_75t_L g16034 ( 
.A(n_16026),
.Y(n_16034)
);

NAND2xp5_ASAP7_75t_L g16035 ( 
.A(n_15916),
.B(n_2745),
.Y(n_16035)
);

HB1xp67_ASAP7_75t_L g16036 ( 
.A(n_15968),
.Y(n_16036)
);

AND2x2_ASAP7_75t_L g16037 ( 
.A(n_15905),
.B(n_2746),
.Y(n_16037)
);

AND2x2_ASAP7_75t_L g16038 ( 
.A(n_15928),
.B(n_15961),
.Y(n_16038)
);

NAND2xp5_ASAP7_75t_L g16039 ( 
.A(n_16019),
.B(n_2747),
.Y(n_16039)
);

NAND4xp25_ASAP7_75t_L g16040 ( 
.A(n_15901),
.B(n_2749),
.C(n_2747),
.D(n_2748),
.Y(n_16040)
);

NAND2xp5_ASAP7_75t_SL g16041 ( 
.A(n_16018),
.B(n_2748),
.Y(n_16041)
);

INVx1_ASAP7_75t_L g16042 ( 
.A(n_16011),
.Y(n_16042)
);

OR2x2_ASAP7_75t_L g16043 ( 
.A(n_15944),
.B(n_2749),
.Y(n_16043)
);

NAND2xp5_ASAP7_75t_L g16044 ( 
.A(n_15903),
.B(n_2750),
.Y(n_16044)
);

NAND2x1_ASAP7_75t_L g16045 ( 
.A(n_16015),
.B(n_2750),
.Y(n_16045)
);

AND2x2_ASAP7_75t_L g16046 ( 
.A(n_15913),
.B(n_2751),
.Y(n_16046)
);

AND2x2_ASAP7_75t_L g16047 ( 
.A(n_15912),
.B(n_2752),
.Y(n_16047)
);

OR2x2_ASAP7_75t_L g16048 ( 
.A(n_16017),
.B(n_2752),
.Y(n_16048)
);

AND2x2_ASAP7_75t_L g16049 ( 
.A(n_15911),
.B(n_2753),
.Y(n_16049)
);

INVx2_ASAP7_75t_L g16050 ( 
.A(n_15946),
.Y(n_16050)
);

AND2x2_ASAP7_75t_L g16051 ( 
.A(n_15942),
.B(n_2753),
.Y(n_16051)
);

INVx1_ASAP7_75t_L g16052 ( 
.A(n_15917),
.Y(n_16052)
);

INVx1_ASAP7_75t_L g16053 ( 
.A(n_15921),
.Y(n_16053)
);

OR2x2_ASAP7_75t_L g16054 ( 
.A(n_15947),
.B(n_2754),
.Y(n_16054)
);

NAND2xp5_ASAP7_75t_L g16055 ( 
.A(n_15907),
.B(n_2754),
.Y(n_16055)
);

NOR2xp33_ASAP7_75t_SL g16056 ( 
.A(n_15920),
.B(n_15953),
.Y(n_16056)
);

AND2x2_ASAP7_75t_L g16057 ( 
.A(n_15941),
.B(n_2755),
.Y(n_16057)
);

INVx1_ASAP7_75t_L g16058 ( 
.A(n_15925),
.Y(n_16058)
);

OR2x2_ASAP7_75t_L g16059 ( 
.A(n_15989),
.B(n_15948),
.Y(n_16059)
);

INVx1_ASAP7_75t_L g16060 ( 
.A(n_15927),
.Y(n_16060)
);

INVx2_ASAP7_75t_L g16061 ( 
.A(n_15940),
.Y(n_16061)
);

INVx1_ASAP7_75t_L g16062 ( 
.A(n_15991),
.Y(n_16062)
);

NAND2xp5_ASAP7_75t_L g16063 ( 
.A(n_15904),
.B(n_2756),
.Y(n_16063)
);

AND2x2_ASAP7_75t_L g16064 ( 
.A(n_15950),
.B(n_2756),
.Y(n_16064)
);

NAND2xp5_ASAP7_75t_L g16065 ( 
.A(n_15923),
.B(n_2757),
.Y(n_16065)
);

INVx1_ASAP7_75t_L g16066 ( 
.A(n_15964),
.Y(n_16066)
);

HB1xp67_ASAP7_75t_L g16067 ( 
.A(n_15969),
.Y(n_16067)
);

INVx2_ASAP7_75t_L g16068 ( 
.A(n_15966),
.Y(n_16068)
);

AND2x2_ASAP7_75t_L g16069 ( 
.A(n_15982),
.B(n_2758),
.Y(n_16069)
);

INVx2_ASAP7_75t_L g16070 ( 
.A(n_15931),
.Y(n_16070)
);

AND2x2_ASAP7_75t_L g16071 ( 
.A(n_15955),
.B(n_2758),
.Y(n_16071)
);

BUFx2_ASAP7_75t_L g16072 ( 
.A(n_15980),
.Y(n_16072)
);

AND2x4_ASAP7_75t_L g16073 ( 
.A(n_15957),
.B(n_2760),
.Y(n_16073)
);

INVx1_ASAP7_75t_L g16074 ( 
.A(n_16021),
.Y(n_16074)
);

INVx2_ASAP7_75t_L g16075 ( 
.A(n_16004),
.Y(n_16075)
);

AND2x2_ASAP7_75t_L g16076 ( 
.A(n_15914),
.B(n_15909),
.Y(n_16076)
);

INVxp67_ASAP7_75t_SL g16077 ( 
.A(n_15943),
.Y(n_16077)
);

HB1xp67_ASAP7_75t_L g16078 ( 
.A(n_15994),
.Y(n_16078)
);

AND2x2_ASAP7_75t_L g16079 ( 
.A(n_15972),
.B(n_2760),
.Y(n_16079)
);

BUFx2_ASAP7_75t_L g16080 ( 
.A(n_15977),
.Y(n_16080)
);

NAND2xp5_ASAP7_75t_L g16081 ( 
.A(n_15995),
.B(n_2761),
.Y(n_16081)
);

AND2x4_ASAP7_75t_SL g16082 ( 
.A(n_15992),
.B(n_2761),
.Y(n_16082)
);

INVx1_ASAP7_75t_L g16083 ( 
.A(n_16024),
.Y(n_16083)
);

AND2x2_ASAP7_75t_L g16084 ( 
.A(n_15908),
.B(n_15915),
.Y(n_16084)
);

OR2x2_ASAP7_75t_L g16085 ( 
.A(n_16025),
.B(n_2762),
.Y(n_16085)
);

AND2x4_ASAP7_75t_L g16086 ( 
.A(n_15960),
.B(n_2762),
.Y(n_16086)
);

AND2x2_ASAP7_75t_L g16087 ( 
.A(n_15938),
.B(n_2763),
.Y(n_16087)
);

AOI22xp33_ASAP7_75t_L g16088 ( 
.A1(n_15902),
.A2(n_2765),
.B1(n_2763),
.B2(n_2764),
.Y(n_16088)
);

HB1xp67_ASAP7_75t_L g16089 ( 
.A(n_15981),
.Y(n_16089)
);

NAND2xp5_ASAP7_75t_L g16090 ( 
.A(n_15939),
.B(n_2764),
.Y(n_16090)
);

AND2x2_ASAP7_75t_L g16091 ( 
.A(n_15974),
.B(n_2765),
.Y(n_16091)
);

AND2x2_ASAP7_75t_L g16092 ( 
.A(n_15976),
.B(n_2766),
.Y(n_16092)
);

INVx1_ASAP7_75t_L g16093 ( 
.A(n_15930),
.Y(n_16093)
);

NAND2xp5_ASAP7_75t_L g16094 ( 
.A(n_15984),
.B(n_2766),
.Y(n_16094)
);

INVx1_ASAP7_75t_L g16095 ( 
.A(n_15934),
.Y(n_16095)
);

AND2x4_ASAP7_75t_L g16096 ( 
.A(n_16009),
.B(n_2767),
.Y(n_16096)
);

NAND2xp67_ASAP7_75t_L g16097 ( 
.A(n_15997),
.B(n_2768),
.Y(n_16097)
);

OR2x2_ASAP7_75t_L g16098 ( 
.A(n_15988),
.B(n_15922),
.Y(n_16098)
);

INVx2_ASAP7_75t_L g16099 ( 
.A(n_16007),
.Y(n_16099)
);

AND2x2_ASAP7_75t_L g16100 ( 
.A(n_15986),
.B(n_2768),
.Y(n_16100)
);

OR2x6_ASAP7_75t_L g16101 ( 
.A(n_16005),
.B(n_2769),
.Y(n_16101)
);

INVx1_ASAP7_75t_L g16102 ( 
.A(n_15952),
.Y(n_16102)
);

INVx1_ASAP7_75t_L g16103 ( 
.A(n_16010),
.Y(n_16103)
);

NAND2xp5_ASAP7_75t_L g16104 ( 
.A(n_15954),
.B(n_2769),
.Y(n_16104)
);

INVx1_ASAP7_75t_L g16105 ( 
.A(n_15932),
.Y(n_16105)
);

NOR2x1_ASAP7_75t_L g16106 ( 
.A(n_15958),
.B(n_15962),
.Y(n_16106)
);

INVxp67_ASAP7_75t_L g16107 ( 
.A(n_15967),
.Y(n_16107)
);

AND2x4_ASAP7_75t_L g16108 ( 
.A(n_15996),
.B(n_2770),
.Y(n_16108)
);

INVx2_ASAP7_75t_L g16109 ( 
.A(n_15985),
.Y(n_16109)
);

INVx1_ASAP7_75t_L g16110 ( 
.A(n_15935),
.Y(n_16110)
);

OR2x2_ASAP7_75t_L g16111 ( 
.A(n_15906),
.B(n_2770),
.Y(n_16111)
);

INVx2_ASAP7_75t_L g16112 ( 
.A(n_15999),
.Y(n_16112)
);

INVx1_ASAP7_75t_L g16113 ( 
.A(n_15971),
.Y(n_16113)
);

NOR2xp33_ASAP7_75t_SL g16114 ( 
.A(n_15990),
.B(n_15924),
.Y(n_16114)
);

OR2x2_ASAP7_75t_L g16115 ( 
.A(n_15993),
.B(n_2771),
.Y(n_16115)
);

AND2x2_ASAP7_75t_L g16116 ( 
.A(n_15918),
.B(n_16014),
.Y(n_16116)
);

INVx1_ASAP7_75t_L g16117 ( 
.A(n_15973),
.Y(n_16117)
);

INVx1_ASAP7_75t_L g16118 ( 
.A(n_15979),
.Y(n_16118)
);

NOR2x1_ASAP7_75t_L g16119 ( 
.A(n_15965),
.B(n_2771),
.Y(n_16119)
);

AND2x2_ASAP7_75t_L g16120 ( 
.A(n_15975),
.B(n_2772),
.Y(n_16120)
);

AND2x2_ASAP7_75t_L g16121 ( 
.A(n_16022),
.B(n_2772),
.Y(n_16121)
);

AND2x2_ASAP7_75t_L g16122 ( 
.A(n_16001),
.B(n_2773),
.Y(n_16122)
);

INVx1_ASAP7_75t_L g16123 ( 
.A(n_15945),
.Y(n_16123)
);

INVxp67_ASAP7_75t_L g16124 ( 
.A(n_15998),
.Y(n_16124)
);

NAND2xp5_ASAP7_75t_L g16125 ( 
.A(n_16013),
.B(n_2773),
.Y(n_16125)
);

INVx2_ASAP7_75t_SL g16126 ( 
.A(n_16008),
.Y(n_16126)
);

OR2x2_ASAP7_75t_L g16127 ( 
.A(n_15956),
.B(n_2774),
.Y(n_16127)
);

HB1xp67_ASAP7_75t_L g16128 ( 
.A(n_16003),
.Y(n_16128)
);

INVx1_ASAP7_75t_L g16129 ( 
.A(n_16006),
.Y(n_16129)
);

NAND2xp5_ASAP7_75t_L g16130 ( 
.A(n_15929),
.B(n_2774),
.Y(n_16130)
);

INVx1_ASAP7_75t_L g16131 ( 
.A(n_15949),
.Y(n_16131)
);

INVx3_ASAP7_75t_SL g16132 ( 
.A(n_16000),
.Y(n_16132)
);

NAND2xp5_ASAP7_75t_SL g16133 ( 
.A(n_15933),
.B(n_16020),
.Y(n_16133)
);

AND2x2_ASAP7_75t_L g16134 ( 
.A(n_15959),
.B(n_2775),
.Y(n_16134)
);

AND2x2_ASAP7_75t_L g16135 ( 
.A(n_16002),
.B(n_2775),
.Y(n_16135)
);

OR2x2_ASAP7_75t_L g16136 ( 
.A(n_15926),
.B(n_2776),
.Y(n_16136)
);

INVx1_ASAP7_75t_L g16137 ( 
.A(n_15970),
.Y(n_16137)
);

INVx1_ASAP7_75t_L g16138 ( 
.A(n_15951),
.Y(n_16138)
);

AND2x4_ASAP7_75t_L g16139 ( 
.A(n_15983),
.B(n_2777),
.Y(n_16139)
);

NAND2xp5_ASAP7_75t_L g16140 ( 
.A(n_15978),
.B(n_15937),
.Y(n_16140)
);

AND2x2_ASAP7_75t_L g16141 ( 
.A(n_15987),
.B(n_2778),
.Y(n_16141)
);

INVx1_ASAP7_75t_L g16142 ( 
.A(n_15936),
.Y(n_16142)
);

AND2x2_ASAP7_75t_L g16143 ( 
.A(n_16023),
.B(n_2779),
.Y(n_16143)
);

AND2x2_ASAP7_75t_L g16144 ( 
.A(n_16023),
.B(n_2779),
.Y(n_16144)
);

AND2x4_ASAP7_75t_L g16145 ( 
.A(n_16023),
.B(n_2780),
.Y(n_16145)
);

OR2x2_ASAP7_75t_L g16146 ( 
.A(n_16016),
.B(n_2780),
.Y(n_16146)
);

INVx2_ASAP7_75t_L g16147 ( 
.A(n_15963),
.Y(n_16147)
);

NAND2xp5_ASAP7_75t_L g16148 ( 
.A(n_16016),
.B(n_2781),
.Y(n_16148)
);

INVx2_ASAP7_75t_L g16149 ( 
.A(n_15963),
.Y(n_16149)
);

BUFx3_ASAP7_75t_L g16150 ( 
.A(n_16023),
.Y(n_16150)
);

INVx1_ASAP7_75t_L g16151 ( 
.A(n_15963),
.Y(n_16151)
);

INVx2_ASAP7_75t_SL g16152 ( 
.A(n_16016),
.Y(n_16152)
);

NAND2xp5_ASAP7_75t_L g16153 ( 
.A(n_16016),
.B(n_2781),
.Y(n_16153)
);

INVx2_ASAP7_75t_L g16154 ( 
.A(n_15963),
.Y(n_16154)
);

NOR2x1_ASAP7_75t_L g16155 ( 
.A(n_15920),
.B(n_2782),
.Y(n_16155)
);

AND2x2_ASAP7_75t_L g16156 ( 
.A(n_16023),
.B(n_2782),
.Y(n_16156)
);

OR2x2_ASAP7_75t_L g16157 ( 
.A(n_16016),
.B(n_2783),
.Y(n_16157)
);

INVx3_ASAP7_75t_L g16158 ( 
.A(n_16023),
.Y(n_16158)
);

NAND2xp5_ASAP7_75t_L g16159 ( 
.A(n_16016),
.B(n_2783),
.Y(n_16159)
);

AND2x4_ASAP7_75t_L g16160 ( 
.A(n_16023),
.B(n_2784),
.Y(n_16160)
);

NAND2xp5_ASAP7_75t_L g16161 ( 
.A(n_16016),
.B(n_2785),
.Y(n_16161)
);

AND2x4_ASAP7_75t_L g16162 ( 
.A(n_16023),
.B(n_2785),
.Y(n_16162)
);

AND2x2_ASAP7_75t_L g16163 ( 
.A(n_16023),
.B(n_2786),
.Y(n_16163)
);

OR2x2_ASAP7_75t_L g16164 ( 
.A(n_16016),
.B(n_2786),
.Y(n_16164)
);

NAND2xp5_ASAP7_75t_L g16165 ( 
.A(n_16016),
.B(n_2787),
.Y(n_16165)
);

OR2x2_ASAP7_75t_L g16166 ( 
.A(n_16016),
.B(n_2788),
.Y(n_16166)
);

INVx1_ASAP7_75t_L g16167 ( 
.A(n_15963),
.Y(n_16167)
);

NAND3xp33_ASAP7_75t_L g16168 ( 
.A(n_15984),
.B(n_2788),
.C(n_2789),
.Y(n_16168)
);

AND2x2_ASAP7_75t_L g16169 ( 
.A(n_16023),
.B(n_2789),
.Y(n_16169)
);

NOR2xp33_ASAP7_75t_L g16170 ( 
.A(n_16016),
.B(n_2791),
.Y(n_16170)
);

NAND2xp5_ASAP7_75t_L g16171 ( 
.A(n_16016),
.B(n_2791),
.Y(n_16171)
);

INVxp67_ASAP7_75t_L g16172 ( 
.A(n_15963),
.Y(n_16172)
);

INVx1_ASAP7_75t_L g16173 ( 
.A(n_15963),
.Y(n_16173)
);

AND2x2_ASAP7_75t_L g16174 ( 
.A(n_16023),
.B(n_2792),
.Y(n_16174)
);

AND2x2_ASAP7_75t_L g16175 ( 
.A(n_16023),
.B(n_2793),
.Y(n_16175)
);

AOI22xp33_ASAP7_75t_L g16176 ( 
.A1(n_16023),
.A2(n_2796),
.B1(n_2794),
.B2(n_2795),
.Y(n_16176)
);

INVx1_ASAP7_75t_L g16177 ( 
.A(n_15963),
.Y(n_16177)
);

AND2x4_ASAP7_75t_SL g16178 ( 
.A(n_16038),
.B(n_2794),
.Y(n_16178)
);

INVx2_ASAP7_75t_L g16179 ( 
.A(n_16150),
.Y(n_16179)
);

INVx1_ASAP7_75t_L g16180 ( 
.A(n_16036),
.Y(n_16180)
);

INVx3_ASAP7_75t_L g16181 ( 
.A(n_16027),
.Y(n_16181)
);

OR2x2_ASAP7_75t_L g16182 ( 
.A(n_16147),
.B(n_2795),
.Y(n_16182)
);

INVx2_ASAP7_75t_L g16183 ( 
.A(n_16149),
.Y(n_16183)
);

AOI22xp5_ASAP7_75t_L g16184 ( 
.A1(n_16056),
.A2(n_2798),
.B1(n_2796),
.B2(n_2797),
.Y(n_16184)
);

AND2x4_ASAP7_75t_L g16185 ( 
.A(n_16154),
.B(n_2797),
.Y(n_16185)
);

NAND2xp5_ASAP7_75t_L g16186 ( 
.A(n_16028),
.B(n_2798),
.Y(n_16186)
);

INVx1_ASAP7_75t_L g16187 ( 
.A(n_16151),
.Y(n_16187)
);

INVx1_ASAP7_75t_L g16188 ( 
.A(n_16167),
.Y(n_16188)
);

INVx2_ASAP7_75t_SL g16189 ( 
.A(n_16082),
.Y(n_16189)
);

HB1xp67_ASAP7_75t_L g16190 ( 
.A(n_16177),
.Y(n_16190)
);

AND2x2_ASAP7_75t_L g16191 ( 
.A(n_16046),
.B(n_2799),
.Y(n_16191)
);

AOI22xp33_ASAP7_75t_L g16192 ( 
.A1(n_16102),
.A2(n_2801),
.B1(n_2799),
.B2(n_2800),
.Y(n_16192)
);

AOI211x1_ASAP7_75t_SL g16193 ( 
.A1(n_16063),
.A2(n_2803),
.B(n_2800),
.C(n_2802),
.Y(n_16193)
);

NAND3xp33_ASAP7_75t_L g16194 ( 
.A(n_16172),
.B(n_2802),
.C(n_2803),
.Y(n_16194)
);

INVx1_ASAP7_75t_L g16195 ( 
.A(n_16173),
.Y(n_16195)
);

INVx1_ASAP7_75t_L g16196 ( 
.A(n_16051),
.Y(n_16196)
);

AOI22xp33_ASAP7_75t_L g16197 ( 
.A1(n_16032),
.A2(n_2806),
.B1(n_2804),
.B2(n_2805),
.Y(n_16197)
);

INVx1_ASAP7_75t_L g16198 ( 
.A(n_16031),
.Y(n_16198)
);

NAND2xp5_ASAP7_75t_L g16199 ( 
.A(n_16152),
.B(n_2804),
.Y(n_16199)
);

INVx1_ASAP7_75t_L g16200 ( 
.A(n_16045),
.Y(n_16200)
);

AOI22xp33_ASAP7_75t_L g16201 ( 
.A1(n_16158),
.A2(n_2808),
.B1(n_2805),
.B2(n_2807),
.Y(n_16201)
);

OR2x2_ASAP7_75t_L g16202 ( 
.A(n_16059),
.B(n_2807),
.Y(n_16202)
);

INVx1_ASAP7_75t_L g16203 ( 
.A(n_16097),
.Y(n_16203)
);

HB1xp67_ASAP7_75t_L g16204 ( 
.A(n_16101),
.Y(n_16204)
);

INVx1_ASAP7_75t_L g16205 ( 
.A(n_16072),
.Y(n_16205)
);

INVx3_ASAP7_75t_L g16206 ( 
.A(n_16029),
.Y(n_16206)
);

INVx3_ASAP7_75t_L g16207 ( 
.A(n_16145),
.Y(n_16207)
);

AOI22xp5_ASAP7_75t_L g16208 ( 
.A1(n_16114),
.A2(n_16030),
.B1(n_16142),
.B2(n_16084),
.Y(n_16208)
);

INVx1_ASAP7_75t_L g16209 ( 
.A(n_16043),
.Y(n_16209)
);

OA21x2_ASAP7_75t_L g16210 ( 
.A1(n_16062),
.A2(n_2808),
.B(n_2809),
.Y(n_16210)
);

INVx1_ASAP7_75t_SL g16211 ( 
.A(n_16047),
.Y(n_16211)
);

INVxp67_ASAP7_75t_L g16212 ( 
.A(n_16170),
.Y(n_16212)
);

OR2x2_ASAP7_75t_L g16213 ( 
.A(n_16055),
.B(n_2810),
.Y(n_16213)
);

HB1xp67_ASAP7_75t_L g16214 ( 
.A(n_16101),
.Y(n_16214)
);

AND2x4_ASAP7_75t_SL g16215 ( 
.A(n_16076),
.B(n_2810),
.Y(n_16215)
);

OAI21xp5_ASAP7_75t_L g16216 ( 
.A1(n_16155),
.A2(n_2811),
.B(n_2812),
.Y(n_16216)
);

INVx1_ASAP7_75t_L g16217 ( 
.A(n_16146),
.Y(n_16217)
);

INVx1_ASAP7_75t_L g16218 ( 
.A(n_16157),
.Y(n_16218)
);

INVx2_ASAP7_75t_L g16219 ( 
.A(n_16164),
.Y(n_16219)
);

HB1xp67_ASAP7_75t_L g16220 ( 
.A(n_16166),
.Y(n_16220)
);

AND2x2_ASAP7_75t_L g16221 ( 
.A(n_16049),
.B(n_2811),
.Y(n_16221)
);

INVx2_ASAP7_75t_L g16222 ( 
.A(n_16160),
.Y(n_16222)
);

AND2x2_ASAP7_75t_L g16223 ( 
.A(n_16037),
.B(n_2813),
.Y(n_16223)
);

INVx1_ASAP7_75t_L g16224 ( 
.A(n_16143),
.Y(n_16224)
);

INVx1_ASAP7_75t_L g16225 ( 
.A(n_16144),
.Y(n_16225)
);

INVx2_ASAP7_75t_L g16226 ( 
.A(n_16162),
.Y(n_16226)
);

INVx2_ASAP7_75t_SL g16227 ( 
.A(n_16108),
.Y(n_16227)
);

NAND2x1p5_ASAP7_75t_L g16228 ( 
.A(n_16042),
.B(n_16156),
.Y(n_16228)
);

AND2x2_ASAP7_75t_L g16229 ( 
.A(n_16163),
.B(n_2813),
.Y(n_16229)
);

OAI21xp33_ASAP7_75t_L g16230 ( 
.A1(n_16140),
.A2(n_2814),
.B(n_2815),
.Y(n_16230)
);

INVx1_ASAP7_75t_L g16231 ( 
.A(n_16169),
.Y(n_16231)
);

INVx1_ASAP7_75t_L g16232 ( 
.A(n_16174),
.Y(n_16232)
);

AND3x2_ASAP7_75t_L g16233 ( 
.A(n_16080),
.B(n_2814),
.C(n_2815),
.Y(n_16233)
);

INVx2_ASAP7_75t_L g16234 ( 
.A(n_16048),
.Y(n_16234)
);

INVx1_ASAP7_75t_L g16235 ( 
.A(n_16175),
.Y(n_16235)
);

NAND4xp75_ASAP7_75t_L g16236 ( 
.A(n_16119),
.B(n_2818),
.C(n_2816),
.D(n_2817),
.Y(n_16236)
);

INVxp67_ASAP7_75t_L g16237 ( 
.A(n_16067),
.Y(n_16237)
);

AOI22xp5_ASAP7_75t_L g16238 ( 
.A1(n_16033),
.A2(n_16034),
.B1(n_16133),
.B2(n_16089),
.Y(n_16238)
);

INVx1_ASAP7_75t_L g16239 ( 
.A(n_16069),
.Y(n_16239)
);

INVx2_ASAP7_75t_L g16240 ( 
.A(n_16086),
.Y(n_16240)
);

NOR2xp33_ASAP7_75t_R g16241 ( 
.A(n_16052),
.B(n_2816),
.Y(n_16241)
);

INVx1_ASAP7_75t_L g16242 ( 
.A(n_16100),
.Y(n_16242)
);

INVx3_ASAP7_75t_L g16243 ( 
.A(n_16073),
.Y(n_16243)
);

NAND2xp5_ASAP7_75t_L g16244 ( 
.A(n_16087),
.B(n_2817),
.Y(n_16244)
);

AND2x2_ASAP7_75t_L g16245 ( 
.A(n_16064),
.B(n_2818),
.Y(n_16245)
);

INVx1_ASAP7_75t_L g16246 ( 
.A(n_16071),
.Y(n_16246)
);

OR2x2_ASAP7_75t_L g16247 ( 
.A(n_16136),
.B(n_2819),
.Y(n_16247)
);

INVx2_ASAP7_75t_L g16248 ( 
.A(n_16054),
.Y(n_16248)
);

INVx1_ASAP7_75t_L g16249 ( 
.A(n_16079),
.Y(n_16249)
);

INVx3_ASAP7_75t_L g16250 ( 
.A(n_16096),
.Y(n_16250)
);

AOI22xp5_ASAP7_75t_L g16251 ( 
.A1(n_16078),
.A2(n_2822),
.B1(n_2820),
.B2(n_2821),
.Y(n_16251)
);

HB1xp67_ASAP7_75t_L g16252 ( 
.A(n_16091),
.Y(n_16252)
);

INVx1_ASAP7_75t_L g16253 ( 
.A(n_16148),
.Y(n_16253)
);

INVx1_ASAP7_75t_SL g16254 ( 
.A(n_16132),
.Y(n_16254)
);

INVx1_ASAP7_75t_SL g16255 ( 
.A(n_16085),
.Y(n_16255)
);

BUFx2_ASAP7_75t_L g16256 ( 
.A(n_16092),
.Y(n_16256)
);

INVx2_ASAP7_75t_L g16257 ( 
.A(n_16057),
.Y(n_16257)
);

INVx4_ASAP7_75t_L g16258 ( 
.A(n_16061),
.Y(n_16258)
);

INVx2_ASAP7_75t_L g16259 ( 
.A(n_16120),
.Y(n_16259)
);

OAI21x1_ASAP7_75t_L g16260 ( 
.A1(n_16106),
.A2(n_16041),
.B(n_16153),
.Y(n_16260)
);

HB1xp67_ASAP7_75t_L g16261 ( 
.A(n_16050),
.Y(n_16261)
);

AND2x2_ASAP7_75t_L g16262 ( 
.A(n_16066),
.B(n_16121),
.Y(n_16262)
);

AND2x2_ASAP7_75t_L g16263 ( 
.A(n_16099),
.B(n_16116),
.Y(n_16263)
);

OAI21xp33_ASAP7_75t_L g16264 ( 
.A1(n_16137),
.A2(n_2821),
.B(n_2822),
.Y(n_16264)
);

OA21x2_ASAP7_75t_L g16265 ( 
.A1(n_16104),
.A2(n_2823),
.B(n_2824),
.Y(n_16265)
);

INVx2_ASAP7_75t_SL g16266 ( 
.A(n_16159),
.Y(n_16266)
);

INVx2_ASAP7_75t_L g16267 ( 
.A(n_16115),
.Y(n_16267)
);

INVx2_ASAP7_75t_L g16268 ( 
.A(n_16122),
.Y(n_16268)
);

INVx1_ASAP7_75t_L g16269 ( 
.A(n_16161),
.Y(n_16269)
);

INVx1_ASAP7_75t_L g16270 ( 
.A(n_16165),
.Y(n_16270)
);

INVx4_ASAP7_75t_L g16271 ( 
.A(n_16068),
.Y(n_16271)
);

INVx1_ASAP7_75t_SL g16272 ( 
.A(n_16098),
.Y(n_16272)
);

BUFx2_ASAP7_75t_L g16273 ( 
.A(n_16171),
.Y(n_16273)
);

OR2x2_ASAP7_75t_L g16274 ( 
.A(n_16040),
.B(n_2823),
.Y(n_16274)
);

INVx1_ASAP7_75t_SL g16275 ( 
.A(n_16111),
.Y(n_16275)
);

INVx3_ASAP7_75t_L g16276 ( 
.A(n_16075),
.Y(n_16276)
);

INVx3_ASAP7_75t_L g16277 ( 
.A(n_16109),
.Y(n_16277)
);

INVx1_ASAP7_75t_L g16278 ( 
.A(n_16090),
.Y(n_16278)
);

AND2x2_ASAP7_75t_L g16279 ( 
.A(n_16103),
.B(n_2824),
.Y(n_16279)
);

AO21x2_ASAP7_75t_L g16280 ( 
.A1(n_16044),
.A2(n_16039),
.B(n_16035),
.Y(n_16280)
);

NAND2xp5_ASAP7_75t_L g16281 ( 
.A(n_16139),
.B(n_2825),
.Y(n_16281)
);

AND2x2_ASAP7_75t_L g16282 ( 
.A(n_16128),
.B(n_2825),
.Y(n_16282)
);

AND3x1_ASAP7_75t_L g16283 ( 
.A(n_16134),
.B(n_2826),
.C(n_2827),
.Y(n_16283)
);

NAND2xp5_ASAP7_75t_SL g16284 ( 
.A(n_16126),
.B(n_2826),
.Y(n_16284)
);

AOI22xp5_ASAP7_75t_L g16285 ( 
.A1(n_16110),
.A2(n_2829),
.B1(n_2827),
.B2(n_2828),
.Y(n_16285)
);

HB1xp67_ASAP7_75t_L g16286 ( 
.A(n_16127),
.Y(n_16286)
);

INVx1_ASAP7_75t_L g16287 ( 
.A(n_16065),
.Y(n_16287)
);

AOI22xp33_ASAP7_75t_L g16288 ( 
.A1(n_16129),
.A2(n_2830),
.B1(n_2828),
.B2(n_2829),
.Y(n_16288)
);

AND2x4_ASAP7_75t_L g16289 ( 
.A(n_16070),
.B(n_16105),
.Y(n_16289)
);

NOR2xp33_ASAP7_75t_L g16290 ( 
.A(n_16168),
.B(n_2831),
.Y(n_16290)
);

AOI21xp5_ASAP7_75t_L g16291 ( 
.A1(n_16094),
.A2(n_2832),
.B(n_2833),
.Y(n_16291)
);

OR2x6_ASAP7_75t_L g16292 ( 
.A(n_16113),
.B(n_2832),
.Y(n_16292)
);

OA21x2_ASAP7_75t_L g16293 ( 
.A1(n_16081),
.A2(n_2833),
.B(n_2834),
.Y(n_16293)
);

INVx1_ASAP7_75t_L g16294 ( 
.A(n_16130),
.Y(n_16294)
);

INVx2_ASAP7_75t_L g16295 ( 
.A(n_16053),
.Y(n_16295)
);

OR2x2_ASAP7_75t_L g16296 ( 
.A(n_16058),
.B(n_16060),
.Y(n_16296)
);

HB1xp67_ASAP7_75t_L g16297 ( 
.A(n_16135),
.Y(n_16297)
);

INVx1_ASAP7_75t_L g16298 ( 
.A(n_16123),
.Y(n_16298)
);

NAND2xp5_ASAP7_75t_L g16299 ( 
.A(n_16088),
.B(n_2834),
.Y(n_16299)
);

OR2x2_ASAP7_75t_L g16300 ( 
.A(n_16131),
.B(n_2835),
.Y(n_16300)
);

INVx4_ASAP7_75t_L g16301 ( 
.A(n_16112),
.Y(n_16301)
);

INVx1_ASAP7_75t_L g16302 ( 
.A(n_16125),
.Y(n_16302)
);

BUFx2_ASAP7_75t_L g16303 ( 
.A(n_16077),
.Y(n_16303)
);

AO21x2_ASAP7_75t_L g16304 ( 
.A1(n_16117),
.A2(n_2836),
.B(n_2837),
.Y(n_16304)
);

BUFx2_ASAP7_75t_L g16305 ( 
.A(n_16138),
.Y(n_16305)
);

BUFx3_ASAP7_75t_L g16306 ( 
.A(n_16118),
.Y(n_16306)
);

INVx1_ASAP7_75t_L g16307 ( 
.A(n_16095),
.Y(n_16307)
);

INVx4_ASAP7_75t_L g16308 ( 
.A(n_16074),
.Y(n_16308)
);

HB1xp67_ASAP7_75t_L g16309 ( 
.A(n_16124),
.Y(n_16309)
);

AND2x2_ASAP7_75t_L g16310 ( 
.A(n_16141),
.B(n_2836),
.Y(n_16310)
);

NOR2xp33_ASAP7_75t_L g16311 ( 
.A(n_16107),
.B(n_2837),
.Y(n_16311)
);

NAND2xp5_ASAP7_75t_L g16312 ( 
.A(n_16083),
.B(n_2838),
.Y(n_16312)
);

INVx2_ASAP7_75t_L g16313 ( 
.A(n_16093),
.Y(n_16313)
);

INVx4_ASAP7_75t_L g16314 ( 
.A(n_16176),
.Y(n_16314)
);

INVx2_ASAP7_75t_L g16315 ( 
.A(n_16150),
.Y(n_16315)
);

AOI22xp33_ASAP7_75t_L g16316 ( 
.A1(n_16102),
.A2(n_2840),
.B1(n_2838),
.B2(n_2839),
.Y(n_16316)
);

INVx1_ASAP7_75t_L g16317 ( 
.A(n_16036),
.Y(n_16317)
);

INVx1_ASAP7_75t_L g16318 ( 
.A(n_16036),
.Y(n_16318)
);

INVx2_ASAP7_75t_L g16319 ( 
.A(n_16150),
.Y(n_16319)
);

AND2x2_ASAP7_75t_L g16320 ( 
.A(n_16038),
.B(n_2839),
.Y(n_16320)
);

INVx1_ASAP7_75t_L g16321 ( 
.A(n_16036),
.Y(n_16321)
);

NAND4xp25_ASAP7_75t_L g16322 ( 
.A(n_16114),
.B(n_2843),
.C(n_2841),
.D(n_2842),
.Y(n_16322)
);

NOR3xp33_ASAP7_75t_L g16323 ( 
.A(n_16258),
.B(n_2841),
.C(n_2842),
.Y(n_16323)
);

INVx1_ASAP7_75t_L g16324 ( 
.A(n_16190),
.Y(n_16324)
);

INVx1_ASAP7_75t_L g16325 ( 
.A(n_16304),
.Y(n_16325)
);

AND2x2_ASAP7_75t_L g16326 ( 
.A(n_16206),
.B(n_2843),
.Y(n_16326)
);

AND2x2_ASAP7_75t_L g16327 ( 
.A(n_16207),
.B(n_2844),
.Y(n_16327)
);

INVx1_ASAP7_75t_L g16328 ( 
.A(n_16204),
.Y(n_16328)
);

INVx1_ASAP7_75t_L g16329 ( 
.A(n_16214),
.Y(n_16329)
);

INVx2_ASAP7_75t_L g16330 ( 
.A(n_16233),
.Y(n_16330)
);

NOR2xp33_ASAP7_75t_L g16331 ( 
.A(n_16181),
.B(n_2844),
.Y(n_16331)
);

NOR2xp33_ASAP7_75t_L g16332 ( 
.A(n_16200),
.B(n_2845),
.Y(n_16332)
);

NAND2xp5_ASAP7_75t_SL g16333 ( 
.A(n_16185),
.B(n_16189),
.Y(n_16333)
);

INVx2_ASAP7_75t_L g16334 ( 
.A(n_16210),
.Y(n_16334)
);

OR2x2_ASAP7_75t_L g16335 ( 
.A(n_16202),
.B(n_2846),
.Y(n_16335)
);

NAND2xp5_ASAP7_75t_L g16336 ( 
.A(n_16320),
.B(n_2847),
.Y(n_16336)
);

AND2x2_ASAP7_75t_L g16337 ( 
.A(n_16179),
.B(n_2847),
.Y(n_16337)
);

NAND2xp5_ASAP7_75t_SL g16338 ( 
.A(n_16283),
.B(n_2848),
.Y(n_16338)
);

NOR2x1_ASAP7_75t_L g16339 ( 
.A(n_16236),
.B(n_16194),
.Y(n_16339)
);

AND2x2_ASAP7_75t_L g16340 ( 
.A(n_16315),
.B(n_2848),
.Y(n_16340)
);

AND2x2_ASAP7_75t_L g16341 ( 
.A(n_16319),
.B(n_16243),
.Y(n_16341)
);

AND2x2_ASAP7_75t_L g16342 ( 
.A(n_16245),
.B(n_2849),
.Y(n_16342)
);

HB1xp67_ASAP7_75t_L g16343 ( 
.A(n_16292),
.Y(n_16343)
);

AND2x2_ASAP7_75t_L g16344 ( 
.A(n_16183),
.B(n_2849),
.Y(n_16344)
);

OR2x6_ASAP7_75t_L g16345 ( 
.A(n_16228),
.B(n_2850),
.Y(n_16345)
);

OR2x2_ASAP7_75t_L g16346 ( 
.A(n_16182),
.B(n_2851),
.Y(n_16346)
);

NOR2xp33_ASAP7_75t_L g16347 ( 
.A(n_16211),
.B(n_16271),
.Y(n_16347)
);

NAND2xp5_ASAP7_75t_L g16348 ( 
.A(n_16178),
.B(n_2851),
.Y(n_16348)
);

NAND2xp5_ASAP7_75t_L g16349 ( 
.A(n_16215),
.B(n_16191),
.Y(n_16349)
);

AND2x2_ASAP7_75t_SL g16350 ( 
.A(n_16256),
.B(n_2852),
.Y(n_16350)
);

AND2x2_ASAP7_75t_L g16351 ( 
.A(n_16222),
.B(n_2852),
.Y(n_16351)
);

INVx1_ASAP7_75t_L g16352 ( 
.A(n_16223),
.Y(n_16352)
);

INVx2_ASAP7_75t_L g16353 ( 
.A(n_16292),
.Y(n_16353)
);

INVx2_ASAP7_75t_L g16354 ( 
.A(n_16221),
.Y(n_16354)
);

NAND2xp5_ASAP7_75t_L g16355 ( 
.A(n_16198),
.B(n_2853),
.Y(n_16355)
);

AND2x2_ASAP7_75t_L g16356 ( 
.A(n_16226),
.B(n_16205),
.Y(n_16356)
);

NAND2xp5_ASAP7_75t_L g16357 ( 
.A(n_16229),
.B(n_2853),
.Y(n_16357)
);

OR2x2_ASAP7_75t_L g16358 ( 
.A(n_16187),
.B(n_2854),
.Y(n_16358)
);

AND2x2_ASAP7_75t_L g16359 ( 
.A(n_16196),
.B(n_2854),
.Y(n_16359)
);

INVx1_ASAP7_75t_L g16360 ( 
.A(n_16220),
.Y(n_16360)
);

AND2x2_ASAP7_75t_L g16361 ( 
.A(n_16305),
.B(n_2855),
.Y(n_16361)
);

INVx1_ASAP7_75t_SL g16362 ( 
.A(n_16241),
.Y(n_16362)
);

AND2x2_ASAP7_75t_L g16363 ( 
.A(n_16227),
.B(n_2855),
.Y(n_16363)
);

AND2x2_ASAP7_75t_L g16364 ( 
.A(n_16242),
.B(n_2856),
.Y(n_16364)
);

INVx1_ASAP7_75t_L g16365 ( 
.A(n_16261),
.Y(n_16365)
);

AND2x2_ASAP7_75t_L g16366 ( 
.A(n_16240),
.B(n_16252),
.Y(n_16366)
);

AND2x4_ASAP7_75t_L g16367 ( 
.A(n_16188),
.B(n_2856),
.Y(n_16367)
);

AND2x2_ASAP7_75t_L g16368 ( 
.A(n_16276),
.B(n_16239),
.Y(n_16368)
);

AND2x2_ASAP7_75t_L g16369 ( 
.A(n_16250),
.B(n_2857),
.Y(n_16369)
);

INVxp67_ASAP7_75t_L g16370 ( 
.A(n_16279),
.Y(n_16370)
);

NAND2xp5_ASAP7_75t_L g16371 ( 
.A(n_16195),
.B(n_2857),
.Y(n_16371)
);

INVx1_ASAP7_75t_L g16372 ( 
.A(n_16199),
.Y(n_16372)
);

NOR2xp33_ASAP7_75t_L g16373 ( 
.A(n_16322),
.B(n_2858),
.Y(n_16373)
);

INVx2_ASAP7_75t_L g16374 ( 
.A(n_16213),
.Y(n_16374)
);

OR2x2_ASAP7_75t_L g16375 ( 
.A(n_16186),
.B(n_2858),
.Y(n_16375)
);

AND2x2_ASAP7_75t_L g16376 ( 
.A(n_16219),
.B(n_2859),
.Y(n_16376)
);

NAND2xp5_ASAP7_75t_L g16377 ( 
.A(n_16203),
.B(n_16282),
.Y(n_16377)
);

OR2x2_ASAP7_75t_L g16378 ( 
.A(n_16247),
.B(n_16209),
.Y(n_16378)
);

INVx2_ASAP7_75t_L g16379 ( 
.A(n_16300),
.Y(n_16379)
);

AND2x2_ASAP7_75t_L g16380 ( 
.A(n_16259),
.B(n_2859),
.Y(n_16380)
);

OR2x2_ASAP7_75t_L g16381 ( 
.A(n_16274),
.B(n_2860),
.Y(n_16381)
);

OR2x2_ASAP7_75t_L g16382 ( 
.A(n_16254),
.B(n_2860),
.Y(n_16382)
);

INVx1_ASAP7_75t_L g16383 ( 
.A(n_16244),
.Y(n_16383)
);

AOI21xp5_ASAP7_75t_L g16384 ( 
.A1(n_16284),
.A2(n_2861),
.B(n_2862),
.Y(n_16384)
);

INVx1_ASAP7_75t_L g16385 ( 
.A(n_16265),
.Y(n_16385)
);

OR2x2_ASAP7_75t_L g16386 ( 
.A(n_16224),
.B(n_2861),
.Y(n_16386)
);

NAND2xp5_ASAP7_75t_L g16387 ( 
.A(n_16193),
.B(n_2862),
.Y(n_16387)
);

NAND2xp5_ASAP7_75t_L g16388 ( 
.A(n_16225),
.B(n_2863),
.Y(n_16388)
);

INVx1_ASAP7_75t_L g16389 ( 
.A(n_16180),
.Y(n_16389)
);

INVx1_ASAP7_75t_SL g16390 ( 
.A(n_16303),
.Y(n_16390)
);

INVx1_ASAP7_75t_L g16391 ( 
.A(n_16317),
.Y(n_16391)
);

NAND2xp5_ASAP7_75t_L g16392 ( 
.A(n_16231),
.B(n_2863),
.Y(n_16392)
);

NAND2xp5_ASAP7_75t_L g16393 ( 
.A(n_16232),
.B(n_2864),
.Y(n_16393)
);

NOR2xp33_ASAP7_75t_L g16394 ( 
.A(n_16314),
.B(n_2864),
.Y(n_16394)
);

INVx1_ASAP7_75t_L g16395 ( 
.A(n_16318),
.Y(n_16395)
);

INVx1_ASAP7_75t_SL g16396 ( 
.A(n_16293),
.Y(n_16396)
);

NOR2x1_ASAP7_75t_L g16397 ( 
.A(n_16321),
.B(n_2865),
.Y(n_16397)
);

INVx1_ASAP7_75t_L g16398 ( 
.A(n_16281),
.Y(n_16398)
);

INVx2_ASAP7_75t_L g16399 ( 
.A(n_16277),
.Y(n_16399)
);

HB1xp67_ASAP7_75t_L g16400 ( 
.A(n_16216),
.Y(n_16400)
);

NAND2xp5_ASAP7_75t_L g16401 ( 
.A(n_16235),
.B(n_2865),
.Y(n_16401)
);

INVx1_ASAP7_75t_L g16402 ( 
.A(n_16310),
.Y(n_16402)
);

INVx2_ASAP7_75t_L g16403 ( 
.A(n_16289),
.Y(n_16403)
);

INVx1_ASAP7_75t_SL g16404 ( 
.A(n_16272),
.Y(n_16404)
);

INVx2_ASAP7_75t_L g16405 ( 
.A(n_16257),
.Y(n_16405)
);

BUFx2_ASAP7_75t_L g16406 ( 
.A(n_16217),
.Y(n_16406)
);

INVx2_ASAP7_75t_L g16407 ( 
.A(n_16306),
.Y(n_16407)
);

INVx1_ASAP7_75t_L g16408 ( 
.A(n_16218),
.Y(n_16408)
);

NOR2x1_ASAP7_75t_R g16409 ( 
.A(n_16301),
.B(n_2866),
.Y(n_16409)
);

NAND2xp5_ASAP7_75t_L g16410 ( 
.A(n_16197),
.B(n_2866),
.Y(n_16410)
);

AND2x2_ASAP7_75t_L g16411 ( 
.A(n_16268),
.B(n_2867),
.Y(n_16411)
);

OR2x2_ASAP7_75t_L g16412 ( 
.A(n_16246),
.B(n_2868),
.Y(n_16412)
);

NAND2xp5_ASAP7_75t_L g16413 ( 
.A(n_16249),
.B(n_2868),
.Y(n_16413)
);

INVx1_ASAP7_75t_L g16414 ( 
.A(n_16309),
.Y(n_16414)
);

AND2x2_ASAP7_75t_L g16415 ( 
.A(n_16263),
.B(n_2869),
.Y(n_16415)
);

OAI22xp5_ASAP7_75t_L g16416 ( 
.A1(n_16237),
.A2(n_2871),
.B1(n_2869),
.B2(n_2870),
.Y(n_16416)
);

CKINVDCx16_ASAP7_75t_R g16417 ( 
.A(n_16208),
.Y(n_16417)
);

OR2x6_ASAP7_75t_L g16418 ( 
.A(n_16234),
.B(n_2870),
.Y(n_16418)
);

AND2x2_ASAP7_75t_L g16419 ( 
.A(n_16262),
.B(n_2872),
.Y(n_16419)
);

INVx2_ASAP7_75t_L g16420 ( 
.A(n_16280),
.Y(n_16420)
);

AND2x2_ASAP7_75t_L g16421 ( 
.A(n_16248),
.B(n_2872),
.Y(n_16421)
);

AND2x4_ASAP7_75t_SL g16422 ( 
.A(n_16308),
.B(n_16267),
.Y(n_16422)
);

NOR2xp67_ASAP7_75t_L g16423 ( 
.A(n_16212),
.B(n_2873),
.Y(n_16423)
);

INVx2_ASAP7_75t_L g16424 ( 
.A(n_16260),
.Y(n_16424)
);

INVx1_ASAP7_75t_L g16425 ( 
.A(n_16297),
.Y(n_16425)
);

OR2x6_ASAP7_75t_L g16426 ( 
.A(n_16266),
.B(n_2874),
.Y(n_16426)
);

INVx1_ASAP7_75t_L g16427 ( 
.A(n_16184),
.Y(n_16427)
);

AND2x2_ASAP7_75t_L g16428 ( 
.A(n_16275),
.B(n_2875),
.Y(n_16428)
);

NAND2xp5_ASAP7_75t_L g16429 ( 
.A(n_16192),
.B(n_2875),
.Y(n_16429)
);

INVx1_ASAP7_75t_L g16430 ( 
.A(n_16251),
.Y(n_16430)
);

AND2x2_ASAP7_75t_L g16431 ( 
.A(n_16255),
.B(n_2876),
.Y(n_16431)
);

INVx1_ASAP7_75t_L g16432 ( 
.A(n_16286),
.Y(n_16432)
);

INVx1_ASAP7_75t_L g16433 ( 
.A(n_16238),
.Y(n_16433)
);

INVx1_ASAP7_75t_L g16434 ( 
.A(n_16312),
.Y(n_16434)
);

AND2x4_ASAP7_75t_L g16435 ( 
.A(n_16298),
.B(n_2876),
.Y(n_16435)
);

INVx1_ASAP7_75t_L g16436 ( 
.A(n_16299),
.Y(n_16436)
);

NAND2x1_ASAP7_75t_L g16437 ( 
.A(n_16273),
.B(n_16295),
.Y(n_16437)
);

AND2x2_ASAP7_75t_L g16438 ( 
.A(n_16313),
.B(n_2877),
.Y(n_16438)
);

NAND2xp5_ASAP7_75t_L g16439 ( 
.A(n_16316),
.B(n_2878),
.Y(n_16439)
);

INVx1_ASAP7_75t_L g16440 ( 
.A(n_16296),
.Y(n_16440)
);

INVx2_ASAP7_75t_L g16441 ( 
.A(n_16278),
.Y(n_16441)
);

OR2x2_ASAP7_75t_L g16442 ( 
.A(n_16307),
.B(n_16253),
.Y(n_16442)
);

NOR2xp33_ASAP7_75t_L g16443 ( 
.A(n_16264),
.B(n_2879),
.Y(n_16443)
);

NAND2xp5_ASAP7_75t_L g16444 ( 
.A(n_16288),
.B(n_2879),
.Y(n_16444)
);

INVx1_ASAP7_75t_L g16445 ( 
.A(n_16311),
.Y(n_16445)
);

NAND2xp5_ASAP7_75t_L g16446 ( 
.A(n_16285),
.B(n_2880),
.Y(n_16446)
);

INVx1_ASAP7_75t_L g16447 ( 
.A(n_16230),
.Y(n_16447)
);

INVx1_ASAP7_75t_L g16448 ( 
.A(n_16290),
.Y(n_16448)
);

AND3x2_ASAP7_75t_L g16449 ( 
.A(n_16269),
.B(n_16270),
.C(n_16302),
.Y(n_16449)
);

INVx1_ASAP7_75t_L g16450 ( 
.A(n_16287),
.Y(n_16450)
);

NOR2xp67_ASAP7_75t_L g16451 ( 
.A(n_16291),
.B(n_2880),
.Y(n_16451)
);

INVx1_ASAP7_75t_L g16452 ( 
.A(n_16294),
.Y(n_16452)
);

NAND3xp33_ASAP7_75t_L g16453 ( 
.A(n_16201),
.B(n_2881),
.C(n_2882),
.Y(n_16453)
);

INVx1_ASAP7_75t_L g16454 ( 
.A(n_16190),
.Y(n_16454)
);

AND2x2_ASAP7_75t_L g16455 ( 
.A(n_16206),
.B(n_2881),
.Y(n_16455)
);

INVxp67_ASAP7_75t_L g16456 ( 
.A(n_16190),
.Y(n_16456)
);

AND2x2_ASAP7_75t_L g16457 ( 
.A(n_16206),
.B(n_2883),
.Y(n_16457)
);

INVx1_ASAP7_75t_L g16458 ( 
.A(n_16190),
.Y(n_16458)
);

OR2x2_ASAP7_75t_L g16459 ( 
.A(n_16345),
.B(n_2883),
.Y(n_16459)
);

NAND2xp5_ASAP7_75t_L g16460 ( 
.A(n_16361),
.B(n_2884),
.Y(n_16460)
);

NAND2xp5_ASAP7_75t_L g16461 ( 
.A(n_16350),
.B(n_2884),
.Y(n_16461)
);

NAND2xp5_ASAP7_75t_L g16462 ( 
.A(n_16423),
.B(n_2885),
.Y(n_16462)
);

INVxp67_ASAP7_75t_L g16463 ( 
.A(n_16409),
.Y(n_16463)
);

INVx1_ASAP7_75t_L g16464 ( 
.A(n_16325),
.Y(n_16464)
);

NAND2xp5_ASAP7_75t_L g16465 ( 
.A(n_16326),
.B(n_2885),
.Y(n_16465)
);

NAND2xp5_ASAP7_75t_L g16466 ( 
.A(n_16327),
.B(n_2886),
.Y(n_16466)
);

NAND2xp5_ASAP7_75t_L g16467 ( 
.A(n_16455),
.B(n_2887),
.Y(n_16467)
);

NAND4xp25_ASAP7_75t_SL g16468 ( 
.A(n_16404),
.B(n_2889),
.C(n_2887),
.D(n_2888),
.Y(n_16468)
);

NAND2xp5_ASAP7_75t_L g16469 ( 
.A(n_16457),
.B(n_2888),
.Y(n_16469)
);

HB1xp67_ASAP7_75t_L g16470 ( 
.A(n_16345),
.Y(n_16470)
);

NAND2xp5_ASAP7_75t_L g16471 ( 
.A(n_16363),
.B(n_2889),
.Y(n_16471)
);

INVx1_ASAP7_75t_L g16472 ( 
.A(n_16343),
.Y(n_16472)
);

NAND2xp5_ASAP7_75t_L g16473 ( 
.A(n_16324),
.B(n_2890),
.Y(n_16473)
);

INVx1_ASAP7_75t_L g16474 ( 
.A(n_16415),
.Y(n_16474)
);

INVx2_ASAP7_75t_L g16475 ( 
.A(n_16426),
.Y(n_16475)
);

OR2x2_ASAP7_75t_L g16476 ( 
.A(n_16396),
.B(n_2891),
.Y(n_16476)
);

NAND2xp5_ASAP7_75t_L g16477 ( 
.A(n_16454),
.B(n_2892),
.Y(n_16477)
);

NAND2xp5_ASAP7_75t_L g16478 ( 
.A(n_16458),
.B(n_2893),
.Y(n_16478)
);

AND2x2_ASAP7_75t_L g16479 ( 
.A(n_16341),
.B(n_2893),
.Y(n_16479)
);

OR2x2_ASAP7_75t_L g16480 ( 
.A(n_16330),
.B(n_2894),
.Y(n_16480)
);

INVx1_ASAP7_75t_L g16481 ( 
.A(n_16369),
.Y(n_16481)
);

INVx1_ASAP7_75t_SL g16482 ( 
.A(n_16422),
.Y(n_16482)
);

NAND2xp33_ASAP7_75t_SL g16483 ( 
.A(n_16437),
.B(n_2895),
.Y(n_16483)
);

AND2x2_ASAP7_75t_L g16484 ( 
.A(n_16356),
.B(n_2895),
.Y(n_16484)
);

AND2x4_ASAP7_75t_L g16485 ( 
.A(n_16397),
.B(n_2896),
.Y(n_16485)
);

INVx1_ASAP7_75t_L g16486 ( 
.A(n_16426),
.Y(n_16486)
);

OAI222xp33_ASAP7_75t_L g16487 ( 
.A1(n_16456),
.A2(n_2898),
.B1(n_2900),
.B2(n_2896),
.C1(n_2897),
.C2(n_2899),
.Y(n_16487)
);

NAND2xp5_ASAP7_75t_L g16488 ( 
.A(n_16367),
.B(n_16435),
.Y(n_16488)
);

INVx2_ASAP7_75t_L g16489 ( 
.A(n_16418),
.Y(n_16489)
);

AND2x2_ASAP7_75t_L g16490 ( 
.A(n_16366),
.B(n_2897),
.Y(n_16490)
);

BUFx2_ASAP7_75t_L g16491 ( 
.A(n_16418),
.Y(n_16491)
);

NAND2xp5_ASAP7_75t_L g16492 ( 
.A(n_16342),
.B(n_2899),
.Y(n_16492)
);

INVx1_ASAP7_75t_L g16493 ( 
.A(n_16334),
.Y(n_16493)
);

INVx1_ASAP7_75t_SL g16494 ( 
.A(n_16390),
.Y(n_16494)
);

INVx2_ASAP7_75t_L g16495 ( 
.A(n_16335),
.Y(n_16495)
);

XOR2x2_ASAP7_75t_L g16496 ( 
.A(n_16333),
.B(n_2900),
.Y(n_16496)
);

INVx1_ASAP7_75t_L g16497 ( 
.A(n_16358),
.Y(n_16497)
);

NOR2xp33_ASAP7_75t_L g16498 ( 
.A(n_16362),
.B(n_16338),
.Y(n_16498)
);

NAND2xp5_ASAP7_75t_L g16499 ( 
.A(n_16419),
.B(n_2901),
.Y(n_16499)
);

NAND2xp5_ASAP7_75t_SL g16500 ( 
.A(n_16417),
.B(n_2901),
.Y(n_16500)
);

NAND2xp5_ASAP7_75t_L g16501 ( 
.A(n_16359),
.B(n_2902),
.Y(n_16501)
);

NAND4xp75_ASAP7_75t_L g16502 ( 
.A(n_16339),
.B(n_16368),
.C(n_16328),
.D(n_16329),
.Y(n_16502)
);

HB1xp67_ASAP7_75t_L g16503 ( 
.A(n_16385),
.Y(n_16503)
);

AND2x2_ASAP7_75t_L g16504 ( 
.A(n_16403),
.B(n_2903),
.Y(n_16504)
);

NAND2xp5_ASAP7_75t_L g16505 ( 
.A(n_16364),
.B(n_2903),
.Y(n_16505)
);

NAND2xp5_ASAP7_75t_L g16506 ( 
.A(n_16351),
.B(n_2904),
.Y(n_16506)
);

AND2x2_ASAP7_75t_L g16507 ( 
.A(n_16406),
.B(n_2904),
.Y(n_16507)
);

NAND2xp5_ASAP7_75t_L g16508 ( 
.A(n_16344),
.B(n_2905),
.Y(n_16508)
);

OR2x2_ASAP7_75t_L g16509 ( 
.A(n_16382),
.B(n_2905),
.Y(n_16509)
);

AND2x2_ASAP7_75t_L g16510 ( 
.A(n_16354),
.B(n_2906),
.Y(n_16510)
);

INVx1_ASAP7_75t_SL g16511 ( 
.A(n_16346),
.Y(n_16511)
);

HB1xp67_ASAP7_75t_L g16512 ( 
.A(n_16451),
.Y(n_16512)
);

NOR2xp33_ASAP7_75t_L g16513 ( 
.A(n_16365),
.B(n_2907),
.Y(n_16513)
);

AND2x2_ASAP7_75t_L g16514 ( 
.A(n_16337),
.B(n_16340),
.Y(n_16514)
);

NAND2xp5_ASAP7_75t_L g16515 ( 
.A(n_16332),
.B(n_2907),
.Y(n_16515)
);

NAND2xp5_ASAP7_75t_L g16516 ( 
.A(n_16380),
.B(n_2908),
.Y(n_16516)
);

NAND2xp5_ASAP7_75t_L g16517 ( 
.A(n_16331),
.B(n_16376),
.Y(n_16517)
);

INVx1_ASAP7_75t_L g16518 ( 
.A(n_16386),
.Y(n_16518)
);

INVx1_ASAP7_75t_L g16519 ( 
.A(n_16412),
.Y(n_16519)
);

HB1xp67_ASAP7_75t_L g16520 ( 
.A(n_16348),
.Y(n_16520)
);

AND2x2_ASAP7_75t_L g16521 ( 
.A(n_16352),
.B(n_2908),
.Y(n_16521)
);

AND2x2_ASAP7_75t_L g16522 ( 
.A(n_16428),
.B(n_2909),
.Y(n_16522)
);

BUFx2_ASAP7_75t_L g16523 ( 
.A(n_16353),
.Y(n_16523)
);

INVx2_ASAP7_75t_L g16524 ( 
.A(n_16375),
.Y(n_16524)
);

INVxp67_ASAP7_75t_L g16525 ( 
.A(n_16347),
.Y(n_16525)
);

NAND3xp33_ASAP7_75t_L g16526 ( 
.A(n_16433),
.B(n_2910),
.C(n_2911),
.Y(n_16526)
);

INVx1_ASAP7_75t_SL g16527 ( 
.A(n_16431),
.Y(n_16527)
);

AND2x2_ASAP7_75t_L g16528 ( 
.A(n_16360),
.B(n_2910),
.Y(n_16528)
);

NAND2xp5_ASAP7_75t_L g16529 ( 
.A(n_16411),
.B(n_2911),
.Y(n_16529)
);

AND3x2_ASAP7_75t_L g16530 ( 
.A(n_16323),
.B(n_2912),
.C(n_2913),
.Y(n_16530)
);

NAND2xp5_ASAP7_75t_L g16531 ( 
.A(n_16421),
.B(n_2912),
.Y(n_16531)
);

INVx1_ASAP7_75t_L g16532 ( 
.A(n_16336),
.Y(n_16532)
);

INVx1_ASAP7_75t_L g16533 ( 
.A(n_16349),
.Y(n_16533)
);

OR2x2_ASAP7_75t_L g16534 ( 
.A(n_16387),
.B(n_2913),
.Y(n_16534)
);

NOR2xp33_ASAP7_75t_L g16535 ( 
.A(n_16370),
.B(n_16402),
.Y(n_16535)
);

AND2x2_ASAP7_75t_L g16536 ( 
.A(n_16407),
.B(n_2914),
.Y(n_16536)
);

INVx1_ASAP7_75t_L g16537 ( 
.A(n_16357),
.Y(n_16537)
);

AND2x2_ASAP7_75t_L g16538 ( 
.A(n_16399),
.B(n_2914),
.Y(n_16538)
);

INVx2_ASAP7_75t_SL g16539 ( 
.A(n_16378),
.Y(n_16539)
);

OR2x2_ASAP7_75t_L g16540 ( 
.A(n_16377),
.B(n_2915),
.Y(n_16540)
);

INVx1_ASAP7_75t_L g16541 ( 
.A(n_16438),
.Y(n_16541)
);

OR2x2_ASAP7_75t_L g16542 ( 
.A(n_16371),
.B(n_2915),
.Y(n_16542)
);

INVx1_ASAP7_75t_L g16543 ( 
.A(n_16355),
.Y(n_16543)
);

INVx2_ASAP7_75t_L g16544 ( 
.A(n_16381),
.Y(n_16544)
);

NOR3xp33_ASAP7_75t_SL g16545 ( 
.A(n_16394),
.B(n_2916),
.C(n_2918),
.Y(n_16545)
);

AND2x2_ASAP7_75t_L g16546 ( 
.A(n_16414),
.B(n_2916),
.Y(n_16546)
);

INVx1_ASAP7_75t_SL g16547 ( 
.A(n_16440),
.Y(n_16547)
);

INVx1_ASAP7_75t_L g16548 ( 
.A(n_16388),
.Y(n_16548)
);

INVx1_ASAP7_75t_L g16549 ( 
.A(n_16392),
.Y(n_16549)
);

OR2x2_ASAP7_75t_L g16550 ( 
.A(n_16393),
.B(n_2918),
.Y(n_16550)
);

AND2x2_ASAP7_75t_L g16551 ( 
.A(n_16405),
.B(n_2919),
.Y(n_16551)
);

AND2x2_ASAP7_75t_L g16552 ( 
.A(n_16425),
.B(n_16432),
.Y(n_16552)
);

HB1xp67_ASAP7_75t_L g16553 ( 
.A(n_16420),
.Y(n_16553)
);

INVx1_ASAP7_75t_L g16554 ( 
.A(n_16401),
.Y(n_16554)
);

AOI22xp5_ASAP7_75t_L g16555 ( 
.A1(n_16373),
.A2(n_2922),
.B1(n_2920),
.B2(n_2921),
.Y(n_16555)
);

INVx1_ASAP7_75t_L g16556 ( 
.A(n_16413),
.Y(n_16556)
);

NAND2xp33_ASAP7_75t_SL g16557 ( 
.A(n_16400),
.B(n_2920),
.Y(n_16557)
);

INVx1_ASAP7_75t_L g16558 ( 
.A(n_16410),
.Y(n_16558)
);

NAND2xp5_ASAP7_75t_L g16559 ( 
.A(n_16389),
.B(n_2921),
.Y(n_16559)
);

INVx2_ASAP7_75t_SL g16560 ( 
.A(n_16449),
.Y(n_16560)
);

INVx1_ASAP7_75t_L g16561 ( 
.A(n_16429),
.Y(n_16561)
);

AND2x2_ASAP7_75t_L g16562 ( 
.A(n_16379),
.B(n_2922),
.Y(n_16562)
);

INVx1_ASAP7_75t_SL g16563 ( 
.A(n_16442),
.Y(n_16563)
);

INVx1_ASAP7_75t_SL g16564 ( 
.A(n_16439),
.Y(n_16564)
);

AND2x2_ASAP7_75t_L g16565 ( 
.A(n_16408),
.B(n_2923),
.Y(n_16565)
);

INVx2_ASAP7_75t_L g16566 ( 
.A(n_16391),
.Y(n_16566)
);

NAND2xp5_ASAP7_75t_L g16567 ( 
.A(n_16395),
.B(n_2923),
.Y(n_16567)
);

OR2x2_ASAP7_75t_L g16568 ( 
.A(n_16444),
.B(n_2924),
.Y(n_16568)
);

OR2x6_ASAP7_75t_L g16569 ( 
.A(n_16424),
.B(n_2925),
.Y(n_16569)
);

INVx1_ASAP7_75t_SL g16570 ( 
.A(n_16446),
.Y(n_16570)
);

NAND2xp5_ASAP7_75t_L g16571 ( 
.A(n_16416),
.B(n_2925),
.Y(n_16571)
);

AND2x2_ASAP7_75t_L g16572 ( 
.A(n_16430),
.B(n_2926),
.Y(n_16572)
);

OR2x2_ASAP7_75t_L g16573 ( 
.A(n_16453),
.B(n_2926),
.Y(n_16573)
);

AND2x2_ASAP7_75t_L g16574 ( 
.A(n_16427),
.B(n_2927),
.Y(n_16574)
);

AOI322xp5_ASAP7_75t_L g16575 ( 
.A1(n_16447),
.A2(n_2934),
.A3(n_2932),
.B1(n_2930),
.B2(n_2928),
.C1(n_2929),
.C2(n_2931),
.Y(n_16575)
);

AND2x2_ASAP7_75t_L g16576 ( 
.A(n_16374),
.B(n_2929),
.Y(n_16576)
);

INVx1_ASAP7_75t_L g16577 ( 
.A(n_16443),
.Y(n_16577)
);

INVx1_ASAP7_75t_L g16578 ( 
.A(n_16441),
.Y(n_16578)
);

INVx1_ASAP7_75t_L g16579 ( 
.A(n_16452),
.Y(n_16579)
);

INVx1_ASAP7_75t_L g16580 ( 
.A(n_16383),
.Y(n_16580)
);

AND2x2_ASAP7_75t_L g16581 ( 
.A(n_16445),
.B(n_2930),
.Y(n_16581)
);

NAND2xp5_ASAP7_75t_SL g16582 ( 
.A(n_16384),
.B(n_2931),
.Y(n_16582)
);

NAND2xp5_ASAP7_75t_L g16583 ( 
.A(n_16398),
.B(n_2932),
.Y(n_16583)
);

INVx1_ASAP7_75t_L g16584 ( 
.A(n_16450),
.Y(n_16584)
);

INVx1_ASAP7_75t_L g16585 ( 
.A(n_16485),
.Y(n_16585)
);

INVx1_ASAP7_75t_SL g16586 ( 
.A(n_16483),
.Y(n_16586)
);

CKINVDCx16_ASAP7_75t_R g16587 ( 
.A(n_16470),
.Y(n_16587)
);

INVx1_ASAP7_75t_SL g16588 ( 
.A(n_16507),
.Y(n_16588)
);

INVx1_ASAP7_75t_SL g16589 ( 
.A(n_16491),
.Y(n_16589)
);

INVx2_ASAP7_75t_SL g16590 ( 
.A(n_16459),
.Y(n_16590)
);

AOI22xp33_ASAP7_75t_L g16591 ( 
.A1(n_16560),
.A2(n_16436),
.B1(n_16448),
.B2(n_16372),
.Y(n_16591)
);

INVx1_ASAP7_75t_L g16592 ( 
.A(n_16485),
.Y(n_16592)
);

NOR2xp33_ASAP7_75t_L g16593 ( 
.A(n_16482),
.B(n_16434),
.Y(n_16593)
);

AOI22xp33_ASAP7_75t_L g16594 ( 
.A1(n_16523),
.A2(n_2937),
.B1(n_2935),
.B2(n_2936),
.Y(n_16594)
);

NAND2xp5_ASAP7_75t_L g16595 ( 
.A(n_16484),
.B(n_2935),
.Y(n_16595)
);

NOR2x1_ASAP7_75t_L g16596 ( 
.A(n_16468),
.B(n_2936),
.Y(n_16596)
);

INVx1_ASAP7_75t_SL g16597 ( 
.A(n_16490),
.Y(n_16597)
);

CKINVDCx16_ASAP7_75t_R g16598 ( 
.A(n_16514),
.Y(n_16598)
);

OAI21x1_ASAP7_75t_SL g16599 ( 
.A1(n_16462),
.A2(n_2937),
.B(n_2938),
.Y(n_16599)
);

INVx1_ASAP7_75t_SL g16600 ( 
.A(n_16479),
.Y(n_16600)
);

INVx1_ASAP7_75t_SL g16601 ( 
.A(n_16557),
.Y(n_16601)
);

INVx4_ASAP7_75t_L g16602 ( 
.A(n_16552),
.Y(n_16602)
);

NAND2xp5_ASAP7_75t_L g16603 ( 
.A(n_16530),
.B(n_2939),
.Y(n_16603)
);

INVx2_ASAP7_75t_L g16604 ( 
.A(n_16480),
.Y(n_16604)
);

AOI22xp33_ASAP7_75t_L g16605 ( 
.A1(n_16472),
.A2(n_2942),
.B1(n_2940),
.B2(n_2941),
.Y(n_16605)
);

INVx2_ASAP7_75t_L g16606 ( 
.A(n_16476),
.Y(n_16606)
);

INVx2_ASAP7_75t_L g16607 ( 
.A(n_16569),
.Y(n_16607)
);

AND2x2_ASAP7_75t_L g16608 ( 
.A(n_16572),
.B(n_2940),
.Y(n_16608)
);

INVx1_ASAP7_75t_L g16609 ( 
.A(n_16521),
.Y(n_16609)
);

OR2x2_ASAP7_75t_L g16610 ( 
.A(n_16461),
.B(n_2941),
.Y(n_16610)
);

INVx1_ASAP7_75t_L g16611 ( 
.A(n_16528),
.Y(n_16611)
);

CKINVDCx16_ASAP7_75t_R g16612 ( 
.A(n_16539),
.Y(n_16612)
);

AOI22xp33_ASAP7_75t_L g16613 ( 
.A1(n_16494),
.A2(n_2945),
.B1(n_2943),
.B2(n_2944),
.Y(n_16613)
);

INVx1_ASAP7_75t_L g16614 ( 
.A(n_16546),
.Y(n_16614)
);

AND2x4_ASAP7_75t_L g16615 ( 
.A(n_16474),
.B(n_2943),
.Y(n_16615)
);

AOI222xp33_ASAP7_75t_L g16616 ( 
.A1(n_16547),
.A2(n_2947),
.B1(n_2949),
.B2(n_2945),
.C1(n_2946),
.C2(n_2948),
.Y(n_16616)
);

NAND2xp5_ASAP7_75t_L g16617 ( 
.A(n_16510),
.B(n_2946),
.Y(n_16617)
);

AND2x2_ASAP7_75t_L g16618 ( 
.A(n_16574),
.B(n_2947),
.Y(n_16618)
);

INVx1_ASAP7_75t_SL g16619 ( 
.A(n_16522),
.Y(n_16619)
);

INVx1_ASAP7_75t_L g16620 ( 
.A(n_16504),
.Y(n_16620)
);

INVx1_ASAP7_75t_L g16621 ( 
.A(n_16565),
.Y(n_16621)
);

NOR2xp33_ASAP7_75t_L g16622 ( 
.A(n_16486),
.B(n_2948),
.Y(n_16622)
);

INVx1_ASAP7_75t_L g16623 ( 
.A(n_16503),
.Y(n_16623)
);

OR2x2_ASAP7_75t_L g16624 ( 
.A(n_16509),
.B(n_2949),
.Y(n_16624)
);

NAND2xp5_ASAP7_75t_L g16625 ( 
.A(n_16551),
.B(n_2950),
.Y(n_16625)
);

OR2x2_ASAP7_75t_L g16626 ( 
.A(n_16540),
.B(n_2950),
.Y(n_16626)
);

INVxp67_ASAP7_75t_L g16627 ( 
.A(n_16513),
.Y(n_16627)
);

HB1xp67_ASAP7_75t_L g16628 ( 
.A(n_16569),
.Y(n_16628)
);

INVx3_ASAP7_75t_L g16629 ( 
.A(n_16475),
.Y(n_16629)
);

NAND2xp33_ASAP7_75t_SL g16630 ( 
.A(n_16545),
.B(n_2951),
.Y(n_16630)
);

AND2x2_ASAP7_75t_L g16631 ( 
.A(n_16536),
.B(n_16563),
.Y(n_16631)
);

INVx1_ASAP7_75t_SL g16632 ( 
.A(n_16562),
.Y(n_16632)
);

INVx1_ASAP7_75t_SL g16633 ( 
.A(n_16576),
.Y(n_16633)
);

AND2x4_ASAP7_75t_L g16634 ( 
.A(n_16481),
.B(n_2951),
.Y(n_16634)
);

INVx1_ASAP7_75t_SL g16635 ( 
.A(n_16581),
.Y(n_16635)
);

INVx1_ASAP7_75t_SL g16636 ( 
.A(n_16538),
.Y(n_16636)
);

OR2x6_ASAP7_75t_L g16637 ( 
.A(n_16502),
.B(n_2952),
.Y(n_16637)
);

INVx1_ASAP7_75t_SL g16638 ( 
.A(n_16534),
.Y(n_16638)
);

INVx1_ASAP7_75t_L g16639 ( 
.A(n_16499),
.Y(n_16639)
);

INVx1_ASAP7_75t_L g16640 ( 
.A(n_16492),
.Y(n_16640)
);

OR2x2_ASAP7_75t_L g16641 ( 
.A(n_16460),
.B(n_2952),
.Y(n_16641)
);

AND2x4_ASAP7_75t_L g16642 ( 
.A(n_16495),
.B(n_16489),
.Y(n_16642)
);

INVx1_ASAP7_75t_L g16643 ( 
.A(n_16465),
.Y(n_16643)
);

INVx1_ASAP7_75t_L g16644 ( 
.A(n_16466),
.Y(n_16644)
);

NAND2xp5_ASAP7_75t_L g16645 ( 
.A(n_16493),
.B(n_2953),
.Y(n_16645)
);

OR2x2_ASAP7_75t_L g16646 ( 
.A(n_16471),
.B(n_2953),
.Y(n_16646)
);

AOI21xp5_ASAP7_75t_L g16647 ( 
.A1(n_16488),
.A2(n_2954),
.B(n_2955),
.Y(n_16647)
);

HB1xp67_ASAP7_75t_L g16648 ( 
.A(n_16512),
.Y(n_16648)
);

INVx2_ASAP7_75t_SL g16649 ( 
.A(n_16496),
.Y(n_16649)
);

INVx1_ASAP7_75t_L g16650 ( 
.A(n_16467),
.Y(n_16650)
);

INVx1_ASAP7_75t_L g16651 ( 
.A(n_16469),
.Y(n_16651)
);

BUFx2_ASAP7_75t_L g16652 ( 
.A(n_16463),
.Y(n_16652)
);

NAND2xp5_ASAP7_75t_SL g16653 ( 
.A(n_16566),
.B(n_2954),
.Y(n_16653)
);

AND2x4_ASAP7_75t_L g16654 ( 
.A(n_16544),
.B(n_2955),
.Y(n_16654)
);

OR2x2_ASAP7_75t_L g16655 ( 
.A(n_16501),
.B(n_2956),
.Y(n_16655)
);

HB1xp67_ASAP7_75t_L g16656 ( 
.A(n_16500),
.Y(n_16656)
);

AND2x2_ASAP7_75t_L g16657 ( 
.A(n_16527),
.B(n_2956),
.Y(n_16657)
);

NAND2xp5_ASAP7_75t_L g16658 ( 
.A(n_16511),
.B(n_2957),
.Y(n_16658)
);

INVx1_ASAP7_75t_L g16659 ( 
.A(n_16505),
.Y(n_16659)
);

AND2x2_ASAP7_75t_L g16660 ( 
.A(n_16541),
.B(n_2957),
.Y(n_16660)
);

INVx4_ASAP7_75t_L g16661 ( 
.A(n_16524),
.Y(n_16661)
);

AND2x4_ASAP7_75t_L g16662 ( 
.A(n_16518),
.B(n_2958),
.Y(n_16662)
);

INVx2_ASAP7_75t_L g16663 ( 
.A(n_16550),
.Y(n_16663)
);

AND2x4_ASAP7_75t_SL g16664 ( 
.A(n_16519),
.B(n_2958),
.Y(n_16664)
);

NAND4xp25_ASAP7_75t_L g16665 ( 
.A(n_16498),
.B(n_2962),
.C(n_2959),
.D(n_2960),
.Y(n_16665)
);

NAND2xp5_ASAP7_75t_L g16666 ( 
.A(n_16497),
.B(n_2959),
.Y(n_16666)
);

NAND2xp5_ASAP7_75t_L g16667 ( 
.A(n_16578),
.B(n_2960),
.Y(n_16667)
);

INVx1_ASAP7_75t_L g16668 ( 
.A(n_16506),
.Y(n_16668)
);

AND2x2_ASAP7_75t_L g16669 ( 
.A(n_16525),
.B(n_16533),
.Y(n_16669)
);

OR2x2_ASAP7_75t_L g16670 ( 
.A(n_16473),
.B(n_2962),
.Y(n_16670)
);

NAND2xp5_ASAP7_75t_L g16671 ( 
.A(n_16555),
.B(n_2963),
.Y(n_16671)
);

INVx2_ASAP7_75t_L g16672 ( 
.A(n_16542),
.Y(n_16672)
);

INVx2_ASAP7_75t_L g16673 ( 
.A(n_16568),
.Y(n_16673)
);

INVx2_ASAP7_75t_L g16674 ( 
.A(n_16573),
.Y(n_16674)
);

HB1xp67_ASAP7_75t_L g16675 ( 
.A(n_16487),
.Y(n_16675)
);

HB1xp67_ASAP7_75t_L g16676 ( 
.A(n_16464),
.Y(n_16676)
);

OR2x2_ASAP7_75t_L g16677 ( 
.A(n_16477),
.B(n_2963),
.Y(n_16677)
);

INVx1_ASAP7_75t_L g16678 ( 
.A(n_16516),
.Y(n_16678)
);

AND2x4_ASAP7_75t_L g16679 ( 
.A(n_16532),
.B(n_2964),
.Y(n_16679)
);

INVx2_ASAP7_75t_L g16680 ( 
.A(n_16529),
.Y(n_16680)
);

INVx1_ASAP7_75t_L g16681 ( 
.A(n_16531),
.Y(n_16681)
);

OR2x2_ASAP7_75t_L g16682 ( 
.A(n_16478),
.B(n_2964),
.Y(n_16682)
);

INVx1_ASAP7_75t_SL g16683 ( 
.A(n_16508),
.Y(n_16683)
);

AND2x2_ASAP7_75t_L g16684 ( 
.A(n_16535),
.B(n_2965),
.Y(n_16684)
);

INVx1_ASAP7_75t_L g16685 ( 
.A(n_16559),
.Y(n_16685)
);

INVx1_ASAP7_75t_SL g16686 ( 
.A(n_16567),
.Y(n_16686)
);

OR2x2_ASAP7_75t_L g16687 ( 
.A(n_16515),
.B(n_16571),
.Y(n_16687)
);

AND2x2_ASAP7_75t_L g16688 ( 
.A(n_16520),
.B(n_2965),
.Y(n_16688)
);

NOR2xp33_ASAP7_75t_R g16689 ( 
.A(n_16579),
.B(n_2966),
.Y(n_16689)
);

INVx1_ASAP7_75t_SL g16690 ( 
.A(n_16583),
.Y(n_16690)
);

NOR2xp33_ASAP7_75t_L g16691 ( 
.A(n_16526),
.B(n_2966),
.Y(n_16691)
);

INVx1_ASAP7_75t_SL g16692 ( 
.A(n_16517),
.Y(n_16692)
);

AND2x2_ASAP7_75t_L g16693 ( 
.A(n_16537),
.B(n_16564),
.Y(n_16693)
);

INVx1_ASAP7_75t_L g16694 ( 
.A(n_16553),
.Y(n_16694)
);

AND2x2_ASAP7_75t_L g16695 ( 
.A(n_16577),
.B(n_2967),
.Y(n_16695)
);

AND2x2_ASAP7_75t_L g16696 ( 
.A(n_16570),
.B(n_2968),
.Y(n_16696)
);

INVx1_ASAP7_75t_L g16697 ( 
.A(n_16584),
.Y(n_16697)
);

AND2x2_ASAP7_75t_L g16698 ( 
.A(n_16580),
.B(n_16561),
.Y(n_16698)
);

INVx1_ASAP7_75t_L g16699 ( 
.A(n_16582),
.Y(n_16699)
);

OR2x2_ASAP7_75t_L g16700 ( 
.A(n_16558),
.B(n_2968),
.Y(n_16700)
);

INVxp67_ASAP7_75t_SL g16701 ( 
.A(n_16548),
.Y(n_16701)
);

NAND2xp5_ASAP7_75t_L g16702 ( 
.A(n_16575),
.B(n_2969),
.Y(n_16702)
);

NAND2xp5_ASAP7_75t_L g16703 ( 
.A(n_16549),
.B(n_2969),
.Y(n_16703)
);

HB1xp67_ASAP7_75t_L g16704 ( 
.A(n_16554),
.Y(n_16704)
);

NOR2x1_ASAP7_75t_L g16705 ( 
.A(n_16556),
.B(n_2970),
.Y(n_16705)
);

INVx1_ASAP7_75t_L g16706 ( 
.A(n_16543),
.Y(n_16706)
);

NAND2xp5_ASAP7_75t_L g16707 ( 
.A(n_16484),
.B(n_2970),
.Y(n_16707)
);

INVx1_ASAP7_75t_SL g16708 ( 
.A(n_16483),
.Y(n_16708)
);

AND2x2_ASAP7_75t_L g16709 ( 
.A(n_16482),
.B(n_2971),
.Y(n_16709)
);

AND2x2_ASAP7_75t_L g16710 ( 
.A(n_16482),
.B(n_2971),
.Y(n_16710)
);

INVx1_ASAP7_75t_L g16711 ( 
.A(n_16485),
.Y(n_16711)
);

INVx1_ASAP7_75t_L g16712 ( 
.A(n_16485),
.Y(n_16712)
);

NOR2xp33_ASAP7_75t_SL g16713 ( 
.A(n_16482),
.B(n_2972),
.Y(n_16713)
);

INVx1_ASAP7_75t_L g16714 ( 
.A(n_16485),
.Y(n_16714)
);

BUFx2_ASAP7_75t_SL g16715 ( 
.A(n_16485),
.Y(n_16715)
);

OR2x2_ASAP7_75t_L g16716 ( 
.A(n_16612),
.B(n_2972),
.Y(n_16716)
);

INVx1_ASAP7_75t_L g16717 ( 
.A(n_16715),
.Y(n_16717)
);

INVx2_ASAP7_75t_L g16718 ( 
.A(n_16602),
.Y(n_16718)
);

NAND2xp5_ASAP7_75t_L g16719 ( 
.A(n_16587),
.B(n_2973),
.Y(n_16719)
);

AOI21xp5_ASAP7_75t_L g16720 ( 
.A1(n_16630),
.A2(n_2974),
.B(n_2975),
.Y(n_16720)
);

INVx1_ASAP7_75t_L g16721 ( 
.A(n_16709),
.Y(n_16721)
);

NAND2xp5_ASAP7_75t_L g16722 ( 
.A(n_16598),
.B(n_2975),
.Y(n_16722)
);

OA21x2_ASAP7_75t_L g16723 ( 
.A1(n_16623),
.A2(n_2976),
.B(n_2977),
.Y(n_16723)
);

NOR2x1p5_ASAP7_75t_SL g16724 ( 
.A(n_16694),
.B(n_2978),
.Y(n_16724)
);

OAI21xp33_ASAP7_75t_L g16725 ( 
.A1(n_16589),
.A2(n_2978),
.B(n_2979),
.Y(n_16725)
);

NOR2x1_ASAP7_75t_L g16726 ( 
.A(n_16705),
.B(n_2979),
.Y(n_16726)
);

AND2x2_ASAP7_75t_L g16727 ( 
.A(n_16710),
.B(n_2980),
.Y(n_16727)
);

OAI21xp33_ASAP7_75t_L g16728 ( 
.A1(n_16593),
.A2(n_2980),
.B(n_2981),
.Y(n_16728)
);

NAND2xp5_ASAP7_75t_L g16729 ( 
.A(n_16654),
.B(n_2981),
.Y(n_16729)
);

NOR2xp33_ASAP7_75t_L g16730 ( 
.A(n_16586),
.B(n_2982),
.Y(n_16730)
);

INVx2_ASAP7_75t_L g16731 ( 
.A(n_16615),
.Y(n_16731)
);

INVx1_ASAP7_75t_L g16732 ( 
.A(n_16664),
.Y(n_16732)
);

OAI21xp5_ASAP7_75t_L g16733 ( 
.A1(n_16596),
.A2(n_2983),
.B(n_2984),
.Y(n_16733)
);

INVxp67_ASAP7_75t_SL g16734 ( 
.A(n_16628),
.Y(n_16734)
);

INVx1_ASAP7_75t_L g16735 ( 
.A(n_16660),
.Y(n_16735)
);

AOI21xp33_ASAP7_75t_L g16736 ( 
.A1(n_16708),
.A2(n_2983),
.B(n_2985),
.Y(n_16736)
);

OAI322xp33_ASAP7_75t_L g16737 ( 
.A1(n_16601),
.A2(n_16697),
.A3(n_16592),
.B1(n_16711),
.B2(n_16714),
.C1(n_16712),
.C2(n_16585),
.Y(n_16737)
);

OAI21xp33_ASAP7_75t_L g16738 ( 
.A1(n_16591),
.A2(n_2985),
.B(n_2986),
.Y(n_16738)
);

XOR2x2_ASAP7_75t_L g16739 ( 
.A(n_16675),
.B(n_2986),
.Y(n_16739)
);

OR2x2_ASAP7_75t_L g16740 ( 
.A(n_16603),
.B(n_2987),
.Y(n_16740)
);

INVxp67_ASAP7_75t_L g16741 ( 
.A(n_16713),
.Y(n_16741)
);

INVx1_ASAP7_75t_L g16742 ( 
.A(n_16608),
.Y(n_16742)
);

INVx2_ASAP7_75t_SL g16743 ( 
.A(n_16634),
.Y(n_16743)
);

INVxp67_ASAP7_75t_L g16744 ( 
.A(n_16622),
.Y(n_16744)
);

OR2x2_ASAP7_75t_L g16745 ( 
.A(n_16624),
.B(n_2987),
.Y(n_16745)
);

OAI22xp5_ASAP7_75t_L g16746 ( 
.A1(n_16613),
.A2(n_2990),
.B1(n_2988),
.B2(n_2989),
.Y(n_16746)
);

INVx1_ASAP7_75t_L g16747 ( 
.A(n_16618),
.Y(n_16747)
);

NOR2xp33_ASAP7_75t_L g16748 ( 
.A(n_16665),
.B(n_2988),
.Y(n_16748)
);

INVx1_ASAP7_75t_L g16749 ( 
.A(n_16700),
.Y(n_16749)
);

NAND3xp33_ASAP7_75t_L g16750 ( 
.A(n_16648),
.B(n_2989),
.C(n_2990),
.Y(n_16750)
);

INVx2_ASAP7_75t_L g16751 ( 
.A(n_16662),
.Y(n_16751)
);

AND2x4_ASAP7_75t_L g16752 ( 
.A(n_16642),
.B(n_2991),
.Y(n_16752)
);

OAI21xp5_ASAP7_75t_L g16753 ( 
.A1(n_16658),
.A2(n_2991),
.B(n_2992),
.Y(n_16753)
);

OAI21xp5_ASAP7_75t_SL g16754 ( 
.A1(n_16597),
.A2(n_2993),
.B(n_2994),
.Y(n_16754)
);

NAND2xp5_ASAP7_75t_L g16755 ( 
.A(n_16695),
.B(n_2993),
.Y(n_16755)
);

NAND2xp33_ASAP7_75t_SL g16756 ( 
.A(n_16689),
.B(n_2994),
.Y(n_16756)
);

AND2x2_ASAP7_75t_L g16757 ( 
.A(n_16657),
.B(n_2995),
.Y(n_16757)
);

OR2x2_ASAP7_75t_L g16758 ( 
.A(n_16595),
.B(n_2995),
.Y(n_16758)
);

INVx1_ASAP7_75t_L g16759 ( 
.A(n_16684),
.Y(n_16759)
);

INVxp67_ASAP7_75t_L g16760 ( 
.A(n_16637),
.Y(n_16760)
);

AOI31xp33_ASAP7_75t_L g16761 ( 
.A1(n_16600),
.A2(n_2998),
.A3(n_2996),
.B(n_2997),
.Y(n_16761)
);

NAND2xp5_ASAP7_75t_SL g16762 ( 
.A(n_16616),
.B(n_16661),
.Y(n_16762)
);

NAND2xp5_ASAP7_75t_L g16763 ( 
.A(n_16688),
.B(n_2996),
.Y(n_16763)
);

AOI22xp5_ASAP7_75t_L g16764 ( 
.A1(n_16652),
.A2(n_2999),
.B1(n_2997),
.B2(n_2998),
.Y(n_16764)
);

AOI222xp33_ASAP7_75t_L g16765 ( 
.A1(n_16676),
.A2(n_3001),
.B1(n_3003),
.B2(n_2999),
.C1(n_3000),
.C2(n_3002),
.Y(n_16765)
);

INVx1_ASAP7_75t_L g16766 ( 
.A(n_16707),
.Y(n_16766)
);

AOI222xp33_ASAP7_75t_L g16767 ( 
.A1(n_16692),
.A2(n_3002),
.B1(n_3004),
.B2(n_3000),
.C1(n_3001),
.C2(n_3003),
.Y(n_16767)
);

INVx1_ASAP7_75t_L g16768 ( 
.A(n_16679),
.Y(n_16768)
);

NAND2xp5_ASAP7_75t_L g16769 ( 
.A(n_16619),
.B(n_3004),
.Y(n_16769)
);

NOR4xp25_ASAP7_75t_SL g16770 ( 
.A(n_16609),
.B(n_16614),
.C(n_16611),
.D(n_16620),
.Y(n_16770)
);

INVx1_ASAP7_75t_L g16771 ( 
.A(n_16637),
.Y(n_16771)
);

AOI222xp33_ASAP7_75t_L g16772 ( 
.A1(n_16588),
.A2(n_3007),
.B1(n_3009),
.B2(n_3005),
.C1(n_3006),
.C2(n_3008),
.Y(n_16772)
);

INVx1_ASAP7_75t_L g16773 ( 
.A(n_16666),
.Y(n_16773)
);

OAI32xp33_ASAP7_75t_L g16774 ( 
.A1(n_16702),
.A2(n_3008),
.A3(n_3005),
.B1(n_3007),
.B2(n_3009),
.Y(n_16774)
);

INVx1_ASAP7_75t_L g16775 ( 
.A(n_16626),
.Y(n_16775)
);

INVx1_ASAP7_75t_L g16776 ( 
.A(n_16696),
.Y(n_16776)
);

AOI22xp5_ASAP7_75t_L g16777 ( 
.A1(n_16629),
.A2(n_3012),
.B1(n_3010),
.B2(n_3011),
.Y(n_16777)
);

INVxp67_ASAP7_75t_SL g16778 ( 
.A(n_16653),
.Y(n_16778)
);

OAI21xp33_ASAP7_75t_L g16779 ( 
.A1(n_16669),
.A2(n_3011),
.B(n_3012),
.Y(n_16779)
);

INVxp67_ASAP7_75t_SL g16780 ( 
.A(n_16617),
.Y(n_16780)
);

INVx1_ASAP7_75t_SL g16781 ( 
.A(n_16631),
.Y(n_16781)
);

AOI22xp5_ASAP7_75t_L g16782 ( 
.A1(n_16649),
.A2(n_3015),
.B1(n_3013),
.B2(n_3014),
.Y(n_16782)
);

AOI22xp5_ASAP7_75t_L g16783 ( 
.A1(n_16635),
.A2(n_3015),
.B1(n_3013),
.B2(n_3014),
.Y(n_16783)
);

NOR2xp33_ASAP7_75t_L g16784 ( 
.A(n_16607),
.B(n_3016),
.Y(n_16784)
);

AOI221xp5_ASAP7_75t_L g16785 ( 
.A1(n_16701),
.A2(n_3018),
.B1(n_3016),
.B2(n_3017),
.C(n_3019),
.Y(n_16785)
);

OAI22xp5_ASAP7_75t_L g16786 ( 
.A1(n_16632),
.A2(n_3020),
.B1(n_3018),
.B2(n_3019),
.Y(n_16786)
);

NAND2xp5_ASAP7_75t_L g16787 ( 
.A(n_16594),
.B(n_3020),
.Y(n_16787)
);

INVxp67_ASAP7_75t_L g16788 ( 
.A(n_16691),
.Y(n_16788)
);

AOI221xp5_ASAP7_75t_L g16789 ( 
.A1(n_16645),
.A2(n_3023),
.B1(n_3021),
.B2(n_3022),
.C(n_3024),
.Y(n_16789)
);

INVx2_ASAP7_75t_L g16790 ( 
.A(n_16599),
.Y(n_16790)
);

OAI21xp5_ASAP7_75t_SL g16791 ( 
.A1(n_16633),
.A2(n_3021),
.B(n_3022),
.Y(n_16791)
);

NAND2xp5_ASAP7_75t_L g16792 ( 
.A(n_16647),
.B(n_3023),
.Y(n_16792)
);

OR2x2_ASAP7_75t_L g16793 ( 
.A(n_16625),
.B(n_3025),
.Y(n_16793)
);

AOI221xp5_ASAP7_75t_SL g16794 ( 
.A1(n_16627),
.A2(n_16636),
.B1(n_16638),
.B2(n_16683),
.C(n_16686),
.Y(n_16794)
);

AND2x2_ASAP7_75t_L g16795 ( 
.A(n_16590),
.B(n_3025),
.Y(n_16795)
);

AOI321xp33_ASAP7_75t_L g16796 ( 
.A1(n_16698),
.A2(n_3028),
.A3(n_3030),
.B1(n_3026),
.B2(n_3027),
.C(n_3029),
.Y(n_16796)
);

OAI21xp33_ASAP7_75t_L g16797 ( 
.A1(n_16693),
.A2(n_3026),
.B(n_3027),
.Y(n_16797)
);

NAND2xp5_ASAP7_75t_L g16798 ( 
.A(n_16605),
.B(n_3028),
.Y(n_16798)
);

AOI22xp33_ASAP7_75t_L g16799 ( 
.A1(n_16704),
.A2(n_3031),
.B1(n_3029),
.B2(n_3030),
.Y(n_16799)
);

INVx1_ASAP7_75t_L g16800 ( 
.A(n_16667),
.Y(n_16800)
);

OAI322xp33_ASAP7_75t_L g16801 ( 
.A1(n_16699),
.A2(n_3037),
.A3(n_3036),
.B1(n_3033),
.B2(n_3031),
.C1(n_3032),
.C2(n_3034),
.Y(n_16801)
);

AND2x2_ASAP7_75t_L g16802 ( 
.A(n_16621),
.B(n_3032),
.Y(n_16802)
);

INVx1_ASAP7_75t_L g16803 ( 
.A(n_16610),
.Y(n_16803)
);

AND2x2_ASAP7_75t_L g16804 ( 
.A(n_16606),
.B(n_3033),
.Y(n_16804)
);

OAI22xp5_ASAP7_75t_L g16805 ( 
.A1(n_16646),
.A2(n_3038),
.B1(n_3034),
.B2(n_3037),
.Y(n_16805)
);

OAI22xp33_ASAP7_75t_L g16806 ( 
.A1(n_16671),
.A2(n_3040),
.B1(n_3038),
.B2(n_3039),
.Y(n_16806)
);

AOI221x1_ASAP7_75t_SL g16807 ( 
.A1(n_16706),
.A2(n_3041),
.B1(n_3039),
.B2(n_3040),
.C(n_3042),
.Y(n_16807)
);

INVx1_ASAP7_75t_L g16808 ( 
.A(n_16641),
.Y(n_16808)
);

OAI22xp5_ASAP7_75t_L g16809 ( 
.A1(n_16655),
.A2(n_3043),
.B1(n_3041),
.B2(n_3042),
.Y(n_16809)
);

NAND4xp75_ASAP7_75t_L g16810 ( 
.A(n_16703),
.B(n_16639),
.C(n_16640),
.D(n_16643),
.Y(n_16810)
);

NAND2xp5_ASAP7_75t_L g16811 ( 
.A(n_16604),
.B(n_3044),
.Y(n_16811)
);

NAND2xp33_ASAP7_75t_L g16812 ( 
.A(n_16656),
.B(n_3045),
.Y(n_16812)
);

OAI322xp33_ASAP7_75t_L g16813 ( 
.A1(n_16690),
.A2(n_16687),
.A3(n_16674),
.B1(n_16685),
.B2(n_16650),
.C1(n_16651),
.C2(n_16644),
.Y(n_16813)
);

AOI221xp5_ASAP7_75t_L g16814 ( 
.A1(n_16659),
.A2(n_3048),
.B1(n_3046),
.B2(n_3047),
.C(n_3049),
.Y(n_16814)
);

OAI22xp5_ASAP7_75t_L g16815 ( 
.A1(n_16670),
.A2(n_3049),
.B1(n_3046),
.B2(n_3048),
.Y(n_16815)
);

INVx2_ASAP7_75t_SL g16816 ( 
.A(n_16677),
.Y(n_16816)
);

NAND2xp5_ASAP7_75t_L g16817 ( 
.A(n_16680),
.B(n_3050),
.Y(n_16817)
);

AND2x2_ASAP7_75t_L g16818 ( 
.A(n_16663),
.B(n_3050),
.Y(n_16818)
);

OAI22xp33_ASAP7_75t_L g16819 ( 
.A1(n_16682),
.A2(n_3053),
.B1(n_3051),
.B2(n_3052),
.Y(n_16819)
);

AOI211xp5_ASAP7_75t_L g16820 ( 
.A1(n_16668),
.A2(n_3053),
.B(n_3051),
.C(n_3052),
.Y(n_16820)
);

OAI21xp5_ASAP7_75t_L g16821 ( 
.A1(n_16678),
.A2(n_16681),
.B(n_16673),
.Y(n_16821)
);

NAND2xp5_ASAP7_75t_L g16822 ( 
.A(n_16672),
.B(n_3054),
.Y(n_16822)
);

INVx1_ASAP7_75t_L g16823 ( 
.A(n_16715),
.Y(n_16823)
);

AND2x2_ASAP7_75t_L g16824 ( 
.A(n_16709),
.B(n_3054),
.Y(n_16824)
);

INVx2_ASAP7_75t_L g16825 ( 
.A(n_16602),
.Y(n_16825)
);

INVx1_ASAP7_75t_L g16826 ( 
.A(n_16715),
.Y(n_16826)
);

INVx2_ASAP7_75t_L g16827 ( 
.A(n_16602),
.Y(n_16827)
);

AOI22xp5_ASAP7_75t_L g16828 ( 
.A1(n_16587),
.A2(n_3057),
.B1(n_3055),
.B2(n_3056),
.Y(n_16828)
);

AOI22xp5_ASAP7_75t_L g16829 ( 
.A1(n_16587),
.A2(n_3057),
.B1(n_3055),
.B2(n_3056),
.Y(n_16829)
);

NAND2xp5_ASAP7_75t_L g16830 ( 
.A(n_16587),
.B(n_3058),
.Y(n_16830)
);

OA21x2_ASAP7_75t_L g16831 ( 
.A1(n_16623),
.A2(n_3059),
.B(n_3060),
.Y(n_16831)
);

O2A1O1Ixp33_ASAP7_75t_SL g16832 ( 
.A1(n_16586),
.A2(n_3061),
.B(n_3059),
.C(n_3060),
.Y(n_16832)
);

NAND2xp5_ASAP7_75t_L g16833 ( 
.A(n_16587),
.B(n_3061),
.Y(n_16833)
);

NAND2xp5_ASAP7_75t_L g16834 ( 
.A(n_16587),
.B(n_3062),
.Y(n_16834)
);

INVx1_ASAP7_75t_L g16835 ( 
.A(n_16715),
.Y(n_16835)
);

INVx1_ASAP7_75t_L g16836 ( 
.A(n_16724),
.Y(n_16836)
);

AOI22xp33_ASAP7_75t_L g16837 ( 
.A1(n_16718),
.A2(n_3065),
.B1(n_3062),
.B2(n_3064),
.Y(n_16837)
);

NOR2xp33_ASAP7_75t_L g16838 ( 
.A(n_16716),
.B(n_3064),
.Y(n_16838)
);

OR2x2_ASAP7_75t_L g16839 ( 
.A(n_16719),
.B(n_3065),
.Y(n_16839)
);

INVx1_ASAP7_75t_L g16840 ( 
.A(n_16727),
.Y(n_16840)
);

INVx1_ASAP7_75t_L g16841 ( 
.A(n_16824),
.Y(n_16841)
);

OAI21xp5_ASAP7_75t_L g16842 ( 
.A1(n_16734),
.A2(n_3066),
.B(n_3067),
.Y(n_16842)
);

INVx1_ASAP7_75t_L g16843 ( 
.A(n_16795),
.Y(n_16843)
);

INVx1_ASAP7_75t_SL g16844 ( 
.A(n_16756),
.Y(n_16844)
);

O2A1O1Ixp33_ASAP7_75t_L g16845 ( 
.A1(n_16832),
.A2(n_3068),
.B(n_3066),
.C(n_3067),
.Y(n_16845)
);

NAND2xp5_ASAP7_75t_L g16846 ( 
.A(n_16752),
.B(n_3069),
.Y(n_16846)
);

BUFx3_ASAP7_75t_L g16847 ( 
.A(n_16825),
.Y(n_16847)
);

INVxp67_ASAP7_75t_L g16848 ( 
.A(n_16726),
.Y(n_16848)
);

OAI32xp33_ASAP7_75t_L g16849 ( 
.A1(n_16830),
.A2(n_3072),
.A3(n_3070),
.B1(n_3071),
.B2(n_3073),
.Y(n_16849)
);

AOI21xp33_ASAP7_75t_L g16850 ( 
.A1(n_16730),
.A2(n_3070),
.B(n_3071),
.Y(n_16850)
);

OAI21xp33_ASAP7_75t_SL g16851 ( 
.A1(n_16833),
.A2(n_3072),
.B(n_3073),
.Y(n_16851)
);

BUFx3_ASAP7_75t_L g16852 ( 
.A(n_16827),
.Y(n_16852)
);

INVx2_ASAP7_75t_L g16853 ( 
.A(n_16723),
.Y(n_16853)
);

INVx1_ASAP7_75t_L g16854 ( 
.A(n_16834),
.Y(n_16854)
);

INVx1_ASAP7_75t_L g16855 ( 
.A(n_16802),
.Y(n_16855)
);

INVx1_ASAP7_75t_L g16856 ( 
.A(n_16757),
.Y(n_16856)
);

AND2x2_ASAP7_75t_L g16857 ( 
.A(n_16731),
.B(n_3074),
.Y(n_16857)
);

INVxp67_ASAP7_75t_L g16858 ( 
.A(n_16784),
.Y(n_16858)
);

OAI32xp33_ASAP7_75t_L g16859 ( 
.A1(n_16722),
.A2(n_3076),
.A3(n_3074),
.B1(n_3075),
.B2(n_3077),
.Y(n_16859)
);

AND2x2_ASAP7_75t_L g16860 ( 
.A(n_16770),
.B(n_3075),
.Y(n_16860)
);

AOI22xp33_ASAP7_75t_L g16861 ( 
.A1(n_16717),
.A2(n_3078),
.B1(n_3076),
.B2(n_3077),
.Y(n_16861)
);

INVx2_ASAP7_75t_L g16862 ( 
.A(n_16723),
.Y(n_16862)
);

AOI221xp5_ASAP7_75t_SL g16863 ( 
.A1(n_16737),
.A2(n_3080),
.B1(n_3078),
.B2(n_3079),
.C(n_3081),
.Y(n_16863)
);

INVx1_ASAP7_75t_L g16864 ( 
.A(n_16804),
.Y(n_16864)
);

INVx1_ASAP7_75t_L g16865 ( 
.A(n_16818),
.Y(n_16865)
);

INVxp67_ASAP7_75t_SL g16866 ( 
.A(n_16831),
.Y(n_16866)
);

INVx2_ASAP7_75t_L g16867 ( 
.A(n_16831),
.Y(n_16867)
);

AND2x2_ASAP7_75t_L g16868 ( 
.A(n_16743),
.B(n_3079),
.Y(n_16868)
);

NOR4xp25_ASAP7_75t_SL g16869 ( 
.A(n_16762),
.B(n_3082),
.C(n_3080),
.D(n_3081),
.Y(n_16869)
);

NAND2xp5_ASAP7_75t_SL g16870 ( 
.A(n_16796),
.B(n_3083),
.Y(n_16870)
);

INVx1_ASAP7_75t_L g16871 ( 
.A(n_16745),
.Y(n_16871)
);

OAI22xp5_ASAP7_75t_L g16872 ( 
.A1(n_16781),
.A2(n_3085),
.B1(n_3083),
.B2(n_3084),
.Y(n_16872)
);

NAND2xp5_ASAP7_75t_L g16873 ( 
.A(n_16807),
.B(n_3084),
.Y(n_16873)
);

NAND2xp5_ASAP7_75t_L g16874 ( 
.A(n_16761),
.B(n_3085),
.Y(n_16874)
);

AND2x2_ASAP7_75t_L g16875 ( 
.A(n_16835),
.B(n_3086),
.Y(n_16875)
);

AOI322xp5_ASAP7_75t_L g16876 ( 
.A1(n_16823),
.A2(n_3092),
.A3(n_3091),
.B1(n_3089),
.B2(n_3086),
.C1(n_3088),
.C2(n_3090),
.Y(n_16876)
);

INVx1_ASAP7_75t_L g16877 ( 
.A(n_16739),
.Y(n_16877)
);

NOR2xp33_ASAP7_75t_L g16878 ( 
.A(n_16738),
.B(n_16725),
.Y(n_16878)
);

INVx1_ASAP7_75t_L g16879 ( 
.A(n_16769),
.Y(n_16879)
);

OAI21xp5_ASAP7_75t_L g16880 ( 
.A1(n_16720),
.A2(n_3089),
.B(n_3090),
.Y(n_16880)
);

OAI22xp5_ASAP7_75t_L g16881 ( 
.A1(n_16760),
.A2(n_3095),
.B1(n_3092),
.B2(n_3093),
.Y(n_16881)
);

INVx1_ASAP7_75t_L g16882 ( 
.A(n_16811),
.Y(n_16882)
);

NAND2xp5_ASAP7_75t_L g16883 ( 
.A(n_16820),
.B(n_3095),
.Y(n_16883)
);

NAND2xp5_ASAP7_75t_SL g16884 ( 
.A(n_16772),
.B(n_3096),
.Y(n_16884)
);

INVx1_ASAP7_75t_L g16885 ( 
.A(n_16763),
.Y(n_16885)
);

HB1xp67_ASAP7_75t_L g16886 ( 
.A(n_16733),
.Y(n_16886)
);

OAI22xp33_ASAP7_75t_SL g16887 ( 
.A1(n_16740),
.A2(n_3098),
.B1(n_3096),
.B2(n_3097),
.Y(n_16887)
);

NAND2xp5_ASAP7_75t_L g16888 ( 
.A(n_16819),
.B(n_3098),
.Y(n_16888)
);

INVx1_ASAP7_75t_L g16889 ( 
.A(n_16822),
.Y(n_16889)
);

OAI211xp5_ASAP7_75t_L g16890 ( 
.A1(n_16754),
.A2(n_3101),
.B(n_3099),
.C(n_3100),
.Y(n_16890)
);

OAI33xp33_ASAP7_75t_L g16891 ( 
.A1(n_16826),
.A2(n_3103),
.A3(n_3105),
.B1(n_3099),
.B2(n_3102),
.B3(n_3104),
.Y(n_16891)
);

NAND2xp5_ASAP7_75t_L g16892 ( 
.A(n_16828),
.B(n_16829),
.Y(n_16892)
);

INVx1_ASAP7_75t_L g16893 ( 
.A(n_16729),
.Y(n_16893)
);

INVx1_ASAP7_75t_L g16894 ( 
.A(n_16755),
.Y(n_16894)
);

NOR2x1_ASAP7_75t_L g16895 ( 
.A(n_16750),
.B(n_3102),
.Y(n_16895)
);

INVx1_ASAP7_75t_L g16896 ( 
.A(n_16817),
.Y(n_16896)
);

NAND3xp33_ASAP7_75t_SL g16897 ( 
.A(n_16791),
.B(n_3103),
.C(n_3104),
.Y(n_16897)
);

OAI22xp5_ASAP7_75t_L g16898 ( 
.A1(n_16741),
.A2(n_3107),
.B1(n_3105),
.B2(n_3106),
.Y(n_16898)
);

AND2x2_ASAP7_75t_L g16899 ( 
.A(n_16751),
.B(n_3106),
.Y(n_16899)
);

AND2x4_ASAP7_75t_SL g16900 ( 
.A(n_16732),
.B(n_3108),
.Y(n_16900)
);

NAND2xp5_ASAP7_75t_L g16901 ( 
.A(n_16779),
.B(n_3108),
.Y(n_16901)
);

AOI22xp33_ASAP7_75t_L g16902 ( 
.A1(n_16771),
.A2(n_3111),
.B1(n_3109),
.B2(n_3110),
.Y(n_16902)
);

AND2x2_ASAP7_75t_L g16903 ( 
.A(n_16742),
.B(n_3109),
.Y(n_16903)
);

OAI22xp5_ASAP7_75t_L g16904 ( 
.A1(n_16787),
.A2(n_3112),
.B1(n_3110),
.B2(n_3111),
.Y(n_16904)
);

NAND2xp33_ASAP7_75t_SL g16905 ( 
.A(n_16790),
.B(n_3112),
.Y(n_16905)
);

INVx2_ASAP7_75t_L g16906 ( 
.A(n_16758),
.Y(n_16906)
);

INVx3_ASAP7_75t_L g16907 ( 
.A(n_16793),
.Y(n_16907)
);

NOR2xp33_ASAP7_75t_L g16908 ( 
.A(n_16797),
.B(n_3113),
.Y(n_16908)
);

OAI21xp33_ASAP7_75t_L g16909 ( 
.A1(n_16721),
.A2(n_3114),
.B(n_3115),
.Y(n_16909)
);

NAND2x1_ASAP7_75t_L g16910 ( 
.A(n_16747),
.B(n_3114),
.Y(n_16910)
);

O2A1O1Ixp33_ASAP7_75t_L g16911 ( 
.A1(n_16812),
.A2(n_3117),
.B(n_3115),
.C(n_3116),
.Y(n_16911)
);

INVx1_ASAP7_75t_L g16912 ( 
.A(n_16792),
.Y(n_16912)
);

INVx1_ASAP7_75t_SL g16913 ( 
.A(n_16798),
.Y(n_16913)
);

OAI221xp5_ASAP7_75t_L g16914 ( 
.A1(n_16794),
.A2(n_3120),
.B1(n_3118),
.B2(n_3119),
.C(n_3121),
.Y(n_16914)
);

AOI32xp33_ASAP7_75t_L g16915 ( 
.A1(n_16759),
.A2(n_3121),
.A3(n_3119),
.B1(n_3120),
.B2(n_3122),
.Y(n_16915)
);

INVx1_ASAP7_75t_L g16916 ( 
.A(n_16728),
.Y(n_16916)
);

INVx1_ASAP7_75t_L g16917 ( 
.A(n_16748),
.Y(n_16917)
);

XNOR2xp5_ASAP7_75t_L g16918 ( 
.A(n_16810),
.B(n_3123),
.Y(n_16918)
);

INVx1_ASAP7_75t_SL g16919 ( 
.A(n_16768),
.Y(n_16919)
);

INVxp67_ASAP7_75t_L g16920 ( 
.A(n_16765),
.Y(n_16920)
);

INVx1_ASAP7_75t_SL g16921 ( 
.A(n_16736),
.Y(n_16921)
);

AOI22xp5_ASAP7_75t_L g16922 ( 
.A1(n_16778),
.A2(n_3125),
.B1(n_3123),
.B2(n_3124),
.Y(n_16922)
);

NOR3xp33_ASAP7_75t_L g16923 ( 
.A(n_16813),
.B(n_3124),
.C(n_3125),
.Y(n_16923)
);

INVxp33_ASAP7_75t_L g16924 ( 
.A(n_16735),
.Y(n_16924)
);

INVx1_ASAP7_75t_L g16925 ( 
.A(n_16753),
.Y(n_16925)
);

AOI22xp5_ASAP7_75t_L g16926 ( 
.A1(n_16776),
.A2(n_16746),
.B1(n_16775),
.B2(n_16744),
.Y(n_16926)
);

OAI22xp33_ASAP7_75t_L g16927 ( 
.A1(n_16782),
.A2(n_3128),
.B1(n_3126),
.B2(n_3127),
.Y(n_16927)
);

INVx1_ASAP7_75t_L g16928 ( 
.A(n_16774),
.Y(n_16928)
);

INVx1_ASAP7_75t_L g16929 ( 
.A(n_16749),
.Y(n_16929)
);

INVx1_ASAP7_75t_L g16930 ( 
.A(n_16805),
.Y(n_16930)
);

NOR2xp33_ASAP7_75t_L g16931 ( 
.A(n_16806),
.B(n_3127),
.Y(n_16931)
);

AND2x2_ASAP7_75t_L g16932 ( 
.A(n_16821),
.B(n_3128),
.Y(n_16932)
);

NAND2xp33_ASAP7_75t_L g16933 ( 
.A(n_16799),
.B(n_3129),
.Y(n_16933)
);

INVx1_ASAP7_75t_L g16934 ( 
.A(n_16809),
.Y(n_16934)
);

OAI32xp33_ASAP7_75t_L g16935 ( 
.A1(n_16788),
.A2(n_3131),
.A3(n_3129),
.B1(n_3130),
.B2(n_3132),
.Y(n_16935)
);

OAI221xp5_ASAP7_75t_SL g16936 ( 
.A1(n_16803),
.A2(n_3134),
.B1(n_3132),
.B2(n_3133),
.C(n_3135),
.Y(n_16936)
);

INVx1_ASAP7_75t_L g16937 ( 
.A(n_16815),
.Y(n_16937)
);

INVx2_ASAP7_75t_L g16938 ( 
.A(n_16816),
.Y(n_16938)
);

AOI21xp33_ASAP7_75t_L g16939 ( 
.A1(n_16780),
.A2(n_3133),
.B(n_3135),
.Y(n_16939)
);

XOR2x2_ASAP7_75t_L g16940 ( 
.A(n_16808),
.B(n_3136),
.Y(n_16940)
);

NAND2xp5_ASAP7_75t_L g16941 ( 
.A(n_16767),
.B(n_3136),
.Y(n_16941)
);

AOI21xp5_ASAP7_75t_L g16942 ( 
.A1(n_16766),
.A2(n_3137),
.B(n_3138),
.Y(n_16942)
);

INVx1_ASAP7_75t_L g16943 ( 
.A(n_16786),
.Y(n_16943)
);

NAND2xp5_ASAP7_75t_SL g16944 ( 
.A(n_16789),
.B(n_3137),
.Y(n_16944)
);

INVx2_ASAP7_75t_SL g16945 ( 
.A(n_16773),
.Y(n_16945)
);

AOI21xp33_ASAP7_75t_L g16946 ( 
.A1(n_16800),
.A2(n_3138),
.B(n_3139),
.Y(n_16946)
);

INVxp67_ASAP7_75t_SL g16947 ( 
.A(n_16783),
.Y(n_16947)
);

INVx1_ASAP7_75t_L g16948 ( 
.A(n_16764),
.Y(n_16948)
);

INVx1_ASAP7_75t_L g16949 ( 
.A(n_16866),
.Y(n_16949)
);

NOR2xp33_ASAP7_75t_L g16950 ( 
.A(n_16914),
.B(n_16801),
.Y(n_16950)
);

INVx1_ASAP7_75t_L g16951 ( 
.A(n_16853),
.Y(n_16951)
);

AND2x2_ASAP7_75t_L g16952 ( 
.A(n_16860),
.B(n_16777),
.Y(n_16952)
);

NAND2xp5_ASAP7_75t_L g16953 ( 
.A(n_16900),
.B(n_16785),
.Y(n_16953)
);

INVx1_ASAP7_75t_L g16954 ( 
.A(n_16862),
.Y(n_16954)
);

AND2x2_ASAP7_75t_L g16955 ( 
.A(n_16932),
.B(n_16919),
.Y(n_16955)
);

INVx2_ASAP7_75t_L g16956 ( 
.A(n_16867),
.Y(n_16956)
);

NAND2xp5_ASAP7_75t_L g16957 ( 
.A(n_16868),
.B(n_16814),
.Y(n_16957)
);

NAND2xp5_ASAP7_75t_L g16958 ( 
.A(n_16875),
.B(n_3139),
.Y(n_16958)
);

INVx1_ASAP7_75t_L g16959 ( 
.A(n_16910),
.Y(n_16959)
);

NAND2xp5_ASAP7_75t_L g16960 ( 
.A(n_16836),
.B(n_3140),
.Y(n_16960)
);

NAND2xp5_ASAP7_75t_L g16961 ( 
.A(n_16903),
.B(n_16863),
.Y(n_16961)
);

INVx1_ASAP7_75t_L g16962 ( 
.A(n_16918),
.Y(n_16962)
);

INVx1_ASAP7_75t_L g16963 ( 
.A(n_16940),
.Y(n_16963)
);

AND2x2_ASAP7_75t_L g16964 ( 
.A(n_16869),
.B(n_3140),
.Y(n_16964)
);

INVx1_ASAP7_75t_L g16965 ( 
.A(n_16839),
.Y(n_16965)
);

AND2x2_ASAP7_75t_L g16966 ( 
.A(n_16847),
.B(n_3141),
.Y(n_16966)
);

INVx1_ASAP7_75t_L g16967 ( 
.A(n_16873),
.Y(n_16967)
);

NAND2xp5_ASAP7_75t_L g16968 ( 
.A(n_16857),
.B(n_3142),
.Y(n_16968)
);

INVx1_ASAP7_75t_L g16969 ( 
.A(n_16874),
.Y(n_16969)
);

AND2x2_ASAP7_75t_L g16970 ( 
.A(n_16852),
.B(n_3142),
.Y(n_16970)
);

NAND2xp5_ASAP7_75t_L g16971 ( 
.A(n_16899),
.B(n_16838),
.Y(n_16971)
);

NAND2xp5_ASAP7_75t_L g16972 ( 
.A(n_16915),
.B(n_16942),
.Y(n_16972)
);

INVx1_ASAP7_75t_L g16973 ( 
.A(n_16846),
.Y(n_16973)
);

AND2x2_ASAP7_75t_L g16974 ( 
.A(n_16840),
.B(n_3143),
.Y(n_16974)
);

INVx2_ASAP7_75t_L g16975 ( 
.A(n_16841),
.Y(n_16975)
);

INVx1_ASAP7_75t_L g16976 ( 
.A(n_16845),
.Y(n_16976)
);

NAND2xp5_ASAP7_75t_L g16977 ( 
.A(n_16923),
.B(n_3143),
.Y(n_16977)
);

INVx1_ASAP7_75t_L g16978 ( 
.A(n_16941),
.Y(n_16978)
);

AND2x4_ASAP7_75t_L g16979 ( 
.A(n_16848),
.B(n_3144),
.Y(n_16979)
);

AND2x4_ASAP7_75t_SL g16980 ( 
.A(n_16856),
.B(n_3144),
.Y(n_16980)
);

INVx1_ASAP7_75t_L g16981 ( 
.A(n_16901),
.Y(n_16981)
);

INVx1_ASAP7_75t_L g16982 ( 
.A(n_16887),
.Y(n_16982)
);

OR2x2_ASAP7_75t_L g16983 ( 
.A(n_16897),
.B(n_3145),
.Y(n_16983)
);

AND2x2_ASAP7_75t_L g16984 ( 
.A(n_16920),
.B(n_3145),
.Y(n_16984)
);

OAI22xp5_ASAP7_75t_L g16985 ( 
.A1(n_16924),
.A2(n_3148),
.B1(n_3146),
.B2(n_3147),
.Y(n_16985)
);

INVx2_ASAP7_75t_L g16986 ( 
.A(n_16907),
.Y(n_16986)
);

OR2x2_ASAP7_75t_L g16987 ( 
.A(n_16870),
.B(n_16888),
.Y(n_16987)
);

OR2x2_ASAP7_75t_L g16988 ( 
.A(n_16844),
.B(n_3146),
.Y(n_16988)
);

NAND2xp5_ASAP7_75t_L g16989 ( 
.A(n_16909),
.B(n_3148),
.Y(n_16989)
);

INVx1_ASAP7_75t_L g16990 ( 
.A(n_16911),
.Y(n_16990)
);

OAI21xp5_ASAP7_75t_L g16991 ( 
.A1(n_16851),
.A2(n_3149),
.B(n_3150),
.Y(n_16991)
);

NAND2xp5_ASAP7_75t_L g16992 ( 
.A(n_16908),
.B(n_3150),
.Y(n_16992)
);

INVx1_ASAP7_75t_L g16993 ( 
.A(n_16883),
.Y(n_16993)
);

AND2x2_ASAP7_75t_L g16994 ( 
.A(n_16928),
.B(n_3151),
.Y(n_16994)
);

INVx1_ASAP7_75t_L g16995 ( 
.A(n_16895),
.Y(n_16995)
);

INVxp67_ASAP7_75t_L g16996 ( 
.A(n_16891),
.Y(n_16996)
);

INVxp33_ASAP7_75t_L g16997 ( 
.A(n_16878),
.Y(n_16997)
);

INVx1_ASAP7_75t_L g16998 ( 
.A(n_16890),
.Y(n_16998)
);

INVx1_ASAP7_75t_L g16999 ( 
.A(n_16880),
.Y(n_16999)
);

NAND2x1_ASAP7_75t_L g17000 ( 
.A(n_16907),
.B(n_3152),
.Y(n_17000)
);

INVx2_ASAP7_75t_L g17001 ( 
.A(n_16855),
.Y(n_17001)
);

NAND2xp5_ASAP7_75t_L g17002 ( 
.A(n_16927),
.B(n_16842),
.Y(n_17002)
);

INVx1_ASAP7_75t_L g17003 ( 
.A(n_16929),
.Y(n_17003)
);

NAND2xp5_ASAP7_75t_L g17004 ( 
.A(n_16871),
.B(n_3152),
.Y(n_17004)
);

NOR3xp33_ASAP7_75t_L g17005 ( 
.A(n_16938),
.B(n_3153),
.C(n_3154),
.Y(n_17005)
);

OAI21xp5_ASAP7_75t_L g17006 ( 
.A1(n_16926),
.A2(n_3153),
.B(n_3155),
.Y(n_17006)
);

AND2x2_ASAP7_75t_L g17007 ( 
.A(n_16843),
.B(n_3155),
.Y(n_17007)
);

INVx1_ASAP7_75t_L g17008 ( 
.A(n_16904),
.Y(n_17008)
);

NAND2xp5_ASAP7_75t_L g17009 ( 
.A(n_16861),
.B(n_16864),
.Y(n_17009)
);

NAND2xp5_ASAP7_75t_L g17010 ( 
.A(n_16865),
.B(n_16902),
.Y(n_17010)
);

INVx1_ASAP7_75t_L g17011 ( 
.A(n_16886),
.Y(n_17011)
);

AND2x2_ASAP7_75t_L g17012 ( 
.A(n_16947),
.B(n_3156),
.Y(n_17012)
);

NAND2xp5_ASAP7_75t_L g17013 ( 
.A(n_16872),
.B(n_3156),
.Y(n_17013)
);

AND2x2_ASAP7_75t_L g17014 ( 
.A(n_16930),
.B(n_3157),
.Y(n_17014)
);

NOR2xp33_ASAP7_75t_L g17015 ( 
.A(n_16850),
.B(n_3157),
.Y(n_17015)
);

INVxp67_ASAP7_75t_SL g17016 ( 
.A(n_16936),
.Y(n_17016)
);

NOR2xp33_ASAP7_75t_L g17017 ( 
.A(n_16884),
.B(n_3158),
.Y(n_17017)
);

INVx1_ASAP7_75t_L g17018 ( 
.A(n_16933),
.Y(n_17018)
);

AND2x2_ASAP7_75t_L g17019 ( 
.A(n_16934),
.B(n_3159),
.Y(n_17019)
);

OR2x2_ASAP7_75t_L g17020 ( 
.A(n_16892),
.B(n_3159),
.Y(n_17020)
);

NAND2xp5_ASAP7_75t_SL g17021 ( 
.A(n_16905),
.B(n_3160),
.Y(n_17021)
);

AND2x2_ASAP7_75t_L g17022 ( 
.A(n_16937),
.B(n_3160),
.Y(n_17022)
);

NAND2xp5_ASAP7_75t_SL g17023 ( 
.A(n_16945),
.B(n_3161),
.Y(n_17023)
);

OAI22xp33_ASAP7_75t_L g17024 ( 
.A1(n_16921),
.A2(n_3163),
.B1(n_3161),
.B2(n_3162),
.Y(n_17024)
);

AND2x2_ASAP7_75t_L g17025 ( 
.A(n_16877),
.B(n_3162),
.Y(n_17025)
);

INVx1_ASAP7_75t_L g17026 ( 
.A(n_16931),
.Y(n_17026)
);

NOR2x1_ASAP7_75t_L g17027 ( 
.A(n_16898),
.B(n_16881),
.Y(n_17027)
);

NAND2xp5_ASAP7_75t_L g17028 ( 
.A(n_16837),
.B(n_3163),
.Y(n_17028)
);

INVx1_ASAP7_75t_L g17029 ( 
.A(n_16943),
.Y(n_17029)
);

HB1xp67_ASAP7_75t_L g17030 ( 
.A(n_16922),
.Y(n_17030)
);

AND2x2_ASAP7_75t_L g17031 ( 
.A(n_16916),
.B(n_3164),
.Y(n_17031)
);

NAND2xp5_ASAP7_75t_L g17032 ( 
.A(n_16939),
.B(n_3165),
.Y(n_17032)
);

OR2x2_ASAP7_75t_L g17033 ( 
.A(n_16948),
.B(n_3165),
.Y(n_17033)
);

INVx1_ASAP7_75t_L g17034 ( 
.A(n_16925),
.Y(n_17034)
);

HB1xp67_ASAP7_75t_L g17035 ( 
.A(n_16935),
.Y(n_17035)
);

NAND2x1p5_ASAP7_75t_L g17036 ( 
.A(n_16906),
.B(n_3166),
.Y(n_17036)
);

OR2x2_ASAP7_75t_L g17037 ( 
.A(n_16879),
.B(n_16854),
.Y(n_17037)
);

NOR2xp33_ASAP7_75t_L g17038 ( 
.A(n_16858),
.B(n_3166),
.Y(n_17038)
);

INVx1_ASAP7_75t_SL g17039 ( 
.A(n_16946),
.Y(n_17039)
);

NAND2xp5_ASAP7_75t_L g17040 ( 
.A(n_16894),
.B(n_3167),
.Y(n_17040)
);

NAND2xp5_ASAP7_75t_SL g17041 ( 
.A(n_16913),
.B(n_3167),
.Y(n_17041)
);

NAND2xp5_ASAP7_75t_L g17042 ( 
.A(n_16885),
.B(n_3169),
.Y(n_17042)
);

INVx1_ASAP7_75t_L g17043 ( 
.A(n_16849),
.Y(n_17043)
);

INVx1_ASAP7_75t_L g17044 ( 
.A(n_16859),
.Y(n_17044)
);

INVx2_ASAP7_75t_L g17045 ( 
.A(n_16893),
.Y(n_17045)
);

NAND2xp33_ASAP7_75t_L g17046 ( 
.A(n_16917),
.B(n_3169),
.Y(n_17046)
);

INVxp67_ASAP7_75t_L g17047 ( 
.A(n_16944),
.Y(n_17047)
);

INVx2_ASAP7_75t_L g17048 ( 
.A(n_16882),
.Y(n_17048)
);

INVx1_ASAP7_75t_L g17049 ( 
.A(n_16912),
.Y(n_17049)
);

AND2x2_ASAP7_75t_L g17050 ( 
.A(n_16889),
.B(n_3170),
.Y(n_17050)
);

NAND2xp5_ASAP7_75t_L g17051 ( 
.A(n_16896),
.B(n_3171),
.Y(n_17051)
);

INVx1_ASAP7_75t_L g17052 ( 
.A(n_16876),
.Y(n_17052)
);

INVx1_ASAP7_75t_L g17053 ( 
.A(n_16866),
.Y(n_17053)
);

INVx1_ASAP7_75t_L g17054 ( 
.A(n_16866),
.Y(n_17054)
);

AND2x2_ASAP7_75t_L g17055 ( 
.A(n_16860),
.B(n_3172),
.Y(n_17055)
);

INVx2_ASAP7_75t_SL g17056 ( 
.A(n_16900),
.Y(n_17056)
);

INVx1_ASAP7_75t_L g17057 ( 
.A(n_16866),
.Y(n_17057)
);

NOR2xp33_ASAP7_75t_L g17058 ( 
.A(n_16914),
.B(n_3172),
.Y(n_17058)
);

INVx1_ASAP7_75t_L g17059 ( 
.A(n_16866),
.Y(n_17059)
);

INVx1_ASAP7_75t_L g17060 ( 
.A(n_16866),
.Y(n_17060)
);

NAND2xp5_ASAP7_75t_L g17061 ( 
.A(n_16900),
.B(n_3173),
.Y(n_17061)
);

AND2x2_ASAP7_75t_L g17062 ( 
.A(n_16860),
.B(n_3173),
.Y(n_17062)
);

NAND2xp5_ASAP7_75t_L g17063 ( 
.A(n_16900),
.B(n_3174),
.Y(n_17063)
);

INVx1_ASAP7_75t_L g17064 ( 
.A(n_16866),
.Y(n_17064)
);

AND2x2_ASAP7_75t_L g17065 ( 
.A(n_16860),
.B(n_3174),
.Y(n_17065)
);

AND2x2_ASAP7_75t_L g17066 ( 
.A(n_16860),
.B(n_3175),
.Y(n_17066)
);

INVx1_ASAP7_75t_L g17067 ( 
.A(n_16866),
.Y(n_17067)
);

NAND2xp5_ASAP7_75t_L g17068 ( 
.A(n_16900),
.B(n_3176),
.Y(n_17068)
);

NOR2xp33_ASAP7_75t_L g17069 ( 
.A(n_16914),
.B(n_3177),
.Y(n_17069)
);

NAND2xp5_ASAP7_75t_L g17070 ( 
.A(n_16900),
.B(n_3177),
.Y(n_17070)
);

INVx1_ASAP7_75t_L g17071 ( 
.A(n_16866),
.Y(n_17071)
);

INVx1_ASAP7_75t_L g17072 ( 
.A(n_16866),
.Y(n_17072)
);

HB1xp67_ASAP7_75t_L g17073 ( 
.A(n_16910),
.Y(n_17073)
);

INVx1_ASAP7_75t_L g17074 ( 
.A(n_16866),
.Y(n_17074)
);

NOR2xp33_ASAP7_75t_SL g17075 ( 
.A(n_16836),
.B(n_3178),
.Y(n_17075)
);

AND2x2_ASAP7_75t_L g17076 ( 
.A(n_16860),
.B(n_3178),
.Y(n_17076)
);

NAND2xp5_ASAP7_75t_L g17077 ( 
.A(n_17055),
.B(n_3179),
.Y(n_17077)
);

XNOR2xp5_ASAP7_75t_L g17078 ( 
.A(n_16997),
.B(n_3179),
.Y(n_17078)
);

INVx1_ASAP7_75t_L g17079 ( 
.A(n_17062),
.Y(n_17079)
);

OAI222xp33_ASAP7_75t_L g17080 ( 
.A1(n_16996),
.A2(n_3182),
.B1(n_3184),
.B2(n_3180),
.C1(n_3181),
.C2(n_3183),
.Y(n_17080)
);

OA21x2_ASAP7_75t_L g17081 ( 
.A1(n_16949),
.A2(n_3181),
.B(n_3182),
.Y(n_17081)
);

AOI211xp5_ASAP7_75t_L g17082 ( 
.A1(n_17058),
.A2(n_3186),
.B(n_3183),
.C(n_3184),
.Y(n_17082)
);

INVx1_ASAP7_75t_L g17083 ( 
.A(n_17065),
.Y(n_17083)
);

AOI222xp33_ASAP7_75t_L g17084 ( 
.A1(n_17053),
.A2(n_3188),
.B1(n_3190),
.B2(n_3186),
.C1(n_3187),
.C2(n_3189),
.Y(n_17084)
);

INVx1_ASAP7_75t_L g17085 ( 
.A(n_17066),
.Y(n_17085)
);

AND2x2_ASAP7_75t_L g17086 ( 
.A(n_16994),
.B(n_3187),
.Y(n_17086)
);

OR2x2_ASAP7_75t_L g17087 ( 
.A(n_16988),
.B(n_3188),
.Y(n_17087)
);

NOR2xp33_ASAP7_75t_L g17088 ( 
.A(n_17076),
.B(n_3189),
.Y(n_17088)
);

AOI31xp33_ASAP7_75t_L g17089 ( 
.A1(n_17073),
.A2(n_16959),
.A3(n_16964),
.B(n_17036),
.Y(n_17089)
);

NAND2xp5_ASAP7_75t_L g17090 ( 
.A(n_16980),
.B(n_3190),
.Y(n_17090)
);

XOR2x2_ASAP7_75t_L g17091 ( 
.A(n_17000),
.B(n_3191),
.Y(n_17091)
);

INVx1_ASAP7_75t_L g17092 ( 
.A(n_16960),
.Y(n_17092)
);

AOI22xp33_ASAP7_75t_L g17093 ( 
.A1(n_17003),
.A2(n_3193),
.B1(n_3191),
.B2(n_3192),
.Y(n_17093)
);

NOR3xp33_ASAP7_75t_L g17094 ( 
.A(n_17011),
.B(n_3192),
.C(n_3193),
.Y(n_17094)
);

INVx1_ASAP7_75t_SL g17095 ( 
.A(n_16966),
.Y(n_17095)
);

XOR2x2_ASAP7_75t_L g17096 ( 
.A(n_17027),
.B(n_3194),
.Y(n_17096)
);

INVx1_ASAP7_75t_L g17097 ( 
.A(n_16970),
.Y(n_17097)
);

INVx1_ASAP7_75t_L g17098 ( 
.A(n_17014),
.Y(n_17098)
);

XNOR2xp5_ASAP7_75t_L g17099 ( 
.A(n_16984),
.B(n_3194),
.Y(n_17099)
);

NAND2xp5_ASAP7_75t_SL g17100 ( 
.A(n_16975),
.B(n_3195),
.Y(n_17100)
);

INVxp67_ASAP7_75t_L g17101 ( 
.A(n_17075),
.Y(n_17101)
);

NAND2xp5_ASAP7_75t_L g17102 ( 
.A(n_17019),
.B(n_3195),
.Y(n_17102)
);

INVx1_ASAP7_75t_L g17103 ( 
.A(n_17022),
.Y(n_17103)
);

INVx1_ASAP7_75t_L g17104 ( 
.A(n_17020),
.Y(n_17104)
);

A2O1A1Ixp33_ASAP7_75t_L g17105 ( 
.A1(n_17069),
.A2(n_17054),
.B(n_17059),
.C(n_17057),
.Y(n_17105)
);

NOR2xp33_ASAP7_75t_L g17106 ( 
.A(n_17061),
.B(n_3196),
.Y(n_17106)
);

INVx1_ASAP7_75t_L g17107 ( 
.A(n_17063),
.Y(n_17107)
);

A2O1A1Ixp33_ASAP7_75t_SL g17108 ( 
.A1(n_17060),
.A2(n_17064),
.B(n_17071),
.C(n_17067),
.Y(n_17108)
);

AOI21xp33_ASAP7_75t_L g17109 ( 
.A1(n_17072),
.A2(n_3196),
.B(n_3197),
.Y(n_17109)
);

NAND2xp5_ASAP7_75t_SL g17110 ( 
.A(n_16986),
.B(n_3197),
.Y(n_17110)
);

INVx2_ASAP7_75t_L g17111 ( 
.A(n_16979),
.Y(n_17111)
);

NAND2xp5_ASAP7_75t_L g17112 ( 
.A(n_17025),
.B(n_3199),
.Y(n_17112)
);

XNOR2x1_ASAP7_75t_L g17113 ( 
.A(n_17012),
.B(n_16955),
.Y(n_17113)
);

NAND2xp5_ASAP7_75t_L g17114 ( 
.A(n_17031),
.B(n_3199),
.Y(n_17114)
);

INVxp67_ASAP7_75t_SL g17115 ( 
.A(n_17068),
.Y(n_17115)
);

INVx1_ASAP7_75t_L g17116 ( 
.A(n_17070),
.Y(n_17116)
);

XNOR2x1_ASAP7_75t_L g17117 ( 
.A(n_16987),
.B(n_3200),
.Y(n_17117)
);

OAI21xp5_ASAP7_75t_SL g17118 ( 
.A1(n_16952),
.A2(n_3200),
.B(n_3201),
.Y(n_17118)
);

AOI322xp5_ASAP7_75t_L g17119 ( 
.A1(n_16950),
.A2(n_3206),
.A3(n_3205),
.B1(n_3203),
.B2(n_3201),
.C1(n_3202),
.C2(n_3204),
.Y(n_17119)
);

O2A1O1Ixp33_ASAP7_75t_L g17120 ( 
.A1(n_17046),
.A2(n_3205),
.B(n_3203),
.C(n_3204),
.Y(n_17120)
);

NAND2xp5_ASAP7_75t_L g17121 ( 
.A(n_17038),
.B(n_3206),
.Y(n_17121)
);

AOI221xp5_ASAP7_75t_L g17122 ( 
.A1(n_17074),
.A2(n_3209),
.B1(n_3207),
.B2(n_3208),
.C(n_3210),
.Y(n_17122)
);

NAND3xp33_ASAP7_75t_L g17123 ( 
.A(n_17006),
.B(n_3208),
.C(n_3209),
.Y(n_17123)
);

NAND2xp5_ASAP7_75t_L g17124 ( 
.A(n_17005),
.B(n_3211),
.Y(n_17124)
);

A2O1A1Ixp33_ASAP7_75t_L g17125 ( 
.A1(n_17015),
.A2(n_3214),
.B(n_3212),
.C(n_3213),
.Y(n_17125)
);

INVx1_ASAP7_75t_L g17126 ( 
.A(n_17004),
.Y(n_17126)
);

CKINVDCx14_ASAP7_75t_R g17127 ( 
.A(n_17035),
.Y(n_17127)
);

OAI21xp33_ASAP7_75t_L g17128 ( 
.A1(n_17029),
.A2(n_3212),
.B(n_3213),
.Y(n_17128)
);

INVx1_ASAP7_75t_L g17129 ( 
.A(n_17033),
.Y(n_17129)
);

A2O1A1Ixp33_ASAP7_75t_L g17130 ( 
.A1(n_17017),
.A2(n_3216),
.B(n_3214),
.C(n_3215),
.Y(n_17130)
);

NAND2xp5_ASAP7_75t_L g17131 ( 
.A(n_17056),
.B(n_3216),
.Y(n_17131)
);

NAND3xp33_ASAP7_75t_L g17132 ( 
.A(n_16977),
.B(n_3217),
.C(n_3218),
.Y(n_17132)
);

INVx3_ASAP7_75t_L g17133 ( 
.A(n_16979),
.Y(n_17133)
);

INVx1_ASAP7_75t_SL g17134 ( 
.A(n_16974),
.Y(n_17134)
);

BUFx3_ASAP7_75t_L g17135 ( 
.A(n_16968),
.Y(n_17135)
);

INVx1_ASAP7_75t_L g17136 ( 
.A(n_17040),
.Y(n_17136)
);

INVx1_ASAP7_75t_L g17137 ( 
.A(n_17042),
.Y(n_17137)
);

INVx1_ASAP7_75t_L g17138 ( 
.A(n_17051),
.Y(n_17138)
);

OAI21xp5_ASAP7_75t_SL g17139 ( 
.A1(n_17034),
.A2(n_3218),
.B(n_3219),
.Y(n_17139)
);

INVx2_ASAP7_75t_L g17140 ( 
.A(n_17007),
.Y(n_17140)
);

OAI21x1_ASAP7_75t_L g17141 ( 
.A1(n_16991),
.A2(n_3219),
.B(n_3220),
.Y(n_17141)
);

INVx1_ASAP7_75t_L g17142 ( 
.A(n_16958),
.Y(n_17142)
);

AOI211xp5_ASAP7_75t_L g17143 ( 
.A1(n_17021),
.A2(n_3223),
.B(n_3221),
.C(n_3222),
.Y(n_17143)
);

INVx1_ASAP7_75t_L g17144 ( 
.A(n_16983),
.Y(n_17144)
);

OAI222xp33_ASAP7_75t_L g17145 ( 
.A1(n_17043),
.A2(n_3224),
.B1(n_3226),
.B2(n_3221),
.C1(n_3222),
.C2(n_3225),
.Y(n_17145)
);

INVx1_ASAP7_75t_SL g17146 ( 
.A(n_17050),
.Y(n_17146)
);

AND2x2_ASAP7_75t_L g17147 ( 
.A(n_16976),
.B(n_3224),
.Y(n_17147)
);

INVx1_ASAP7_75t_L g17148 ( 
.A(n_17023),
.Y(n_17148)
);

NAND2xp5_ASAP7_75t_L g17149 ( 
.A(n_16956),
.B(n_3225),
.Y(n_17149)
);

NAND2xp5_ASAP7_75t_L g17150 ( 
.A(n_16951),
.B(n_3226),
.Y(n_17150)
);

AOI22xp5_ASAP7_75t_L g17151 ( 
.A1(n_17001),
.A2(n_3229),
.B1(n_3227),
.B2(n_3228),
.Y(n_17151)
);

INVx1_ASAP7_75t_L g17152 ( 
.A(n_16989),
.Y(n_17152)
);

OAI22xp5_ASAP7_75t_L g17153 ( 
.A1(n_17052),
.A2(n_3231),
.B1(n_3228),
.B2(n_3230),
.Y(n_17153)
);

INVx2_ASAP7_75t_L g17154 ( 
.A(n_16954),
.Y(n_17154)
);

NOR2xp33_ASAP7_75t_L g17155 ( 
.A(n_16982),
.B(n_3230),
.Y(n_17155)
);

INVx1_ASAP7_75t_L g17156 ( 
.A(n_17041),
.Y(n_17156)
);

INVx1_ASAP7_75t_L g17157 ( 
.A(n_17013),
.Y(n_17157)
);

INVx1_ASAP7_75t_L g17158 ( 
.A(n_17032),
.Y(n_17158)
);

AOI21xp5_ASAP7_75t_L g17159 ( 
.A1(n_16961),
.A2(n_3232),
.B(n_3233),
.Y(n_17159)
);

O2A1O1Ixp33_ASAP7_75t_L g17160 ( 
.A1(n_16992),
.A2(n_3234),
.B(n_3232),
.C(n_3233),
.Y(n_17160)
);

AND2x2_ASAP7_75t_SL g17161 ( 
.A(n_17044),
.B(n_3234),
.Y(n_17161)
);

HB1xp67_ASAP7_75t_L g17162 ( 
.A(n_16985),
.Y(n_17162)
);

CKINVDCx20_ASAP7_75t_R g17163 ( 
.A(n_16963),
.Y(n_17163)
);

INVx1_ASAP7_75t_L g17164 ( 
.A(n_17028),
.Y(n_17164)
);

INVx2_ASAP7_75t_L g17165 ( 
.A(n_17037),
.Y(n_17165)
);

O2A1O1Ixp33_ASAP7_75t_L g17166 ( 
.A1(n_16995),
.A2(n_3237),
.B(n_3235),
.C(n_3236),
.Y(n_17166)
);

INVx1_ASAP7_75t_L g17167 ( 
.A(n_16953),
.Y(n_17167)
);

INVx1_ASAP7_75t_L g17168 ( 
.A(n_16998),
.Y(n_17168)
);

XNOR2x1_ASAP7_75t_L g17169 ( 
.A(n_16962),
.B(n_3235),
.Y(n_17169)
);

XNOR2xp5_ASAP7_75t_L g17170 ( 
.A(n_17030),
.B(n_3236),
.Y(n_17170)
);

NAND2xp5_ASAP7_75t_L g17171 ( 
.A(n_17024),
.B(n_3237),
.Y(n_17171)
);

AND2x2_ASAP7_75t_L g17172 ( 
.A(n_17016),
.B(n_3238),
.Y(n_17172)
);

INVx1_ASAP7_75t_L g17173 ( 
.A(n_16972),
.Y(n_17173)
);

OAI21xp5_ASAP7_75t_L g17174 ( 
.A1(n_17047),
.A2(n_3238),
.B(n_3239),
.Y(n_17174)
);

INVx1_ASAP7_75t_SL g17175 ( 
.A(n_16957),
.Y(n_17175)
);

INVx1_ASAP7_75t_L g17176 ( 
.A(n_16971),
.Y(n_17176)
);

OR2x2_ASAP7_75t_L g17177 ( 
.A(n_16990),
.B(n_3239),
.Y(n_17177)
);

INVx1_ASAP7_75t_L g17178 ( 
.A(n_17010),
.Y(n_17178)
);

NAND2xp5_ASAP7_75t_L g17179 ( 
.A(n_16999),
.B(n_16965),
.Y(n_17179)
);

AND2x2_ASAP7_75t_L g17180 ( 
.A(n_17018),
.B(n_3240),
.Y(n_17180)
);

AOI21xp33_ASAP7_75t_SL g17181 ( 
.A1(n_17009),
.A2(n_3240),
.B(n_3241),
.Y(n_17181)
);

NAND2xp5_ASAP7_75t_L g17182 ( 
.A(n_16973),
.B(n_3241),
.Y(n_17182)
);

OA21x2_ASAP7_75t_L g17183 ( 
.A1(n_17049),
.A2(n_3242),
.B(n_3243),
.Y(n_17183)
);

AND2x2_ASAP7_75t_L g17184 ( 
.A(n_17045),
.B(n_3242),
.Y(n_17184)
);

INVx1_ASAP7_75t_L g17185 ( 
.A(n_17002),
.Y(n_17185)
);

OAI21xp5_ASAP7_75t_SL g17186 ( 
.A1(n_17039),
.A2(n_3243),
.B(n_3244),
.Y(n_17186)
);

AND2x2_ASAP7_75t_L g17187 ( 
.A(n_17048),
.B(n_3244),
.Y(n_17187)
);

INVx1_ASAP7_75t_L g17188 ( 
.A(n_17026),
.Y(n_17188)
);

INVx1_ASAP7_75t_L g17189 ( 
.A(n_16967),
.Y(n_17189)
);

OAI21xp5_ASAP7_75t_SL g17190 ( 
.A1(n_17008),
.A2(n_3245),
.B(n_3246),
.Y(n_17190)
);

NAND2xp33_ASAP7_75t_SL g17191 ( 
.A(n_16969),
.B(n_3245),
.Y(n_17191)
);

AOI21xp5_ASAP7_75t_L g17192 ( 
.A1(n_16978),
.A2(n_3246),
.B(n_3247),
.Y(n_17192)
);

NAND2xp5_ASAP7_75t_L g17193 ( 
.A(n_16981),
.B(n_3247),
.Y(n_17193)
);

NAND2xp5_ASAP7_75t_L g17194 ( 
.A(n_16993),
.B(n_3248),
.Y(n_17194)
);

INVx2_ASAP7_75t_L g17195 ( 
.A(n_16979),
.Y(n_17195)
);

AOI222xp33_ASAP7_75t_L g17196 ( 
.A1(n_16949),
.A2(n_3250),
.B1(n_3252),
.B2(n_3248),
.C1(n_3249),
.C2(n_3251),
.Y(n_17196)
);

OAI22xp5_ASAP7_75t_L g17197 ( 
.A1(n_16996),
.A2(n_3251),
.B1(n_3249),
.B2(n_3250),
.Y(n_17197)
);

INVx1_ASAP7_75t_L g17198 ( 
.A(n_17055),
.Y(n_17198)
);

NAND2xp5_ASAP7_75t_L g17199 ( 
.A(n_17055),
.B(n_3253),
.Y(n_17199)
);

INVx1_ASAP7_75t_L g17200 ( 
.A(n_17177),
.Y(n_17200)
);

AOI221x1_ASAP7_75t_L g17201 ( 
.A1(n_17191),
.A2(n_3255),
.B1(n_3253),
.B2(n_3254),
.C(n_3256),
.Y(n_17201)
);

AOI211xp5_ASAP7_75t_L g17202 ( 
.A1(n_17181),
.A2(n_3257),
.B(n_3254),
.C(n_3255),
.Y(n_17202)
);

XNOR2x2_ASAP7_75t_L g17203 ( 
.A(n_17096),
.B(n_3257),
.Y(n_17203)
);

AND2x2_ASAP7_75t_L g17204 ( 
.A(n_17172),
.B(n_3258),
.Y(n_17204)
);

NAND2xp5_ASAP7_75t_L g17205 ( 
.A(n_17086),
.B(n_3259),
.Y(n_17205)
);

AOI211xp5_ASAP7_75t_L g17206 ( 
.A1(n_17186),
.A2(n_3261),
.B(n_3259),
.C(n_3260),
.Y(n_17206)
);

INVx1_ASAP7_75t_L g17207 ( 
.A(n_17131),
.Y(n_17207)
);

NAND2xp5_ASAP7_75t_L g17208 ( 
.A(n_17161),
.B(n_3261),
.Y(n_17208)
);

NAND4xp25_ASAP7_75t_SL g17209 ( 
.A(n_17082),
.B(n_3264),
.C(n_3262),
.D(n_3263),
.Y(n_17209)
);

INVx1_ASAP7_75t_L g17210 ( 
.A(n_17099),
.Y(n_17210)
);

OAI21xp5_ASAP7_75t_L g17211 ( 
.A1(n_17105),
.A2(n_3263),
.B(n_3264),
.Y(n_17211)
);

OAI22xp33_ASAP7_75t_L g17212 ( 
.A1(n_17089),
.A2(n_3267),
.B1(n_3265),
.B2(n_3266),
.Y(n_17212)
);

NOR2xp33_ASAP7_75t_L g17213 ( 
.A(n_17087),
.B(n_3265),
.Y(n_17213)
);

NAND3xp33_ASAP7_75t_L g17214 ( 
.A(n_17143),
.B(n_3266),
.C(n_3267),
.Y(n_17214)
);

OAI22xp33_ASAP7_75t_SL g17215 ( 
.A1(n_17077),
.A2(n_3270),
.B1(n_3268),
.B2(n_3269),
.Y(n_17215)
);

AOI21xp5_ASAP7_75t_L g17216 ( 
.A1(n_17108),
.A2(n_3268),
.B(n_3271),
.Y(n_17216)
);

INVxp67_ASAP7_75t_L g17217 ( 
.A(n_17155),
.Y(n_17217)
);

OAI21xp33_ASAP7_75t_L g17218 ( 
.A1(n_17127),
.A2(n_3271),
.B(n_3272),
.Y(n_17218)
);

OAI21xp33_ASAP7_75t_SL g17219 ( 
.A1(n_17141),
.A2(n_3272),
.B(n_3273),
.Y(n_17219)
);

OA22x2_ASAP7_75t_L g17220 ( 
.A1(n_17118),
.A2(n_17190),
.B1(n_17139),
.B2(n_17147),
.Y(n_17220)
);

AOI221xp5_ASAP7_75t_L g17221 ( 
.A1(n_17168),
.A2(n_3275),
.B1(n_3273),
.B2(n_3274),
.C(n_3276),
.Y(n_17221)
);

O2A1O1Ixp33_ASAP7_75t_L g17222 ( 
.A1(n_17199),
.A2(n_3276),
.B(n_3274),
.C(n_3275),
.Y(n_17222)
);

O2A1O1Ixp33_ASAP7_75t_L g17223 ( 
.A1(n_17154),
.A2(n_17165),
.B(n_17102),
.C(n_17114),
.Y(n_17223)
);

AOI22xp33_ASAP7_75t_SL g17224 ( 
.A1(n_17163),
.A2(n_3280),
.B1(n_3277),
.B2(n_3279),
.Y(n_17224)
);

AOI322xp5_ASAP7_75t_L g17225 ( 
.A1(n_17175),
.A2(n_3283),
.A3(n_3282),
.B1(n_3280),
.B2(n_3277),
.C1(n_3279),
.C2(n_3281),
.Y(n_17225)
);

AOI21xp5_ASAP7_75t_L g17226 ( 
.A1(n_17091),
.A2(n_3281),
.B(n_3282),
.Y(n_17226)
);

AOI22xp5_ASAP7_75t_L g17227 ( 
.A1(n_17178),
.A2(n_3285),
.B1(n_3283),
.B2(n_3284),
.Y(n_17227)
);

AOI322xp5_ASAP7_75t_L g17228 ( 
.A1(n_17185),
.A2(n_3289),
.A3(n_3288),
.B1(n_3286),
.B2(n_3284),
.C1(n_3285),
.C2(n_3287),
.Y(n_17228)
);

AOI21xp33_ASAP7_75t_L g17229 ( 
.A1(n_17120),
.A2(n_3286),
.B(n_3287),
.Y(n_17229)
);

AOI211xp5_ASAP7_75t_L g17230 ( 
.A1(n_17123),
.A2(n_3291),
.B(n_3289),
.C(n_3290),
.Y(n_17230)
);

OA22x2_ASAP7_75t_L g17231 ( 
.A1(n_17079),
.A2(n_3292),
.B1(n_3290),
.B2(n_3291),
.Y(n_17231)
);

HB1xp67_ASAP7_75t_L g17232 ( 
.A(n_17183),
.Y(n_17232)
);

AOI21xp5_ASAP7_75t_L g17233 ( 
.A1(n_17179),
.A2(n_3292),
.B(n_3293),
.Y(n_17233)
);

INVx2_ASAP7_75t_L g17234 ( 
.A(n_17183),
.Y(n_17234)
);

OAI22xp5_ASAP7_75t_L g17235 ( 
.A1(n_17132),
.A2(n_3295),
.B1(n_3293),
.B2(n_3294),
.Y(n_17235)
);

INVx2_ASAP7_75t_SL g17236 ( 
.A(n_17133),
.Y(n_17236)
);

INVx1_ASAP7_75t_L g17237 ( 
.A(n_17170),
.Y(n_17237)
);

OAI22xp33_ASAP7_75t_SL g17238 ( 
.A1(n_17171),
.A2(n_3296),
.B1(n_3294),
.B2(n_3295),
.Y(n_17238)
);

NAND2xp5_ASAP7_75t_L g17239 ( 
.A(n_17088),
.B(n_3297),
.Y(n_17239)
);

NAND3xp33_ASAP7_75t_SL g17240 ( 
.A(n_17134),
.B(n_3297),
.C(n_3298),
.Y(n_17240)
);

AND2x2_ASAP7_75t_L g17241 ( 
.A(n_17083),
.B(n_17085),
.Y(n_17241)
);

AOI22xp33_ASAP7_75t_L g17242 ( 
.A1(n_17167),
.A2(n_3300),
.B1(n_3298),
.B2(n_3299),
.Y(n_17242)
);

AOI322xp5_ASAP7_75t_L g17243 ( 
.A1(n_17173),
.A2(n_3304),
.A3(n_3303),
.B1(n_3301),
.B2(n_3299),
.C1(n_3300),
.C2(n_3302),
.Y(n_17243)
);

AOI221xp5_ASAP7_75t_L g17244 ( 
.A1(n_17101),
.A2(n_3303),
.B1(n_3301),
.B2(n_3302),
.C(n_3304),
.Y(n_17244)
);

AOI322xp5_ASAP7_75t_L g17245 ( 
.A1(n_17095),
.A2(n_3310),
.A3(n_3309),
.B1(n_3307),
.B2(n_3305),
.C1(n_3306),
.C2(n_3308),
.Y(n_17245)
);

INVxp33_ASAP7_75t_SL g17246 ( 
.A(n_17162),
.Y(n_17246)
);

OAI21xp33_ASAP7_75t_SL g17247 ( 
.A1(n_17113),
.A2(n_3305),
.B(n_3306),
.Y(n_17247)
);

INVx1_ASAP7_75t_L g17248 ( 
.A(n_17117),
.Y(n_17248)
);

NAND2xp5_ASAP7_75t_L g17249 ( 
.A(n_17094),
.B(n_3308),
.Y(n_17249)
);

AOI22xp5_ASAP7_75t_L g17250 ( 
.A1(n_17188),
.A2(n_3311),
.B1(n_3309),
.B2(n_3310),
.Y(n_17250)
);

OAI22xp5_ASAP7_75t_L g17251 ( 
.A1(n_17169),
.A2(n_17112),
.B1(n_17090),
.B2(n_17130),
.Y(n_17251)
);

AOI22xp5_ASAP7_75t_L g17252 ( 
.A1(n_17198),
.A2(n_3313),
.B1(n_3311),
.B2(n_3312),
.Y(n_17252)
);

OAI22xp5_ASAP7_75t_L g17253 ( 
.A1(n_17124),
.A2(n_3314),
.B1(n_3312),
.B2(n_3313),
.Y(n_17253)
);

INVx1_ASAP7_75t_L g17254 ( 
.A(n_17150),
.Y(n_17254)
);

OAI22xp5_ASAP7_75t_L g17255 ( 
.A1(n_17125),
.A2(n_17121),
.B1(n_17195),
.B2(n_17111),
.Y(n_17255)
);

AOI22xp5_ASAP7_75t_L g17256 ( 
.A1(n_17189),
.A2(n_3318),
.B1(n_3315),
.B2(n_3317),
.Y(n_17256)
);

AOI32xp33_ASAP7_75t_L g17257 ( 
.A1(n_17146),
.A2(n_3319),
.A3(n_3315),
.B1(n_3318),
.B2(n_3320),
.Y(n_17257)
);

AOI221xp5_ASAP7_75t_L g17258 ( 
.A1(n_17148),
.A2(n_3321),
.B1(n_3319),
.B2(n_3320),
.C(n_3322),
.Y(n_17258)
);

INVx1_ASAP7_75t_L g17259 ( 
.A(n_17149),
.Y(n_17259)
);

NAND2xp5_ASAP7_75t_L g17260 ( 
.A(n_17106),
.B(n_3321),
.Y(n_17260)
);

AOI32xp33_ASAP7_75t_L g17261 ( 
.A1(n_17176),
.A2(n_3324),
.A3(n_3322),
.B1(n_3323),
.B2(n_3325),
.Y(n_17261)
);

NAND2xp5_ASAP7_75t_L g17262 ( 
.A(n_17078),
.B(n_3323),
.Y(n_17262)
);

AOI221xp5_ASAP7_75t_L g17263 ( 
.A1(n_17156),
.A2(n_17103),
.B1(n_17098),
.B2(n_17144),
.C(n_17097),
.Y(n_17263)
);

AOI322xp5_ASAP7_75t_L g17264 ( 
.A1(n_17115),
.A2(n_3330),
.A3(n_3329),
.B1(n_3327),
.B2(n_3325),
.C1(n_3326),
.C2(n_3328),
.Y(n_17264)
);

INVx1_ASAP7_75t_L g17265 ( 
.A(n_17110),
.Y(n_17265)
);

INVxp67_ASAP7_75t_L g17266 ( 
.A(n_17184),
.Y(n_17266)
);

AOI221xp5_ASAP7_75t_L g17267 ( 
.A1(n_17160),
.A2(n_17159),
.B1(n_17129),
.B2(n_17164),
.C(n_17152),
.Y(n_17267)
);

OAI22x1_ASAP7_75t_L g17268 ( 
.A1(n_17140),
.A2(n_3328),
.B1(n_3326),
.B2(n_3327),
.Y(n_17268)
);

OAI22xp5_ASAP7_75t_L g17269 ( 
.A1(n_17104),
.A2(n_3332),
.B1(n_3330),
.B2(n_3331),
.Y(n_17269)
);

OAI22xp5_ASAP7_75t_SL g17270 ( 
.A1(n_17081),
.A2(n_3333),
.B1(n_3331),
.B2(n_3332),
.Y(n_17270)
);

OAI222xp33_ASAP7_75t_L g17271 ( 
.A1(n_17107),
.A2(n_3335),
.B1(n_3337),
.B2(n_3333),
.C1(n_3334),
.C2(n_3336),
.Y(n_17271)
);

OAI21xp5_ASAP7_75t_L g17272 ( 
.A1(n_17092),
.A2(n_17126),
.B(n_17136),
.Y(n_17272)
);

OAI31xp33_ASAP7_75t_L g17273 ( 
.A1(n_17145),
.A2(n_17080),
.A3(n_17153),
.B(n_17116),
.Y(n_17273)
);

INVx1_ASAP7_75t_L g17274 ( 
.A(n_17193),
.Y(n_17274)
);

INVx1_ASAP7_75t_L g17275 ( 
.A(n_17194),
.Y(n_17275)
);

NOR2xp33_ASAP7_75t_L g17276 ( 
.A(n_17100),
.B(n_3334),
.Y(n_17276)
);

NOR3xp33_ASAP7_75t_L g17277 ( 
.A(n_17142),
.B(n_3335),
.C(n_3336),
.Y(n_17277)
);

NAND4xp25_ASAP7_75t_SL g17278 ( 
.A(n_17166),
.B(n_3340),
.C(n_3338),
.D(n_3339),
.Y(n_17278)
);

OAI222xp33_ASAP7_75t_L g17279 ( 
.A1(n_17157),
.A2(n_3342),
.B1(n_3344),
.B2(n_3340),
.C1(n_3341),
.C2(n_3343),
.Y(n_17279)
);

AOI21xp33_ASAP7_75t_SL g17280 ( 
.A1(n_17197),
.A2(n_3341),
.B(n_3342),
.Y(n_17280)
);

INVx1_ASAP7_75t_L g17281 ( 
.A(n_17182),
.Y(n_17281)
);

O2A1O1Ixp33_ASAP7_75t_L g17282 ( 
.A1(n_17109),
.A2(n_3346),
.B(n_3344),
.C(n_3345),
.Y(n_17282)
);

INVx1_ASAP7_75t_SL g17283 ( 
.A(n_17180),
.Y(n_17283)
);

OAI221xp5_ASAP7_75t_L g17284 ( 
.A1(n_17128),
.A2(n_3348),
.B1(n_3346),
.B2(n_3347),
.C(n_3349),
.Y(n_17284)
);

NOR2xp33_ASAP7_75t_L g17285 ( 
.A(n_17135),
.B(n_3347),
.Y(n_17285)
);

AOI22xp5_ASAP7_75t_L g17286 ( 
.A1(n_17137),
.A2(n_3352),
.B1(n_3349),
.B2(n_3351),
.Y(n_17286)
);

AOI221xp5_ASAP7_75t_L g17287 ( 
.A1(n_17158),
.A2(n_3354),
.B1(n_3352),
.B2(n_3353),
.C(n_3355),
.Y(n_17287)
);

AOI22xp5_ASAP7_75t_L g17288 ( 
.A1(n_17138),
.A2(n_3356),
.B1(n_3354),
.B2(n_3355),
.Y(n_17288)
);

AOI222xp33_ASAP7_75t_L g17289 ( 
.A1(n_17174),
.A2(n_3358),
.B1(n_3360),
.B2(n_3356),
.C1(n_3357),
.C2(n_3359),
.Y(n_17289)
);

INVx1_ASAP7_75t_L g17290 ( 
.A(n_17081),
.Y(n_17290)
);

NAND2xp5_ASAP7_75t_L g17291 ( 
.A(n_17192),
.B(n_3357),
.Y(n_17291)
);

OAI21xp5_ASAP7_75t_SL g17292 ( 
.A1(n_17084),
.A2(n_17196),
.B(n_17151),
.Y(n_17292)
);

AND2x2_ASAP7_75t_L g17293 ( 
.A(n_17187),
.B(n_17093),
.Y(n_17293)
);

AOI221xp5_ASAP7_75t_L g17294 ( 
.A1(n_17122),
.A2(n_3361),
.B1(n_3358),
.B2(n_3359),
.C(n_3362),
.Y(n_17294)
);

OAI21xp33_ASAP7_75t_L g17295 ( 
.A1(n_17119),
.A2(n_3361),
.B(n_3362),
.Y(n_17295)
);

NOR3x1_ASAP7_75t_L g17296 ( 
.A(n_17186),
.B(n_3363),
.C(n_3364),
.Y(n_17296)
);

AOI21xp33_ASAP7_75t_L g17297 ( 
.A1(n_17108),
.A2(n_3363),
.B(n_3364),
.Y(n_17297)
);

OAI322xp33_ASAP7_75t_SL g17298 ( 
.A1(n_17179),
.A2(n_3370),
.A3(n_3369),
.B1(n_3367),
.B2(n_3365),
.C1(n_3366),
.C2(n_3368),
.Y(n_17298)
);

OAI21xp33_ASAP7_75t_SL g17299 ( 
.A1(n_17089),
.A2(n_3365),
.B(n_3366),
.Y(n_17299)
);

AOI22xp5_ASAP7_75t_L g17300 ( 
.A1(n_17127),
.A2(n_3372),
.B1(n_3369),
.B2(n_3371),
.Y(n_17300)
);

A2O1A1Ixp33_ASAP7_75t_L g17301 ( 
.A1(n_17160),
.A2(n_3373),
.B(n_3371),
.C(n_3372),
.Y(n_17301)
);

INVxp67_ASAP7_75t_L g17302 ( 
.A(n_17155),
.Y(n_17302)
);

AOI22xp5_ASAP7_75t_L g17303 ( 
.A1(n_17127),
.A2(n_3376),
.B1(n_3374),
.B2(n_3375),
.Y(n_17303)
);

INVx1_ASAP7_75t_L g17304 ( 
.A(n_17177),
.Y(n_17304)
);

O2A1O1Ixp33_ASAP7_75t_L g17305 ( 
.A1(n_17108),
.A2(n_3378),
.B(n_3375),
.C(n_3377),
.Y(n_17305)
);

AND2x2_ASAP7_75t_L g17306 ( 
.A(n_17172),
.B(n_3377),
.Y(n_17306)
);

NAND2xp5_ASAP7_75t_L g17307 ( 
.A(n_17086),
.B(n_3378),
.Y(n_17307)
);

INVx2_ASAP7_75t_L g17308 ( 
.A(n_17183),
.Y(n_17308)
);

AOI221xp5_ASAP7_75t_L g17309 ( 
.A1(n_17089),
.A2(n_3381),
.B1(n_3379),
.B2(n_3380),
.C(n_3382),
.Y(n_17309)
);

INVx1_ASAP7_75t_L g17310 ( 
.A(n_17177),
.Y(n_17310)
);

AND2x2_ASAP7_75t_L g17311 ( 
.A(n_17172),
.B(n_3379),
.Y(n_17311)
);

INVx1_ASAP7_75t_SL g17312 ( 
.A(n_17086),
.Y(n_17312)
);

AOI211xp5_ASAP7_75t_L g17313 ( 
.A1(n_17181),
.A2(n_3383),
.B(n_3380),
.C(n_3381),
.Y(n_17313)
);

AOI22xp5_ASAP7_75t_L g17314 ( 
.A1(n_17127),
.A2(n_3385),
.B1(n_3383),
.B2(n_3384),
.Y(n_17314)
);

OAI22xp33_ASAP7_75t_L g17315 ( 
.A1(n_17089),
.A2(n_3386),
.B1(n_3384),
.B2(n_3385),
.Y(n_17315)
);

INVx1_ASAP7_75t_L g17316 ( 
.A(n_17177),
.Y(n_17316)
);

OAI221xp5_ASAP7_75t_L g17317 ( 
.A1(n_17108),
.A2(n_3388),
.B1(n_3386),
.B2(n_3387),
.C(n_3389),
.Y(n_17317)
);

OAI221xp5_ASAP7_75t_L g17318 ( 
.A1(n_17108),
.A2(n_3391),
.B1(n_3387),
.B2(n_3390),
.C(n_3392),
.Y(n_17318)
);

NOR2xp33_ASAP7_75t_L g17319 ( 
.A(n_17131),
.B(n_3390),
.Y(n_17319)
);

XOR2xp5_ASAP7_75t_L g17320 ( 
.A(n_17246),
.B(n_3392),
.Y(n_17320)
);

NAND2xp5_ASAP7_75t_SL g17321 ( 
.A(n_17238),
.B(n_3393),
.Y(n_17321)
);

INVx2_ASAP7_75t_SL g17322 ( 
.A(n_17234),
.Y(n_17322)
);

INVx1_ASAP7_75t_L g17323 ( 
.A(n_17232),
.Y(n_17323)
);

HB1xp67_ASAP7_75t_L g17324 ( 
.A(n_17268),
.Y(n_17324)
);

NOR2x1_ASAP7_75t_L g17325 ( 
.A(n_17290),
.B(n_3393),
.Y(n_17325)
);

INVx2_ASAP7_75t_SL g17326 ( 
.A(n_17308),
.Y(n_17326)
);

NAND2xp5_ASAP7_75t_L g17327 ( 
.A(n_17204),
.B(n_3394),
.Y(n_17327)
);

INVxp67_ASAP7_75t_SL g17328 ( 
.A(n_17270),
.Y(n_17328)
);

INVx1_ASAP7_75t_L g17329 ( 
.A(n_17205),
.Y(n_17329)
);

HB1xp67_ASAP7_75t_L g17330 ( 
.A(n_17231),
.Y(n_17330)
);

NOR3xp33_ASAP7_75t_L g17331 ( 
.A(n_17263),
.B(n_3394),
.C(n_3395),
.Y(n_17331)
);

AND2x2_ASAP7_75t_L g17332 ( 
.A(n_17241),
.B(n_3396),
.Y(n_17332)
);

NAND2xp5_ASAP7_75t_SL g17333 ( 
.A(n_17212),
.B(n_3396),
.Y(n_17333)
);

INVx1_ASAP7_75t_SL g17334 ( 
.A(n_17306),
.Y(n_17334)
);

NAND2xp5_ASAP7_75t_L g17335 ( 
.A(n_17311),
.B(n_3397),
.Y(n_17335)
);

XNOR2x1_ASAP7_75t_L g17336 ( 
.A(n_17203),
.B(n_3397),
.Y(n_17336)
);

NAND2xp5_ASAP7_75t_L g17337 ( 
.A(n_17216),
.B(n_3398),
.Y(n_17337)
);

OAI21xp33_ASAP7_75t_L g17338 ( 
.A1(n_17236),
.A2(n_3398),
.B(n_3399),
.Y(n_17338)
);

NAND2xp5_ASAP7_75t_SL g17339 ( 
.A(n_17315),
.B(n_17289),
.Y(n_17339)
);

AND2x2_ASAP7_75t_L g17340 ( 
.A(n_17296),
.B(n_3399),
.Y(n_17340)
);

NOR2xp33_ASAP7_75t_L g17341 ( 
.A(n_17299),
.B(n_3400),
.Y(n_17341)
);

NAND2xp5_ASAP7_75t_L g17342 ( 
.A(n_17218),
.B(n_3400),
.Y(n_17342)
);

NOR2xp33_ASAP7_75t_L g17343 ( 
.A(n_17247),
.B(n_3401),
.Y(n_17343)
);

INVx1_ASAP7_75t_L g17344 ( 
.A(n_17307),
.Y(n_17344)
);

NAND2xp5_ASAP7_75t_SL g17345 ( 
.A(n_17206),
.B(n_3401),
.Y(n_17345)
);

INVx1_ASAP7_75t_L g17346 ( 
.A(n_17305),
.Y(n_17346)
);

INVx1_ASAP7_75t_L g17347 ( 
.A(n_17208),
.Y(n_17347)
);

NAND2xp5_ASAP7_75t_L g17348 ( 
.A(n_17213),
.B(n_3402),
.Y(n_17348)
);

NAND2xp5_ASAP7_75t_SL g17349 ( 
.A(n_17309),
.B(n_3402),
.Y(n_17349)
);

NAND2xp5_ASAP7_75t_L g17350 ( 
.A(n_17319),
.B(n_3403),
.Y(n_17350)
);

NAND2xp5_ASAP7_75t_L g17351 ( 
.A(n_17202),
.B(n_3403),
.Y(n_17351)
);

NAND2xp5_ASAP7_75t_L g17352 ( 
.A(n_17313),
.B(n_3404),
.Y(n_17352)
);

AND2x2_ASAP7_75t_L g17353 ( 
.A(n_17211),
.B(n_3404),
.Y(n_17353)
);

NAND2xp5_ASAP7_75t_L g17354 ( 
.A(n_17277),
.B(n_3405),
.Y(n_17354)
);

AOI21xp5_ASAP7_75t_L g17355 ( 
.A1(n_17297),
.A2(n_3405),
.B(n_3407),
.Y(n_17355)
);

NOR2xp33_ASAP7_75t_L g17356 ( 
.A(n_17219),
.B(n_17317),
.Y(n_17356)
);

INVx2_ASAP7_75t_L g17357 ( 
.A(n_17220),
.Y(n_17357)
);

NAND2xp5_ASAP7_75t_L g17358 ( 
.A(n_17233),
.B(n_17300),
.Y(n_17358)
);

NAND2xp33_ASAP7_75t_SL g17359 ( 
.A(n_17291),
.B(n_3407),
.Y(n_17359)
);

INVx1_ASAP7_75t_SL g17360 ( 
.A(n_17262),
.Y(n_17360)
);

AND2x2_ASAP7_75t_L g17361 ( 
.A(n_17312),
.B(n_3408),
.Y(n_17361)
);

INVx1_ASAP7_75t_L g17362 ( 
.A(n_17318),
.Y(n_17362)
);

INVx1_ASAP7_75t_L g17363 ( 
.A(n_17239),
.Y(n_17363)
);

INVx1_ASAP7_75t_L g17364 ( 
.A(n_17249),
.Y(n_17364)
);

NAND2xp5_ASAP7_75t_L g17365 ( 
.A(n_17303),
.B(n_3408),
.Y(n_17365)
);

NAND2xp5_ASAP7_75t_L g17366 ( 
.A(n_17314),
.B(n_17215),
.Y(n_17366)
);

AND2x2_ASAP7_75t_L g17367 ( 
.A(n_17283),
.B(n_3409),
.Y(n_17367)
);

NAND2xp5_ASAP7_75t_L g17368 ( 
.A(n_17226),
.B(n_3410),
.Y(n_17368)
);

NAND2xp5_ASAP7_75t_L g17369 ( 
.A(n_17280),
.B(n_3410),
.Y(n_17369)
);

OAI211xp5_ASAP7_75t_L g17370 ( 
.A1(n_17273),
.A2(n_3413),
.B(n_3411),
.C(n_3412),
.Y(n_17370)
);

INVx2_ASAP7_75t_SL g17371 ( 
.A(n_17293),
.Y(n_17371)
);

NAND2xp33_ASAP7_75t_SL g17372 ( 
.A(n_17260),
.B(n_3412),
.Y(n_17372)
);

AOI221xp5_ASAP7_75t_SL g17373 ( 
.A1(n_17295),
.A2(n_3416),
.B1(n_3414),
.B2(n_3415),
.C(n_3417),
.Y(n_17373)
);

NAND3xp33_ASAP7_75t_L g17374 ( 
.A(n_17230),
.B(n_3414),
.C(n_3415),
.Y(n_17374)
);

NOR2xp33_ASAP7_75t_L g17375 ( 
.A(n_17209),
.B(n_3416),
.Y(n_17375)
);

INVxp67_ASAP7_75t_L g17376 ( 
.A(n_17285),
.Y(n_17376)
);

NAND2xp5_ASAP7_75t_L g17377 ( 
.A(n_17201),
.B(n_3417),
.Y(n_17377)
);

NOR2xp33_ASAP7_75t_L g17378 ( 
.A(n_17278),
.B(n_17276),
.Y(n_17378)
);

INVx1_ASAP7_75t_SL g17379 ( 
.A(n_17224),
.Y(n_17379)
);

NOR2x1_ASAP7_75t_SL g17380 ( 
.A(n_17240),
.B(n_3418),
.Y(n_17380)
);

INVx1_ASAP7_75t_L g17381 ( 
.A(n_17282),
.Y(n_17381)
);

INVx1_ASAP7_75t_SL g17382 ( 
.A(n_17253),
.Y(n_17382)
);

NAND2xp5_ASAP7_75t_L g17383 ( 
.A(n_17257),
.B(n_3418),
.Y(n_17383)
);

NAND2xp5_ASAP7_75t_L g17384 ( 
.A(n_17261),
.B(n_3419),
.Y(n_17384)
);

NOR3xp33_ASAP7_75t_L g17385 ( 
.A(n_17255),
.B(n_3419),
.C(n_3420),
.Y(n_17385)
);

NAND2xp5_ASAP7_75t_L g17386 ( 
.A(n_17301),
.B(n_3421),
.Y(n_17386)
);

NOR2x1_ASAP7_75t_L g17387 ( 
.A(n_17265),
.B(n_3421),
.Y(n_17387)
);

NAND2xp5_ASAP7_75t_SL g17388 ( 
.A(n_17294),
.B(n_3422),
.Y(n_17388)
);

NAND2xp5_ASAP7_75t_L g17389 ( 
.A(n_17235),
.B(n_3422),
.Y(n_17389)
);

NOR3xp33_ASAP7_75t_L g17390 ( 
.A(n_17223),
.B(n_3423),
.C(n_3424),
.Y(n_17390)
);

INVx1_ASAP7_75t_L g17391 ( 
.A(n_17214),
.Y(n_17391)
);

NAND2xp5_ASAP7_75t_L g17392 ( 
.A(n_17222),
.B(n_3423),
.Y(n_17392)
);

INVx1_ASAP7_75t_L g17393 ( 
.A(n_17284),
.Y(n_17393)
);

OAI22xp5_ASAP7_75t_L g17394 ( 
.A1(n_17266),
.A2(n_3426),
.B1(n_3424),
.B2(n_3425),
.Y(n_17394)
);

AND2x4_ASAP7_75t_SL g17395 ( 
.A(n_17237),
.B(n_3426),
.Y(n_17395)
);

INVx1_ASAP7_75t_SL g17396 ( 
.A(n_17229),
.Y(n_17396)
);

AND2x2_ASAP7_75t_L g17397 ( 
.A(n_17200),
.B(n_3427),
.Y(n_17397)
);

INVx1_ASAP7_75t_L g17398 ( 
.A(n_17304),
.Y(n_17398)
);

NAND2xp5_ASAP7_75t_L g17399 ( 
.A(n_17310),
.B(n_17316),
.Y(n_17399)
);

NAND2xp5_ASAP7_75t_L g17400 ( 
.A(n_17242),
.B(n_3427),
.Y(n_17400)
);

NAND2xp5_ASAP7_75t_L g17401 ( 
.A(n_17292),
.B(n_3428),
.Y(n_17401)
);

OR2x2_ASAP7_75t_L g17402 ( 
.A(n_17210),
.B(n_3428),
.Y(n_17402)
);

NAND2xp5_ASAP7_75t_L g17403 ( 
.A(n_17227),
.B(n_3429),
.Y(n_17403)
);

INVxp67_ASAP7_75t_L g17404 ( 
.A(n_17256),
.Y(n_17404)
);

INVx1_ASAP7_75t_L g17405 ( 
.A(n_17248),
.Y(n_17405)
);

NOR2xp33_ASAP7_75t_L g17406 ( 
.A(n_17217),
.B(n_3430),
.Y(n_17406)
);

NAND2xp5_ASAP7_75t_L g17407 ( 
.A(n_17302),
.B(n_3430),
.Y(n_17407)
);

AND2x2_ASAP7_75t_L g17408 ( 
.A(n_17207),
.B(n_3431),
.Y(n_17408)
);

NOR2xp67_ASAP7_75t_SL g17409 ( 
.A(n_17259),
.B(n_3431),
.Y(n_17409)
);

INVx2_ASAP7_75t_SL g17410 ( 
.A(n_17254),
.Y(n_17410)
);

CKINVDCx20_ASAP7_75t_R g17411 ( 
.A(n_17251),
.Y(n_17411)
);

NAND2xp33_ASAP7_75t_L g17412 ( 
.A(n_17274),
.B(n_3432),
.Y(n_17412)
);

NAND2xp5_ASAP7_75t_L g17413 ( 
.A(n_17221),
.B(n_3432),
.Y(n_17413)
);

NAND2x1_ASAP7_75t_SL g17414 ( 
.A(n_17252),
.B(n_3433),
.Y(n_17414)
);

INVx1_ASAP7_75t_L g17415 ( 
.A(n_17275),
.Y(n_17415)
);

NAND2xp5_ASAP7_75t_L g17416 ( 
.A(n_17244),
.B(n_3434),
.Y(n_17416)
);

NOR2xp33_ASAP7_75t_L g17417 ( 
.A(n_17281),
.B(n_3435),
.Y(n_17417)
);

INVx1_ASAP7_75t_L g17418 ( 
.A(n_17250),
.Y(n_17418)
);

INVx1_ASAP7_75t_L g17419 ( 
.A(n_17286),
.Y(n_17419)
);

A2O1A1Ixp33_ASAP7_75t_L g17420 ( 
.A1(n_17267),
.A2(n_3438),
.B(n_3436),
.C(n_3437),
.Y(n_17420)
);

OAI31xp33_ASAP7_75t_L g17421 ( 
.A1(n_17279),
.A2(n_3439),
.A3(n_3436),
.B(n_3437),
.Y(n_17421)
);

INVx1_ASAP7_75t_L g17422 ( 
.A(n_17288),
.Y(n_17422)
);

OR2x2_ASAP7_75t_L g17423 ( 
.A(n_17272),
.B(n_3440),
.Y(n_17423)
);

NAND2xp5_ASAP7_75t_L g17424 ( 
.A(n_17287),
.B(n_3441),
.Y(n_17424)
);

NAND2xp5_ASAP7_75t_SL g17425 ( 
.A(n_17258),
.B(n_3441),
.Y(n_17425)
);

INVxp67_ASAP7_75t_L g17426 ( 
.A(n_17269),
.Y(n_17426)
);

OAI221xp5_ASAP7_75t_L g17427 ( 
.A1(n_17225),
.A2(n_3444),
.B1(n_3442),
.B2(n_3443),
.C(n_3445),
.Y(n_17427)
);

NOR2xp33_ASAP7_75t_L g17428 ( 
.A(n_17271),
.B(n_3442),
.Y(n_17428)
);

OR2x2_ASAP7_75t_L g17429 ( 
.A(n_17298),
.B(n_3443),
.Y(n_17429)
);

NAND2xp5_ASAP7_75t_L g17430 ( 
.A(n_17245),
.B(n_3444),
.Y(n_17430)
);

INVxp67_ASAP7_75t_L g17431 ( 
.A(n_17228),
.Y(n_17431)
);

INVx2_ASAP7_75t_L g17432 ( 
.A(n_17243),
.Y(n_17432)
);

OAI21xp5_ASAP7_75t_SL g17433 ( 
.A1(n_17264),
.A2(n_3445),
.B(n_3446),
.Y(n_17433)
);

NAND2xp5_ASAP7_75t_L g17434 ( 
.A(n_17204),
.B(n_3446),
.Y(n_17434)
);

NAND2xp5_ASAP7_75t_L g17435 ( 
.A(n_17204),
.B(n_3447),
.Y(n_17435)
);

AND2x2_ASAP7_75t_L g17436 ( 
.A(n_17241),
.B(n_3447),
.Y(n_17436)
);

INVx1_ASAP7_75t_L g17437 ( 
.A(n_17232),
.Y(n_17437)
);

NAND2xp5_ASAP7_75t_L g17438 ( 
.A(n_17204),
.B(n_3448),
.Y(n_17438)
);

NAND2xp5_ASAP7_75t_L g17439 ( 
.A(n_17204),
.B(n_3448),
.Y(n_17439)
);

INVx1_ASAP7_75t_L g17440 ( 
.A(n_17232),
.Y(n_17440)
);

NAND2xp5_ASAP7_75t_L g17441 ( 
.A(n_17204),
.B(n_3449),
.Y(n_17441)
);

NAND4xp75_ASAP7_75t_L g17442 ( 
.A(n_17401),
.B(n_3451),
.C(n_3449),
.D(n_3450),
.Y(n_17442)
);

INVxp67_ASAP7_75t_L g17443 ( 
.A(n_17409),
.Y(n_17443)
);

NAND4xp25_ASAP7_75t_L g17444 ( 
.A(n_17421),
.B(n_3453),
.C(n_3450),
.D(n_3452),
.Y(n_17444)
);

NAND2xp5_ASAP7_75t_SL g17445 ( 
.A(n_17373),
.B(n_3452),
.Y(n_17445)
);

NAND3xp33_ASAP7_75t_SL g17446 ( 
.A(n_17370),
.B(n_3454),
.C(n_3455),
.Y(n_17446)
);

NAND2xp5_ASAP7_75t_L g17447 ( 
.A(n_17395),
.B(n_3454),
.Y(n_17447)
);

INVx1_ASAP7_75t_L g17448 ( 
.A(n_17325),
.Y(n_17448)
);

INVxp67_ASAP7_75t_SL g17449 ( 
.A(n_17387),
.Y(n_17449)
);

NAND3xp33_ASAP7_75t_L g17450 ( 
.A(n_17331),
.B(n_3455),
.C(n_3456),
.Y(n_17450)
);

NAND3xp33_ASAP7_75t_L g17451 ( 
.A(n_17390),
.B(n_3456),
.C(n_3457),
.Y(n_17451)
);

INVx2_ASAP7_75t_L g17452 ( 
.A(n_17332),
.Y(n_17452)
);

NAND3xp33_ASAP7_75t_L g17453 ( 
.A(n_17412),
.B(n_3457),
.C(n_3458),
.Y(n_17453)
);

NAND3xp33_ASAP7_75t_L g17454 ( 
.A(n_17385),
.B(n_3458),
.C(n_3459),
.Y(n_17454)
);

NOR2xp33_ASAP7_75t_L g17455 ( 
.A(n_17327),
.B(n_3459),
.Y(n_17455)
);

OAI322xp33_ASAP7_75t_L g17456 ( 
.A1(n_17323),
.A2(n_3465),
.A3(n_3464),
.B1(n_3462),
.B2(n_3460),
.C1(n_3461),
.C2(n_3463),
.Y(n_17456)
);

NAND3xp33_ASAP7_75t_SL g17457 ( 
.A(n_17411),
.B(n_3460),
.C(n_3461),
.Y(n_17457)
);

AOI21xp33_ASAP7_75t_L g17458 ( 
.A1(n_17322),
.A2(n_3462),
.B(n_3463),
.Y(n_17458)
);

NOR4xp25_ASAP7_75t_L g17459 ( 
.A(n_17437),
.B(n_17440),
.C(n_17326),
.D(n_17379),
.Y(n_17459)
);

NAND3xp33_ASAP7_75t_SL g17460 ( 
.A(n_17334),
.B(n_3464),
.C(n_3465),
.Y(n_17460)
);

NOR3xp33_ASAP7_75t_L g17461 ( 
.A(n_17399),
.B(n_17371),
.C(n_17398),
.Y(n_17461)
);

NOR2xp33_ASAP7_75t_L g17462 ( 
.A(n_17335),
.B(n_3466),
.Y(n_17462)
);

NAND4xp25_ASAP7_75t_SL g17463 ( 
.A(n_17355),
.B(n_3468),
.C(n_3466),
.D(n_3467),
.Y(n_17463)
);

NAND2xp5_ASAP7_75t_L g17464 ( 
.A(n_17341),
.B(n_3467),
.Y(n_17464)
);

NOR3xp33_ASAP7_75t_SL g17465 ( 
.A(n_17359),
.B(n_3468),
.C(n_3469),
.Y(n_17465)
);

NAND4xp25_ASAP7_75t_L g17466 ( 
.A(n_17375),
.B(n_3471),
.C(n_3469),
.D(n_3470),
.Y(n_17466)
);

NOR2x1_ASAP7_75t_SL g17467 ( 
.A(n_17377),
.B(n_3470),
.Y(n_17467)
);

O2A1O1Ixp5_ASAP7_75t_L g17468 ( 
.A1(n_17333),
.A2(n_3473),
.B(n_3471),
.C(n_3472),
.Y(n_17468)
);

NAND2xp5_ASAP7_75t_L g17469 ( 
.A(n_17340),
.B(n_3473),
.Y(n_17469)
);

NOR4xp25_ASAP7_75t_L g17470 ( 
.A(n_17346),
.B(n_3477),
.C(n_3475),
.D(n_3476),
.Y(n_17470)
);

NAND3xp33_ASAP7_75t_L g17471 ( 
.A(n_17372),
.B(n_3476),
.C(n_3477),
.Y(n_17471)
);

NAND2xp5_ASAP7_75t_SL g17472 ( 
.A(n_17357),
.B(n_3478),
.Y(n_17472)
);

NOR2xp67_ASAP7_75t_L g17473 ( 
.A(n_17427),
.B(n_3478),
.Y(n_17473)
);

NOR4xp25_ASAP7_75t_L g17474 ( 
.A(n_17431),
.B(n_3481),
.C(n_3479),
.D(n_3480),
.Y(n_17474)
);

NOR2x1_ASAP7_75t_L g17475 ( 
.A(n_17423),
.B(n_3479),
.Y(n_17475)
);

OAI211xp5_ASAP7_75t_L g17476 ( 
.A1(n_17337),
.A2(n_3483),
.B(n_3481),
.C(n_3482),
.Y(n_17476)
);

NAND3xp33_ASAP7_75t_SL g17477 ( 
.A(n_17396),
.B(n_3482),
.C(n_3483),
.Y(n_17477)
);

NAND3xp33_ASAP7_75t_L g17478 ( 
.A(n_17336),
.B(n_3484),
.C(n_3485),
.Y(n_17478)
);

OAI211xp5_ASAP7_75t_L g17479 ( 
.A1(n_17430),
.A2(n_3486),
.B(n_3487),
.C(n_3485),
.Y(n_17479)
);

NOR2xp33_ASAP7_75t_L g17480 ( 
.A(n_17434),
.B(n_4311),
.Y(n_17480)
);

OR2x2_ASAP7_75t_L g17481 ( 
.A(n_17429),
.B(n_3484),
.Y(n_17481)
);

NOR2xp33_ASAP7_75t_L g17482 ( 
.A(n_17435),
.B(n_4312),
.Y(n_17482)
);

O2A1O1Ixp33_ASAP7_75t_L g17483 ( 
.A1(n_17324),
.A2(n_3489),
.B(n_3486),
.C(n_3488),
.Y(n_17483)
);

NAND3xp33_ASAP7_75t_SL g17484 ( 
.A(n_17348),
.B(n_3489),
.C(n_3490),
.Y(n_17484)
);

OAI21xp33_ASAP7_75t_L g17485 ( 
.A1(n_17405),
.A2(n_17432),
.B(n_17362),
.Y(n_17485)
);

OA22x2_ASAP7_75t_L g17486 ( 
.A1(n_17433),
.A2(n_3493),
.B1(n_3491),
.B2(n_3492),
.Y(n_17486)
);

AND4x1_ASAP7_75t_L g17487 ( 
.A(n_17378),
.B(n_3493),
.C(n_3491),
.D(n_3492),
.Y(n_17487)
);

NOR3xp33_ASAP7_75t_SL g17488 ( 
.A(n_17328),
.B(n_3494),
.C(n_3495),
.Y(n_17488)
);

NAND4xp25_ASAP7_75t_L g17489 ( 
.A(n_17374),
.B(n_3497),
.C(n_3494),
.D(n_3496),
.Y(n_17489)
);

NAND2xp5_ASAP7_75t_L g17490 ( 
.A(n_17320),
.B(n_3498),
.Y(n_17490)
);

NOR4xp25_ASAP7_75t_L g17491 ( 
.A(n_17426),
.B(n_4322),
.C(n_3500),
.D(n_3496),
.Y(n_17491)
);

NAND2xp5_ASAP7_75t_SL g17492 ( 
.A(n_17342),
.B(n_3499),
.Y(n_17492)
);

NOR3x1_ASAP7_75t_L g17493 ( 
.A(n_17383),
.B(n_3499),
.C(n_3500),
.Y(n_17493)
);

NOR4xp25_ASAP7_75t_L g17494 ( 
.A(n_17382),
.B(n_4317),
.C(n_4310),
.D(n_3503),
.Y(n_17494)
);

INVx1_ASAP7_75t_SL g17495 ( 
.A(n_17361),
.Y(n_17495)
);

NAND4xp25_ASAP7_75t_L g17496 ( 
.A(n_17356),
.B(n_3504),
.C(n_3501),
.D(n_3502),
.Y(n_17496)
);

AOI22xp33_ASAP7_75t_L g17497 ( 
.A1(n_17410),
.A2(n_3505),
.B1(n_3501),
.B2(n_3504),
.Y(n_17497)
);

NAND4xp25_ASAP7_75t_L g17498 ( 
.A(n_17428),
.B(n_3507),
.C(n_3505),
.D(n_3506),
.Y(n_17498)
);

XOR2x2_ASAP7_75t_L g17499 ( 
.A(n_17380),
.B(n_3506),
.Y(n_17499)
);

AOI211x1_ASAP7_75t_L g17500 ( 
.A1(n_17321),
.A2(n_3509),
.B(n_3507),
.C(n_3508),
.Y(n_17500)
);

O2A1O1Ixp33_ASAP7_75t_L g17501 ( 
.A1(n_17330),
.A2(n_3512),
.B(n_3510),
.C(n_3511),
.Y(n_17501)
);

NAND3xp33_ASAP7_75t_L g17502 ( 
.A(n_17368),
.B(n_17343),
.C(n_17350),
.Y(n_17502)
);

NOR2x1_ASAP7_75t_L g17503 ( 
.A(n_17438),
.B(n_3511),
.Y(n_17503)
);

NOR3xp33_ASAP7_75t_SL g17504 ( 
.A(n_17384),
.B(n_3510),
.C(n_3512),
.Y(n_17504)
);

NOR3xp33_ASAP7_75t_L g17505 ( 
.A(n_17415),
.B(n_3513),
.C(n_3514),
.Y(n_17505)
);

NOR2x1_ASAP7_75t_L g17506 ( 
.A(n_17439),
.B(n_3514),
.Y(n_17506)
);

OAI22xp5_ASAP7_75t_L g17507 ( 
.A1(n_17441),
.A2(n_4324),
.B1(n_3516),
.B2(n_3513),
.Y(n_17507)
);

NAND2xp5_ASAP7_75t_L g17508 ( 
.A(n_17367),
.B(n_3516),
.Y(n_17508)
);

AOI21xp5_ASAP7_75t_SL g17509 ( 
.A1(n_17420),
.A2(n_3518),
.B(n_3517),
.Y(n_17509)
);

XNOR2xp5_ASAP7_75t_L g17510 ( 
.A(n_17353),
.B(n_3515),
.Y(n_17510)
);

NOR3xp33_ASAP7_75t_L g17511 ( 
.A(n_17381),
.B(n_3515),
.C(n_3517),
.Y(n_17511)
);

NOR2x1_ASAP7_75t_L g17512 ( 
.A(n_17402),
.B(n_3519),
.Y(n_17512)
);

NAND4xp25_ASAP7_75t_L g17513 ( 
.A(n_17351),
.B(n_3520),
.C(n_3518),
.D(n_3519),
.Y(n_17513)
);

NAND2xp5_ASAP7_75t_L g17514 ( 
.A(n_17338),
.B(n_3521),
.Y(n_17514)
);

NAND3xp33_ASAP7_75t_SL g17515 ( 
.A(n_17360),
.B(n_3520),
.C(n_3522),
.Y(n_17515)
);

NAND2xp5_ASAP7_75t_SL g17516 ( 
.A(n_17369),
.B(n_3522),
.Y(n_17516)
);

NOR3x1_ASAP7_75t_SL g17517 ( 
.A(n_17376),
.B(n_3523),
.C(n_3524),
.Y(n_17517)
);

NOR2xp33_ASAP7_75t_SL g17518 ( 
.A(n_17406),
.B(n_3523),
.Y(n_17518)
);

AOI211xp5_ASAP7_75t_L g17519 ( 
.A1(n_17345),
.A2(n_3526),
.B(n_3524),
.C(n_3525),
.Y(n_17519)
);

NAND2xp5_ASAP7_75t_L g17520 ( 
.A(n_17414),
.B(n_3527),
.Y(n_17520)
);

AOI221x1_ASAP7_75t_L g17521 ( 
.A1(n_17391),
.A2(n_3528),
.B1(n_3525),
.B2(n_3527),
.C(n_3529),
.Y(n_17521)
);

NAND2xp5_ASAP7_75t_L g17522 ( 
.A(n_17352),
.B(n_3529),
.Y(n_17522)
);

NOR3xp33_ASAP7_75t_L g17523 ( 
.A(n_17347),
.B(n_3528),
.C(n_3531),
.Y(n_17523)
);

NAND2xp5_ASAP7_75t_SL g17524 ( 
.A(n_17400),
.B(n_3531),
.Y(n_17524)
);

NAND2xp5_ASAP7_75t_L g17525 ( 
.A(n_17329),
.B(n_3533),
.Y(n_17525)
);

NOR2xp67_ASAP7_75t_L g17526 ( 
.A(n_17394),
.B(n_3533),
.Y(n_17526)
);

AND4x1_ASAP7_75t_L g17527 ( 
.A(n_17344),
.B(n_3535),
.C(n_3532),
.D(n_3534),
.Y(n_17527)
);

OAI211xp5_ASAP7_75t_L g17528 ( 
.A1(n_17389),
.A2(n_3536),
.B(n_3537),
.C(n_3535),
.Y(n_17528)
);

NAND2xp5_ASAP7_75t_L g17529 ( 
.A(n_17407),
.B(n_17365),
.Y(n_17529)
);

AOI21xp5_ASAP7_75t_L g17530 ( 
.A1(n_17349),
.A2(n_3532),
.B(n_3536),
.Y(n_17530)
);

NAND2xp5_ASAP7_75t_L g17531 ( 
.A(n_17354),
.B(n_3538),
.Y(n_17531)
);

AOI21xp5_ASAP7_75t_L g17532 ( 
.A1(n_17392),
.A2(n_3537),
.B(n_3538),
.Y(n_17532)
);

NOR3xp33_ASAP7_75t_L g17533 ( 
.A(n_17393),
.B(n_3539),
.C(n_3540),
.Y(n_17533)
);

AOI211xp5_ASAP7_75t_L g17534 ( 
.A1(n_17425),
.A2(n_3541),
.B(n_3539),
.C(n_3540),
.Y(n_17534)
);

INVx1_ASAP7_75t_L g17535 ( 
.A(n_17403),
.Y(n_17535)
);

A2O1A1Ixp33_ASAP7_75t_L g17536 ( 
.A1(n_17404),
.A2(n_17386),
.B(n_17416),
.C(n_17413),
.Y(n_17536)
);

NAND4xp25_ASAP7_75t_SL g17537 ( 
.A(n_17424),
.B(n_3543),
.C(n_3541),
.D(n_3542),
.Y(n_17537)
);

NOR3xp33_ASAP7_75t_L g17538 ( 
.A(n_17418),
.B(n_3542),
.C(n_3543),
.Y(n_17538)
);

NOR2xp33_ASAP7_75t_L g17539 ( 
.A(n_17366),
.B(n_4319),
.Y(n_17539)
);

NAND4xp75_ASAP7_75t_L g17540 ( 
.A(n_17419),
.B(n_3546),
.C(n_3544),
.D(n_3545),
.Y(n_17540)
);

OAI21xp33_ASAP7_75t_L g17541 ( 
.A1(n_17363),
.A2(n_3546),
.B(n_3547),
.Y(n_17541)
);

NAND4xp25_ASAP7_75t_L g17542 ( 
.A(n_17358),
.B(n_3549),
.C(n_3547),
.D(n_3548),
.Y(n_17542)
);

AOI22xp5_ASAP7_75t_L g17543 ( 
.A1(n_17422),
.A2(n_17339),
.B1(n_17364),
.B2(n_17388),
.Y(n_17543)
);

NOR4xp25_ASAP7_75t_L g17544 ( 
.A(n_17417),
.B(n_4316),
.C(n_4309),
.D(n_3551),
.Y(n_17544)
);

INVx1_ASAP7_75t_L g17545 ( 
.A(n_17436),
.Y(n_17545)
);

NOR2x1_ASAP7_75t_L g17546 ( 
.A(n_17397),
.B(n_3550),
.Y(n_17546)
);

NOR2x1_ASAP7_75t_L g17547 ( 
.A(n_17408),
.B(n_3550),
.Y(n_17547)
);

AOI33xp33_ASAP7_75t_L g17548 ( 
.A1(n_17323),
.A2(n_3552),
.A3(n_3554),
.B1(n_3548),
.B2(n_3551),
.B3(n_3553),
.Y(n_17548)
);

AOI222xp33_ASAP7_75t_L g17549 ( 
.A1(n_17323),
.A2(n_3554),
.B1(n_3556),
.B2(n_3552),
.C1(n_3553),
.C2(n_3555),
.Y(n_17549)
);

NAND2xp5_ASAP7_75t_L g17550 ( 
.A(n_17395),
.B(n_3556),
.Y(n_17550)
);

NAND3xp33_ASAP7_75t_L g17551 ( 
.A(n_17331),
.B(n_3555),
.C(n_3557),
.Y(n_17551)
);

NAND3xp33_ASAP7_75t_SL g17552 ( 
.A(n_17370),
.B(n_3557),
.C(n_3558),
.Y(n_17552)
);

NOR2xp33_ASAP7_75t_R g17553 ( 
.A(n_17359),
.B(n_3558),
.Y(n_17553)
);

OAI21xp5_ASAP7_75t_L g17554 ( 
.A1(n_17355),
.A2(n_3559),
.B(n_3560),
.Y(n_17554)
);

AOI211xp5_ASAP7_75t_L g17555 ( 
.A1(n_17370),
.A2(n_3562),
.B(n_3559),
.C(n_3561),
.Y(n_17555)
);

NOR3xp33_ASAP7_75t_L g17556 ( 
.A(n_17401),
.B(n_3561),
.C(n_3562),
.Y(n_17556)
);

AOI211xp5_ASAP7_75t_L g17557 ( 
.A1(n_17370),
.A2(n_3565),
.B(n_3563),
.C(n_3564),
.Y(n_17557)
);

NAND3xp33_ASAP7_75t_L g17558 ( 
.A(n_17331),
.B(n_3563),
.C(n_3565),
.Y(n_17558)
);

INVx1_ASAP7_75t_L g17559 ( 
.A(n_17325),
.Y(n_17559)
);

NOR2x1_ASAP7_75t_L g17560 ( 
.A(n_17325),
.B(n_3567),
.Y(n_17560)
);

NOR2x1_ASAP7_75t_L g17561 ( 
.A(n_17325),
.B(n_3568),
.Y(n_17561)
);

NOR3x1_ASAP7_75t_L g17562 ( 
.A(n_17370),
.B(n_3566),
.C(n_3568),
.Y(n_17562)
);

NOR3xp33_ASAP7_75t_SL g17563 ( 
.A(n_17401),
.B(n_3569),
.C(n_3570),
.Y(n_17563)
);

NOR2x1_ASAP7_75t_L g17564 ( 
.A(n_17325),
.B(n_3571),
.Y(n_17564)
);

AOI22xp5_ASAP7_75t_L g17565 ( 
.A1(n_17411),
.A2(n_3572),
.B1(n_3569),
.B2(n_3571),
.Y(n_17565)
);

O2A1O1Ixp33_ASAP7_75t_L g17566 ( 
.A1(n_17401),
.A2(n_3576),
.B(n_3573),
.C(n_3574),
.Y(n_17566)
);

AOI22xp5_ASAP7_75t_L g17567 ( 
.A1(n_17411),
.A2(n_3578),
.B1(n_3576),
.B2(n_3577),
.Y(n_17567)
);

INVx1_ASAP7_75t_L g17568 ( 
.A(n_17325),
.Y(n_17568)
);

BUFx3_ASAP7_75t_L g17569 ( 
.A(n_17398),
.Y(n_17569)
);

NAND4xp25_ASAP7_75t_SL g17570 ( 
.A(n_17373),
.B(n_3579),
.C(n_3577),
.D(n_3578),
.Y(n_17570)
);

NAND4xp25_ASAP7_75t_L g17571 ( 
.A(n_17401),
.B(n_3581),
.C(n_3579),
.D(n_3580),
.Y(n_17571)
);

NOR3xp33_ASAP7_75t_L g17572 ( 
.A(n_17401),
.B(n_3580),
.C(n_3581),
.Y(n_17572)
);

NAND3xp33_ASAP7_75t_L g17573 ( 
.A(n_17331),
.B(n_3582),
.C(n_3583),
.Y(n_17573)
);

NAND2xp5_ASAP7_75t_L g17574 ( 
.A(n_17395),
.B(n_3583),
.Y(n_17574)
);

INVx1_ASAP7_75t_L g17575 ( 
.A(n_17325),
.Y(n_17575)
);

NOR3xp33_ASAP7_75t_SL g17576 ( 
.A(n_17401),
.B(n_3582),
.C(n_3584),
.Y(n_17576)
);

AOI21xp5_ASAP7_75t_L g17577 ( 
.A1(n_17401),
.A2(n_3584),
.B(n_3585),
.Y(n_17577)
);

AOI221xp5_ASAP7_75t_L g17578 ( 
.A1(n_17427),
.A2(n_3587),
.B1(n_3585),
.B2(n_3586),
.C(n_3588),
.Y(n_17578)
);

NOR4xp25_ASAP7_75t_L g17579 ( 
.A(n_17401),
.B(n_4323),
.C(n_4314),
.D(n_3588),
.Y(n_17579)
);

NAND4xp25_ASAP7_75t_L g17580 ( 
.A(n_17401),
.B(n_3589),
.C(n_3586),
.D(n_3587),
.Y(n_17580)
);

NAND4xp25_ASAP7_75t_L g17581 ( 
.A(n_17401),
.B(n_3591),
.C(n_3589),
.D(n_3590),
.Y(n_17581)
);

NOR2x1_ASAP7_75t_L g17582 ( 
.A(n_17325),
.B(n_3592),
.Y(n_17582)
);

NOR2xp67_ASAP7_75t_SL g17583 ( 
.A(n_17398),
.B(n_3591),
.Y(n_17583)
);

O2A1O1Ixp33_ASAP7_75t_L g17584 ( 
.A1(n_17401),
.A2(n_3594),
.B(n_3592),
.C(n_3593),
.Y(n_17584)
);

NAND2xp5_ASAP7_75t_L g17585 ( 
.A(n_17395),
.B(n_3594),
.Y(n_17585)
);

NAND4xp25_ASAP7_75t_L g17586 ( 
.A(n_17401),
.B(n_3596),
.C(n_3593),
.D(n_3595),
.Y(n_17586)
);

NAND4xp25_ASAP7_75t_L g17587 ( 
.A(n_17401),
.B(n_3597),
.C(n_3595),
.D(n_3596),
.Y(n_17587)
);

INVxp33_ASAP7_75t_SL g17588 ( 
.A(n_17330),
.Y(n_17588)
);

AOI21xp5_ASAP7_75t_L g17589 ( 
.A1(n_17401),
.A2(n_3598),
.B(n_3599),
.Y(n_17589)
);

OAI21xp33_ASAP7_75t_L g17590 ( 
.A1(n_17401),
.A2(n_3600),
.B(n_3601),
.Y(n_17590)
);

NOR2x1_ASAP7_75t_L g17591 ( 
.A(n_17325),
.B(n_3601),
.Y(n_17591)
);

NAND3xp33_ASAP7_75t_SL g17592 ( 
.A(n_17370),
.B(n_3600),
.C(n_3602),
.Y(n_17592)
);

OA211x2_ASAP7_75t_L g17593 ( 
.A1(n_17341),
.A2(n_3604),
.B(n_3602),
.C(n_3603),
.Y(n_17593)
);

INVx1_ASAP7_75t_L g17594 ( 
.A(n_17325),
.Y(n_17594)
);

OAI221xp5_ASAP7_75t_L g17595 ( 
.A1(n_17421),
.A2(n_3605),
.B1(n_3603),
.B2(n_3604),
.C(n_3606),
.Y(n_17595)
);

NAND3xp33_ASAP7_75t_SL g17596 ( 
.A(n_17370),
.B(n_3605),
.C(n_3606),
.Y(n_17596)
);

NAND4xp75_ASAP7_75t_L g17597 ( 
.A(n_17401),
.B(n_3609),
.C(n_3607),
.D(n_3608),
.Y(n_17597)
);

NOR2xp33_ASAP7_75t_SL g17598 ( 
.A(n_17361),
.B(n_3607),
.Y(n_17598)
);

O2A1O1Ixp33_ASAP7_75t_L g17599 ( 
.A1(n_17401),
.A2(n_3611),
.B(n_3608),
.C(n_3610),
.Y(n_17599)
);

AOI22xp5_ASAP7_75t_L g17600 ( 
.A1(n_17588),
.A2(n_3613),
.B1(n_3610),
.B2(n_3612),
.Y(n_17600)
);

AOI31xp33_ASAP7_75t_L g17601 ( 
.A1(n_17481),
.A2(n_3614),
.A3(n_3612),
.B(n_3613),
.Y(n_17601)
);

AOI22xp5_ASAP7_75t_L g17602 ( 
.A1(n_17461),
.A2(n_3616),
.B1(n_3614),
.B2(n_3615),
.Y(n_17602)
);

INVx1_ASAP7_75t_L g17603 ( 
.A(n_17517),
.Y(n_17603)
);

INVx1_ASAP7_75t_L g17604 ( 
.A(n_17447),
.Y(n_17604)
);

AOI22xp5_ASAP7_75t_L g17605 ( 
.A1(n_17539),
.A2(n_3618),
.B1(n_3616),
.B2(n_3617),
.Y(n_17605)
);

NOR2x1_ASAP7_75t_L g17606 ( 
.A(n_17560),
.B(n_4314),
.Y(n_17606)
);

AOI22xp5_ASAP7_75t_L g17607 ( 
.A1(n_17598),
.A2(n_3619),
.B1(n_3617),
.B2(n_3618),
.Y(n_17607)
);

AOI22xp5_ASAP7_75t_L g17608 ( 
.A1(n_17485),
.A2(n_3622),
.B1(n_3620),
.B2(n_3621),
.Y(n_17608)
);

NOR4xp25_ASAP7_75t_L g17609 ( 
.A(n_17536),
.B(n_3622),
.C(n_3620),
.D(n_3621),
.Y(n_17609)
);

INVx2_ASAP7_75t_L g17610 ( 
.A(n_17540),
.Y(n_17610)
);

O2A1O1Ixp33_ASAP7_75t_L g17611 ( 
.A1(n_17472),
.A2(n_3631),
.B(n_3639),
.C(n_3623),
.Y(n_17611)
);

AOI22xp5_ASAP7_75t_L g17612 ( 
.A1(n_17556),
.A2(n_17572),
.B1(n_17537),
.B2(n_17518),
.Y(n_17612)
);

AO22x2_ASAP7_75t_L g17613 ( 
.A1(n_17448),
.A2(n_3625),
.B1(n_3623),
.B2(n_3624),
.Y(n_17613)
);

INVx1_ASAP7_75t_L g17614 ( 
.A(n_17550),
.Y(n_17614)
);

AOI22xp5_ASAP7_75t_L g17615 ( 
.A1(n_17457),
.A2(n_3626),
.B1(n_3624),
.B2(n_3625),
.Y(n_17615)
);

OA22x2_ASAP7_75t_L g17616 ( 
.A1(n_17510),
.A2(n_3628),
.B1(n_3626),
.B2(n_3627),
.Y(n_17616)
);

INVx1_ASAP7_75t_L g17617 ( 
.A(n_17574),
.Y(n_17617)
);

A2O1A1Ixp33_ASAP7_75t_L g17618 ( 
.A1(n_17566),
.A2(n_3629),
.B(n_3627),
.C(n_3628),
.Y(n_17618)
);

INVxp67_ASAP7_75t_L g17619 ( 
.A(n_17583),
.Y(n_17619)
);

AOI22xp5_ASAP7_75t_L g17620 ( 
.A1(n_17570),
.A2(n_3631),
.B1(n_3629),
.B2(n_3630),
.Y(n_17620)
);

AOI22xp33_ASAP7_75t_L g17621 ( 
.A1(n_17569),
.A2(n_3633),
.B1(n_3630),
.B2(n_3632),
.Y(n_17621)
);

NAND2xp5_ASAP7_75t_L g17622 ( 
.A(n_17579),
.B(n_3632),
.Y(n_17622)
);

AOI221xp5_ASAP7_75t_L g17623 ( 
.A1(n_17459),
.A2(n_3635),
.B1(n_3633),
.B2(n_3634),
.C(n_3636),
.Y(n_17623)
);

NAND2xp5_ASAP7_75t_L g17624 ( 
.A(n_17455),
.B(n_3634),
.Y(n_17624)
);

AO22x2_ASAP7_75t_L g17625 ( 
.A1(n_17559),
.A2(n_3637),
.B1(n_3635),
.B2(n_3636),
.Y(n_17625)
);

OAI22xp5_ASAP7_75t_L g17626 ( 
.A1(n_17478),
.A2(n_3641),
.B1(n_3638),
.B2(n_3639),
.Y(n_17626)
);

AOI22xp5_ASAP7_75t_L g17627 ( 
.A1(n_17463),
.A2(n_3642),
.B1(n_3638),
.B2(n_3641),
.Y(n_17627)
);

INVxp67_ASAP7_75t_SL g17628 ( 
.A(n_17561),
.Y(n_17628)
);

INVx1_ASAP7_75t_L g17629 ( 
.A(n_17585),
.Y(n_17629)
);

AOI22xp5_ASAP7_75t_L g17630 ( 
.A1(n_17460),
.A2(n_3644),
.B1(n_3642),
.B2(n_3643),
.Y(n_17630)
);

AO22x2_ASAP7_75t_L g17631 ( 
.A1(n_17568),
.A2(n_3645),
.B1(n_3643),
.B2(n_3644),
.Y(n_17631)
);

AOI221xp5_ASAP7_75t_L g17632 ( 
.A1(n_17595),
.A2(n_3648),
.B1(n_3646),
.B2(n_3647),
.C(n_3649),
.Y(n_17632)
);

AOI22xp5_ASAP7_75t_L g17633 ( 
.A1(n_17477),
.A2(n_3648),
.B1(n_3646),
.B2(n_3647),
.Y(n_17633)
);

INVxp67_ASAP7_75t_SL g17634 ( 
.A(n_17564),
.Y(n_17634)
);

NAND2xp5_ASAP7_75t_L g17635 ( 
.A(n_17462),
.B(n_3649),
.Y(n_17635)
);

AOI22xp5_ASAP7_75t_L g17636 ( 
.A1(n_17515),
.A2(n_3652),
.B1(n_3650),
.B2(n_3651),
.Y(n_17636)
);

INVx2_ASAP7_75t_L g17637 ( 
.A(n_17442),
.Y(n_17637)
);

AOI22xp5_ASAP7_75t_L g17638 ( 
.A1(n_17498),
.A2(n_3653),
.B1(n_3650),
.B2(n_3652),
.Y(n_17638)
);

AOI31xp33_ASAP7_75t_L g17639 ( 
.A1(n_17443),
.A2(n_3655),
.A3(n_3653),
.B(n_3654),
.Y(n_17639)
);

NOR2xp33_ASAP7_75t_L g17640 ( 
.A(n_17444),
.B(n_3654),
.Y(n_17640)
);

AOI221xp5_ASAP7_75t_L g17641 ( 
.A1(n_17500),
.A2(n_3657),
.B1(n_3655),
.B2(n_3656),
.C(n_3658),
.Y(n_17641)
);

AOI22xp5_ASAP7_75t_L g17642 ( 
.A1(n_17593),
.A2(n_3658),
.B1(n_3656),
.B2(n_3657),
.Y(n_17642)
);

OAI22x1_ASAP7_75t_L g17643 ( 
.A1(n_17471),
.A2(n_3661),
.B1(n_3659),
.B2(n_3660),
.Y(n_17643)
);

NOR2xp33_ASAP7_75t_L g17644 ( 
.A(n_17466),
.B(n_3659),
.Y(n_17644)
);

INVxp67_ASAP7_75t_SL g17645 ( 
.A(n_17582),
.Y(n_17645)
);

NOR2x1_ASAP7_75t_L g17646 ( 
.A(n_17591),
.B(n_4310),
.Y(n_17646)
);

INVxp67_ASAP7_75t_L g17647 ( 
.A(n_17480),
.Y(n_17647)
);

NOR2x1_ASAP7_75t_L g17648 ( 
.A(n_17575),
.B(n_4311),
.Y(n_17648)
);

OAI22xp5_ASAP7_75t_L g17649 ( 
.A1(n_17490),
.A2(n_3664),
.B1(n_3662),
.B2(n_3663),
.Y(n_17649)
);

NOR4xp25_ASAP7_75t_L g17650 ( 
.A(n_17464),
.B(n_3664),
.C(n_3662),
.D(n_3663),
.Y(n_17650)
);

INVxp67_ASAP7_75t_SL g17651 ( 
.A(n_17547),
.Y(n_17651)
);

NOR4xp25_ASAP7_75t_L g17652 ( 
.A(n_17495),
.B(n_3667),
.C(n_3665),
.D(n_3666),
.Y(n_17652)
);

INVx1_ASAP7_75t_L g17653 ( 
.A(n_17546),
.Y(n_17653)
);

OAI22xp5_ASAP7_75t_L g17654 ( 
.A1(n_17469),
.A2(n_3670),
.B1(n_3668),
.B2(n_3669),
.Y(n_17654)
);

NOR2xp33_ASAP7_75t_L g17655 ( 
.A(n_17479),
.B(n_3669),
.Y(n_17655)
);

NOR2x1_ASAP7_75t_L g17656 ( 
.A(n_17594),
.B(n_4321),
.Y(n_17656)
);

INVx1_ASAP7_75t_L g17657 ( 
.A(n_17512),
.Y(n_17657)
);

XNOR2x1_ASAP7_75t_L g17658 ( 
.A(n_17499),
.B(n_17503),
.Y(n_17658)
);

INVx1_ASAP7_75t_L g17659 ( 
.A(n_17506),
.Y(n_17659)
);

INVx1_ASAP7_75t_L g17660 ( 
.A(n_17486),
.Y(n_17660)
);

INVx1_ASAP7_75t_L g17661 ( 
.A(n_17520),
.Y(n_17661)
);

NOR2x1_ASAP7_75t_L g17662 ( 
.A(n_17597),
.B(n_4321),
.Y(n_17662)
);

NAND2xp5_ASAP7_75t_L g17663 ( 
.A(n_17482),
.B(n_3670),
.Y(n_17663)
);

AOI22xp5_ASAP7_75t_L g17664 ( 
.A1(n_17484),
.A2(n_3673),
.B1(n_3671),
.B2(n_3672),
.Y(n_17664)
);

NAND2xp5_ASAP7_75t_SL g17665 ( 
.A(n_17474),
.B(n_3671),
.Y(n_17665)
);

INVx2_ASAP7_75t_L g17666 ( 
.A(n_17562),
.Y(n_17666)
);

INVx1_ASAP7_75t_L g17667 ( 
.A(n_17508),
.Y(n_17667)
);

NOR2xp33_ASAP7_75t_L g17668 ( 
.A(n_17489),
.B(n_3673),
.Y(n_17668)
);

AOI22xp5_ASAP7_75t_L g17669 ( 
.A1(n_17446),
.A2(n_3677),
.B1(n_3675),
.B2(n_3676),
.Y(n_17669)
);

INVx1_ASAP7_75t_L g17670 ( 
.A(n_17475),
.Y(n_17670)
);

AOI221xp5_ASAP7_75t_L g17671 ( 
.A1(n_17552),
.A2(n_3679),
.B1(n_3676),
.B2(n_3678),
.C(n_3680),
.Y(n_17671)
);

AOI22xp5_ASAP7_75t_L g17672 ( 
.A1(n_17592),
.A2(n_3681),
.B1(n_3678),
.B2(n_3680),
.Y(n_17672)
);

NOR2xp33_ASAP7_75t_L g17673 ( 
.A(n_17596),
.B(n_3681),
.Y(n_17673)
);

OR2x2_ASAP7_75t_L g17674 ( 
.A(n_17544),
.B(n_3684),
.Y(n_17674)
);

INVx1_ASAP7_75t_L g17675 ( 
.A(n_17467),
.Y(n_17675)
);

NOR2x1_ASAP7_75t_L g17676 ( 
.A(n_17453),
.B(n_4315),
.Y(n_17676)
);

INVx1_ASAP7_75t_L g17677 ( 
.A(n_17488),
.Y(n_17677)
);

INVx1_ASAP7_75t_L g17678 ( 
.A(n_17531),
.Y(n_17678)
);

INVxp67_ASAP7_75t_L g17679 ( 
.A(n_17525),
.Y(n_17679)
);

AO22x2_ASAP7_75t_L g17680 ( 
.A1(n_17545),
.A2(n_3685),
.B1(n_3683),
.B2(n_3684),
.Y(n_17680)
);

AOI22xp5_ASAP7_75t_L g17681 ( 
.A1(n_17473),
.A2(n_3687),
.B1(n_3683),
.B2(n_3686),
.Y(n_17681)
);

OAI22xp5_ASAP7_75t_L g17682 ( 
.A1(n_17451),
.A2(n_3690),
.B1(n_3688),
.B2(n_3689),
.Y(n_17682)
);

AOI22xp5_ASAP7_75t_L g17683 ( 
.A1(n_17533),
.A2(n_3690),
.B1(n_3688),
.B2(n_3689),
.Y(n_17683)
);

AOI22xp5_ASAP7_75t_L g17684 ( 
.A1(n_17578),
.A2(n_3693),
.B1(n_3691),
.B2(n_3692),
.Y(n_17684)
);

INVx1_ASAP7_75t_L g17685 ( 
.A(n_17514),
.Y(n_17685)
);

INVx1_ASAP7_75t_L g17686 ( 
.A(n_17522),
.Y(n_17686)
);

NAND2xp5_ASAP7_75t_L g17687 ( 
.A(n_17511),
.B(n_17590),
.Y(n_17687)
);

INVx1_ASAP7_75t_L g17688 ( 
.A(n_17563),
.Y(n_17688)
);

A2O1A1Ixp33_ASAP7_75t_SL g17689 ( 
.A1(n_17543),
.A2(n_3693),
.B(n_3691),
.C(n_3692),
.Y(n_17689)
);

OAI22xp5_ASAP7_75t_SL g17690 ( 
.A1(n_17449),
.A2(n_3696),
.B1(n_3694),
.B2(n_3695),
.Y(n_17690)
);

AO22x2_ASAP7_75t_L g17691 ( 
.A1(n_17452),
.A2(n_3697),
.B1(n_3695),
.B2(n_3696),
.Y(n_17691)
);

NOR2x1_ASAP7_75t_L g17692 ( 
.A(n_17571),
.B(n_4313),
.Y(n_17692)
);

INVx1_ASAP7_75t_L g17693 ( 
.A(n_17576),
.Y(n_17693)
);

NOR4xp25_ASAP7_75t_L g17694 ( 
.A(n_17502),
.B(n_3699),
.C(n_3697),
.D(n_3698),
.Y(n_17694)
);

AOI22xp5_ASAP7_75t_L g17695 ( 
.A1(n_17476),
.A2(n_3701),
.B1(n_3699),
.B2(n_3700),
.Y(n_17695)
);

NOR2xp33_ASAP7_75t_L g17696 ( 
.A(n_17450),
.B(n_3701),
.Y(n_17696)
);

NAND2xp5_ASAP7_75t_L g17697 ( 
.A(n_17555),
.B(n_3702),
.Y(n_17697)
);

NOR2x1_ASAP7_75t_L g17698 ( 
.A(n_17580),
.B(n_17581),
.Y(n_17698)
);

INVx1_ASAP7_75t_L g17699 ( 
.A(n_17454),
.Y(n_17699)
);

INVx1_ASAP7_75t_L g17700 ( 
.A(n_17468),
.Y(n_17700)
);

INVx1_ASAP7_75t_L g17701 ( 
.A(n_17493),
.Y(n_17701)
);

AOI22xp5_ASAP7_75t_L g17702 ( 
.A1(n_17551),
.A2(n_3704),
.B1(n_3702),
.B2(n_3703),
.Y(n_17702)
);

INVx1_ASAP7_75t_L g17703 ( 
.A(n_17558),
.Y(n_17703)
);

INVx2_ASAP7_75t_L g17704 ( 
.A(n_17565),
.Y(n_17704)
);

INVx1_ASAP7_75t_L g17705 ( 
.A(n_17573),
.Y(n_17705)
);

AOI22xp5_ASAP7_75t_L g17706 ( 
.A1(n_17492),
.A2(n_3707),
.B1(n_3705),
.B2(n_3706),
.Y(n_17706)
);

AO22x2_ASAP7_75t_L g17707 ( 
.A1(n_17535),
.A2(n_3707),
.B1(n_3705),
.B2(n_3706),
.Y(n_17707)
);

NOR4xp25_ASAP7_75t_L g17708 ( 
.A(n_17524),
.B(n_3710),
.C(n_3708),
.D(n_3709),
.Y(n_17708)
);

AOI22xp5_ASAP7_75t_L g17709 ( 
.A1(n_17516),
.A2(n_3711),
.B1(n_3709),
.B2(n_3710),
.Y(n_17709)
);

NAND2xp5_ASAP7_75t_L g17710 ( 
.A(n_17557),
.B(n_3711),
.Y(n_17710)
);

AOI22xp5_ASAP7_75t_L g17711 ( 
.A1(n_17445),
.A2(n_3715),
.B1(n_3713),
.B2(n_3714),
.Y(n_17711)
);

INVxp67_ASAP7_75t_SL g17712 ( 
.A(n_17584),
.Y(n_17712)
);

AOI22xp5_ASAP7_75t_L g17713 ( 
.A1(n_17526),
.A2(n_3715),
.B1(n_3713),
.B2(n_3714),
.Y(n_17713)
);

INVx1_ASAP7_75t_L g17714 ( 
.A(n_17465),
.Y(n_17714)
);

AOI22xp5_ASAP7_75t_L g17715 ( 
.A1(n_17528),
.A2(n_3718),
.B1(n_3716),
.B2(n_3717),
.Y(n_17715)
);

NOR2x1_ASAP7_75t_L g17716 ( 
.A(n_17586),
.B(n_4315),
.Y(n_17716)
);

AO22x1_ASAP7_75t_L g17717 ( 
.A1(n_17538),
.A2(n_3718),
.B1(n_3716),
.B2(n_3717),
.Y(n_17717)
);

AOI22xp5_ASAP7_75t_L g17718 ( 
.A1(n_17519),
.A2(n_17534),
.B1(n_17504),
.B2(n_17513),
.Y(n_17718)
);

INVx1_ASAP7_75t_L g17719 ( 
.A(n_17487),
.Y(n_17719)
);

AOI22xp5_ASAP7_75t_L g17720 ( 
.A1(n_17587),
.A2(n_3721),
.B1(n_3719),
.B2(n_3720),
.Y(n_17720)
);

AOI22xp5_ASAP7_75t_L g17721 ( 
.A1(n_17505),
.A2(n_3721),
.B1(n_3719),
.B2(n_3720),
.Y(n_17721)
);

INVx1_ASAP7_75t_L g17722 ( 
.A(n_17554),
.Y(n_17722)
);

AOI31xp33_ASAP7_75t_L g17723 ( 
.A1(n_17532),
.A2(n_3724),
.A3(n_3722),
.B(n_3723),
.Y(n_17723)
);

NAND2xp5_ASAP7_75t_L g17724 ( 
.A(n_17717),
.B(n_17577),
.Y(n_17724)
);

BUFx2_ASAP7_75t_L g17725 ( 
.A(n_17648),
.Y(n_17725)
);

NOR3xp33_ASAP7_75t_L g17726 ( 
.A(n_17603),
.B(n_17529),
.C(n_17530),
.Y(n_17726)
);

HB1xp67_ASAP7_75t_L g17727 ( 
.A(n_17656),
.Y(n_17727)
);

NOR2x1p5_ASAP7_75t_L g17728 ( 
.A(n_17622),
.B(n_17496),
.Y(n_17728)
);

AOI21xp5_ASAP7_75t_L g17729 ( 
.A1(n_17651),
.A2(n_17589),
.B(n_17509),
.Y(n_17729)
);

BUFx4f_ASAP7_75t_SL g17730 ( 
.A(n_17675),
.Y(n_17730)
);

NAND2xp5_ASAP7_75t_L g17731 ( 
.A(n_17650),
.B(n_17491),
.Y(n_17731)
);

NAND2xp33_ASAP7_75t_SL g17732 ( 
.A(n_17674),
.B(n_17553),
.Y(n_17732)
);

NAND2xp5_ASAP7_75t_L g17733 ( 
.A(n_17623),
.B(n_17470),
.Y(n_17733)
);

INVxp67_ASAP7_75t_L g17734 ( 
.A(n_17624),
.Y(n_17734)
);

INVx1_ASAP7_75t_SL g17735 ( 
.A(n_17635),
.Y(n_17735)
);

NAND2xp5_ASAP7_75t_L g17736 ( 
.A(n_17713),
.B(n_17523),
.Y(n_17736)
);

INVx1_ASAP7_75t_L g17737 ( 
.A(n_17642),
.Y(n_17737)
);

AND3x1_ASAP7_75t_L g17738 ( 
.A(n_17606),
.B(n_17494),
.C(n_17599),
.Y(n_17738)
);

NAND2xp5_ASAP7_75t_L g17739 ( 
.A(n_17627),
.B(n_17541),
.Y(n_17739)
);

NAND3xp33_ASAP7_75t_L g17740 ( 
.A(n_17681),
.B(n_17501),
.C(n_17483),
.Y(n_17740)
);

AND2x2_ASAP7_75t_L g17741 ( 
.A(n_17692),
.B(n_17458),
.Y(n_17741)
);

AND2x2_ASAP7_75t_L g17742 ( 
.A(n_17716),
.B(n_17527),
.Y(n_17742)
);

OR2x2_ASAP7_75t_L g17743 ( 
.A(n_17609),
.B(n_17694),
.Y(n_17743)
);

CKINVDCx20_ASAP7_75t_R g17744 ( 
.A(n_17612),
.Y(n_17744)
);

AOI311xp33_ASAP7_75t_L g17745 ( 
.A1(n_17673),
.A2(n_17507),
.A3(n_17521),
.B(n_17548),
.C(n_17542),
.Y(n_17745)
);

INVx1_ASAP7_75t_SL g17746 ( 
.A(n_17663),
.Y(n_17746)
);

NAND2xp5_ASAP7_75t_SL g17747 ( 
.A(n_17638),
.B(n_17549),
.Y(n_17747)
);

INVxp67_ASAP7_75t_L g17748 ( 
.A(n_17640),
.Y(n_17748)
);

NAND2xp5_ASAP7_75t_L g17749 ( 
.A(n_17695),
.B(n_17715),
.Y(n_17749)
);

AND2x2_ASAP7_75t_L g17750 ( 
.A(n_17662),
.B(n_17567),
.Y(n_17750)
);

NAND3xp33_ASAP7_75t_L g17751 ( 
.A(n_17711),
.B(n_17671),
.C(n_17619),
.Y(n_17751)
);

INVx1_ASAP7_75t_L g17752 ( 
.A(n_17646),
.Y(n_17752)
);

NOR2x1_ASAP7_75t_L g17753 ( 
.A(n_17653),
.B(n_17456),
.Y(n_17753)
);

AOI22xp5_ASAP7_75t_L g17754 ( 
.A1(n_17644),
.A2(n_17497),
.B1(n_3726),
.B2(n_3722),
.Y(n_17754)
);

NAND2xp5_ASAP7_75t_L g17755 ( 
.A(n_17720),
.B(n_3725),
.Y(n_17755)
);

NAND2xp5_ASAP7_75t_L g17756 ( 
.A(n_17620),
.B(n_3725),
.Y(n_17756)
);

NAND2xp5_ASAP7_75t_L g17757 ( 
.A(n_17630),
.B(n_3726),
.Y(n_17757)
);

INVx1_ASAP7_75t_L g17758 ( 
.A(n_17616),
.Y(n_17758)
);

INVx1_ASAP7_75t_L g17759 ( 
.A(n_17643),
.Y(n_17759)
);

NOR3xp33_ASAP7_75t_L g17760 ( 
.A(n_17628),
.B(n_3727),
.C(n_3728),
.Y(n_17760)
);

INVx1_ASAP7_75t_L g17761 ( 
.A(n_17669),
.Y(n_17761)
);

AND2x2_ASAP7_75t_L g17762 ( 
.A(n_17668),
.B(n_3728),
.Y(n_17762)
);

NOR3xp33_ASAP7_75t_L g17763 ( 
.A(n_17634),
.B(n_17645),
.C(n_17657),
.Y(n_17763)
);

NAND2xp5_ASAP7_75t_L g17764 ( 
.A(n_17633),
.B(n_3729),
.Y(n_17764)
);

AOI221xp5_ASAP7_75t_L g17765 ( 
.A1(n_17708),
.A2(n_3731),
.B1(n_3729),
.B2(n_3730),
.C(n_3732),
.Y(n_17765)
);

NAND2xp5_ASAP7_75t_L g17766 ( 
.A(n_17723),
.B(n_3730),
.Y(n_17766)
);

NOR2x1_ASAP7_75t_L g17767 ( 
.A(n_17659),
.B(n_3731),
.Y(n_17767)
);

OAI21xp5_ASAP7_75t_L g17768 ( 
.A1(n_17618),
.A2(n_3732),
.B(n_3734),
.Y(n_17768)
);

NAND3xp33_ASAP7_75t_L g17769 ( 
.A(n_17660),
.B(n_3742),
.C(n_3734),
.Y(n_17769)
);

AOI22xp5_ASAP7_75t_L g17770 ( 
.A1(n_17719),
.A2(n_17626),
.B1(n_17682),
.B2(n_17696),
.Y(n_17770)
);

INVx1_ASAP7_75t_L g17771 ( 
.A(n_17672),
.Y(n_17771)
);

NAND2xp5_ASAP7_75t_L g17772 ( 
.A(n_17636),
.B(n_3735),
.Y(n_17772)
);

INVx1_ASAP7_75t_L g17773 ( 
.A(n_17665),
.Y(n_17773)
);

NAND3xp33_ASAP7_75t_L g17774 ( 
.A(n_17700),
.B(n_3744),
.C(n_3735),
.Y(n_17774)
);

INVx2_ASAP7_75t_L g17775 ( 
.A(n_17691),
.Y(n_17775)
);

INVx1_ASAP7_75t_L g17776 ( 
.A(n_17697),
.Y(n_17776)
);

AND3x1_ASAP7_75t_L g17777 ( 
.A(n_17610),
.B(n_3736),
.C(n_3737),
.Y(n_17777)
);

NAND2xp5_ASAP7_75t_L g17778 ( 
.A(n_17615),
.B(n_3736),
.Y(n_17778)
);

INVx1_ASAP7_75t_L g17779 ( 
.A(n_17710),
.Y(n_17779)
);

INVx1_ASAP7_75t_L g17780 ( 
.A(n_17664),
.Y(n_17780)
);

NAND2x2_ASAP7_75t_L g17781 ( 
.A(n_17687),
.B(n_3737),
.Y(n_17781)
);

NOR2x1_ASAP7_75t_L g17782 ( 
.A(n_17670),
.B(n_3738),
.Y(n_17782)
);

INVx1_ASAP7_75t_L g17783 ( 
.A(n_17676),
.Y(n_17783)
);

NOR2xp33_ASAP7_75t_L g17784 ( 
.A(n_17655),
.B(n_3739),
.Y(n_17784)
);

NOR3x1_ASAP7_75t_L g17785 ( 
.A(n_17689),
.B(n_17712),
.C(n_17677),
.Y(n_17785)
);

INVx1_ASAP7_75t_L g17786 ( 
.A(n_17601),
.Y(n_17786)
);

NAND2xp5_ASAP7_75t_L g17787 ( 
.A(n_17702),
.B(n_3739),
.Y(n_17787)
);

NAND2xp5_ASAP7_75t_L g17788 ( 
.A(n_17641),
.B(n_3740),
.Y(n_17788)
);

NAND2xp5_ASAP7_75t_L g17789 ( 
.A(n_17632),
.B(n_3740),
.Y(n_17789)
);

AND2x2_ASAP7_75t_L g17790 ( 
.A(n_17637),
.B(n_3741),
.Y(n_17790)
);

NOR3x1_ASAP7_75t_L g17791 ( 
.A(n_17688),
.B(n_4306),
.C(n_4305),
.Y(n_17791)
);

NOR2xp33_ASAP7_75t_L g17792 ( 
.A(n_17666),
.B(n_3743),
.Y(n_17792)
);

INVx1_ASAP7_75t_SL g17793 ( 
.A(n_17658),
.Y(n_17793)
);

HB1xp67_ASAP7_75t_L g17794 ( 
.A(n_17652),
.Y(n_17794)
);

XNOR2x2_ASAP7_75t_L g17795 ( 
.A(n_17701),
.B(n_3743),
.Y(n_17795)
);

INVxp67_ASAP7_75t_L g17796 ( 
.A(n_17698),
.Y(n_17796)
);

BUFx2_ASAP7_75t_L g17797 ( 
.A(n_17706),
.Y(n_17797)
);

NOR2xp67_ASAP7_75t_SL g17798 ( 
.A(n_17661),
.B(n_17604),
.Y(n_17798)
);

NAND3xp33_ASAP7_75t_L g17799 ( 
.A(n_17714),
.B(n_3754),
.C(n_3744),
.Y(n_17799)
);

OR2x2_ASAP7_75t_L g17800 ( 
.A(n_17721),
.B(n_3746),
.Y(n_17800)
);

OR2x2_ASAP7_75t_L g17801 ( 
.A(n_17683),
.B(n_3746),
.Y(n_17801)
);

AOI21xp5_ASAP7_75t_L g17802 ( 
.A1(n_17693),
.A2(n_3747),
.B(n_3748),
.Y(n_17802)
);

INVx1_ASAP7_75t_L g17803 ( 
.A(n_17611),
.Y(n_17803)
);

OAI221xp5_ASAP7_75t_SL g17804 ( 
.A1(n_17684),
.A2(n_17718),
.B1(n_17705),
.B2(n_17703),
.C(n_17699),
.Y(n_17804)
);

OAI221xp5_ASAP7_75t_L g17805 ( 
.A1(n_17607),
.A2(n_3749),
.B1(n_3747),
.B2(n_3748),
.C(n_3750),
.Y(n_17805)
);

AOI21xp5_ASAP7_75t_L g17806 ( 
.A1(n_17679),
.A2(n_3750),
.B(n_3751),
.Y(n_17806)
);

AND2x2_ASAP7_75t_L g17807 ( 
.A(n_17704),
.B(n_3751),
.Y(n_17807)
);

NOR3xp33_ASAP7_75t_L g17808 ( 
.A(n_17614),
.B(n_3753),
.C(n_3754),
.Y(n_17808)
);

NAND2xp5_ASAP7_75t_L g17809 ( 
.A(n_17709),
.B(n_3753),
.Y(n_17809)
);

NAND3x1_ASAP7_75t_SL g17810 ( 
.A(n_17639),
.B(n_3755),
.C(n_3756),
.Y(n_17810)
);

NAND2xp5_ASAP7_75t_L g17811 ( 
.A(n_17608),
.B(n_3755),
.Y(n_17811)
);

BUFx6f_ASAP7_75t_L g17812 ( 
.A(n_17617),
.Y(n_17812)
);

INVx2_ASAP7_75t_L g17813 ( 
.A(n_17691),
.Y(n_17813)
);

NAND2x1p5_ASAP7_75t_L g17814 ( 
.A(n_17785),
.B(n_17722),
.Y(n_17814)
);

INVx2_ASAP7_75t_L g17815 ( 
.A(n_17791),
.Y(n_17815)
);

NOR2x1p5_ASAP7_75t_L g17816 ( 
.A(n_17766),
.B(n_17629),
.Y(n_17816)
);

OAI221xp5_ASAP7_75t_L g17817 ( 
.A1(n_17765),
.A2(n_17647),
.B1(n_17602),
.B2(n_17685),
.C(n_17667),
.Y(n_17817)
);

AOI22xp5_ASAP7_75t_L g17818 ( 
.A1(n_17744),
.A2(n_17686),
.B1(n_17678),
.B2(n_17690),
.Y(n_17818)
);

OA22x2_ASAP7_75t_L g17819 ( 
.A1(n_17754),
.A2(n_17605),
.B1(n_17600),
.B2(n_17649),
.Y(n_17819)
);

O2A1O1Ixp33_ASAP7_75t_L g17820 ( 
.A1(n_17727),
.A2(n_17654),
.B(n_17621),
.C(n_17680),
.Y(n_17820)
);

AND2x4_ASAP7_75t_L g17821 ( 
.A(n_17790),
.B(n_17753),
.Y(n_17821)
);

NOR2x1_ASAP7_75t_L g17822 ( 
.A(n_17767),
.B(n_17680),
.Y(n_17822)
);

NOR2xp33_ASAP7_75t_L g17823 ( 
.A(n_17756),
.B(n_17613),
.Y(n_17823)
);

AOI221x1_ASAP7_75t_L g17824 ( 
.A1(n_17763),
.A2(n_17726),
.B1(n_17732),
.B2(n_17752),
.C(n_17773),
.Y(n_17824)
);

INVx1_ASAP7_75t_L g17825 ( 
.A(n_17795),
.Y(n_17825)
);

NAND2xp5_ASAP7_75t_L g17826 ( 
.A(n_17782),
.B(n_17613),
.Y(n_17826)
);

OAI22xp5_ASAP7_75t_L g17827 ( 
.A1(n_17781),
.A2(n_17631),
.B1(n_17625),
.B2(n_17707),
.Y(n_17827)
);

AOI222xp33_ASAP7_75t_L g17828 ( 
.A1(n_17730),
.A2(n_17631),
.B1(n_17625),
.B2(n_17707),
.C1(n_3758),
.C2(n_3760),
.Y(n_17828)
);

NOR3xp33_ASAP7_75t_L g17829 ( 
.A(n_17804),
.B(n_3756),
.C(n_3757),
.Y(n_17829)
);

AO21x1_ASAP7_75t_L g17830 ( 
.A1(n_17784),
.A2(n_3760),
.B(n_3759),
.Y(n_17830)
);

INVx1_ASAP7_75t_L g17831 ( 
.A(n_17810),
.Y(n_17831)
);

NOR2xp33_ASAP7_75t_L g17832 ( 
.A(n_17762),
.B(n_3757),
.Y(n_17832)
);

INVx2_ASAP7_75t_L g17833 ( 
.A(n_17807),
.Y(n_17833)
);

NAND3xp33_ASAP7_75t_SL g17834 ( 
.A(n_17793),
.B(n_3759),
.C(n_3761),
.Y(n_17834)
);

NAND2xp5_ASAP7_75t_L g17835 ( 
.A(n_17802),
.B(n_3761),
.Y(n_17835)
);

NAND2xp5_ASAP7_75t_L g17836 ( 
.A(n_17760),
.B(n_3762),
.Y(n_17836)
);

OAI321xp33_ASAP7_75t_L g17837 ( 
.A1(n_17796),
.A2(n_3764),
.A3(n_3766),
.B1(n_3767),
.B2(n_3763),
.C(n_3765),
.Y(n_17837)
);

INVx1_ASAP7_75t_L g17838 ( 
.A(n_17777),
.Y(n_17838)
);

INVx1_ASAP7_75t_L g17839 ( 
.A(n_17811),
.Y(n_17839)
);

NOR2x1_ASAP7_75t_L g17840 ( 
.A(n_17813),
.B(n_3762),
.Y(n_17840)
);

NOR3xp33_ASAP7_75t_SL g17841 ( 
.A(n_17751),
.B(n_3771),
.C(n_3763),
.Y(n_17841)
);

OAI21xp33_ASAP7_75t_L g17842 ( 
.A1(n_17735),
.A2(n_3764),
.B(n_3765),
.Y(n_17842)
);

AOI211xp5_ASAP7_75t_L g17843 ( 
.A1(n_17805),
.A2(n_3768),
.B(n_3766),
.C(n_3767),
.Y(n_17843)
);

NAND3xp33_ASAP7_75t_SL g17844 ( 
.A(n_17725),
.B(n_17729),
.C(n_17770),
.Y(n_17844)
);

NAND3x1_ASAP7_75t_SL g17845 ( 
.A(n_17742),
.B(n_3768),
.C(n_3769),
.Y(n_17845)
);

INVxp67_ASAP7_75t_L g17846 ( 
.A(n_17792),
.Y(n_17846)
);

NOR3xp33_ASAP7_75t_L g17847 ( 
.A(n_17783),
.B(n_3769),
.C(n_3770),
.Y(n_17847)
);

INVx1_ASAP7_75t_SL g17848 ( 
.A(n_17743),
.Y(n_17848)
);

NAND2xp33_ASAP7_75t_SL g17849 ( 
.A(n_17731),
.B(n_3770),
.Y(n_17849)
);

NOR2x1_ASAP7_75t_L g17850 ( 
.A(n_17775),
.B(n_3772),
.Y(n_17850)
);

AOI22xp33_ASAP7_75t_L g17851 ( 
.A1(n_17812),
.A2(n_3774),
.B1(n_3772),
.B2(n_3773),
.Y(n_17851)
);

INVx2_ASAP7_75t_L g17852 ( 
.A(n_17800),
.Y(n_17852)
);

AOI22xp5_ASAP7_75t_L g17853 ( 
.A1(n_17758),
.A2(n_3776),
.B1(n_3777),
.B2(n_3774),
.Y(n_17853)
);

INVx1_ASAP7_75t_L g17854 ( 
.A(n_17755),
.Y(n_17854)
);

AND2x2_ASAP7_75t_L g17855 ( 
.A(n_17745),
.B(n_3773),
.Y(n_17855)
);

NOR3xp33_ASAP7_75t_L g17856 ( 
.A(n_17786),
.B(n_3776),
.C(n_3778),
.Y(n_17856)
);

OAI211xp5_ASAP7_75t_L g17857 ( 
.A1(n_17794),
.A2(n_3780),
.B(n_3778),
.C(n_3779),
.Y(n_17857)
);

NAND3x1_ASAP7_75t_SL g17858 ( 
.A(n_17750),
.B(n_3779),
.C(n_3780),
.Y(n_17858)
);

AND3x1_ASAP7_75t_L g17859 ( 
.A(n_17737),
.B(n_3781),
.C(n_3782),
.Y(n_17859)
);

OAI22xp33_ASAP7_75t_L g17860 ( 
.A1(n_17787),
.A2(n_3783),
.B1(n_3781),
.B2(n_3782),
.Y(n_17860)
);

NAND2xp5_ASAP7_75t_L g17861 ( 
.A(n_17808),
.B(n_3783),
.Y(n_17861)
);

NAND3xp33_ASAP7_75t_L g17862 ( 
.A(n_17798),
.B(n_3784),
.C(n_3785),
.Y(n_17862)
);

NAND2xp5_ASAP7_75t_L g17863 ( 
.A(n_17806),
.B(n_3785),
.Y(n_17863)
);

AO22x2_ASAP7_75t_L g17864 ( 
.A1(n_17759),
.A2(n_3788),
.B1(n_3789),
.B2(n_3787),
.Y(n_17864)
);

NOR3xp33_ASAP7_75t_L g17865 ( 
.A(n_17748),
.B(n_3786),
.C(n_3787),
.Y(n_17865)
);

AOI221xp5_ASAP7_75t_L g17866 ( 
.A1(n_17768),
.A2(n_3790),
.B1(n_3786),
.B2(n_3789),
.C(n_3791),
.Y(n_17866)
);

OAI211xp5_ASAP7_75t_L g17867 ( 
.A1(n_17724),
.A2(n_17803),
.B(n_17780),
.C(n_17761),
.Y(n_17867)
);

OR2x2_ASAP7_75t_L g17868 ( 
.A(n_17757),
.B(n_3790),
.Y(n_17868)
);

INVx2_ASAP7_75t_SL g17869 ( 
.A(n_17728),
.Y(n_17869)
);

OAI221xp5_ASAP7_75t_L g17870 ( 
.A1(n_17809),
.A2(n_3793),
.B1(n_3791),
.B2(n_3792),
.C(n_3794),
.Y(n_17870)
);

AOI222xp33_ASAP7_75t_L g17871 ( 
.A1(n_17778),
.A2(n_3795),
.B1(n_3798),
.B2(n_3792),
.C1(n_3793),
.C2(n_3796),
.Y(n_17871)
);

NAND3xp33_ASAP7_75t_L g17872 ( 
.A(n_17812),
.B(n_3795),
.C(n_3796),
.Y(n_17872)
);

NAND3x1_ASAP7_75t_L g17873 ( 
.A(n_17741),
.B(n_3798),
.C(n_3800),
.Y(n_17873)
);

INVx1_ASAP7_75t_L g17874 ( 
.A(n_17764),
.Y(n_17874)
);

HB1xp67_ASAP7_75t_L g17875 ( 
.A(n_17774),
.Y(n_17875)
);

NAND2xp5_ASAP7_75t_L g17876 ( 
.A(n_17769),
.B(n_3800),
.Y(n_17876)
);

AOI21xp5_ASAP7_75t_L g17877 ( 
.A1(n_17747),
.A2(n_17733),
.B(n_17738),
.Y(n_17877)
);

NAND3x1_ASAP7_75t_L g17878 ( 
.A(n_17771),
.B(n_3801),
.C(n_3802),
.Y(n_17878)
);

NOR2x1_ASAP7_75t_L g17879 ( 
.A(n_17799),
.B(n_3802),
.Y(n_17879)
);

NAND2x1p5_ASAP7_75t_L g17880 ( 
.A(n_17812),
.B(n_3803),
.Y(n_17880)
);

NAND2xp5_ASAP7_75t_L g17881 ( 
.A(n_17772),
.B(n_3803),
.Y(n_17881)
);

XNOR2x1_ASAP7_75t_L g17882 ( 
.A(n_17855),
.B(n_17746),
.Y(n_17882)
);

AND2x4_ASAP7_75t_L g17883 ( 
.A(n_17815),
.B(n_17824),
.Y(n_17883)
);

NOR2xp33_ASAP7_75t_SL g17884 ( 
.A(n_17848),
.B(n_17797),
.Y(n_17884)
);

HB1xp67_ASAP7_75t_L g17885 ( 
.A(n_17880),
.Y(n_17885)
);

NOR3xp33_ASAP7_75t_L g17886 ( 
.A(n_17844),
.B(n_17734),
.C(n_17776),
.Y(n_17886)
);

AOI221xp5_ASAP7_75t_L g17887 ( 
.A1(n_17849),
.A2(n_17740),
.B1(n_17788),
.B2(n_17789),
.C(n_17749),
.Y(n_17887)
);

NAND2xp5_ASAP7_75t_L g17888 ( 
.A(n_17829),
.B(n_17801),
.Y(n_17888)
);

AND2x2_ASAP7_75t_L g17889 ( 
.A(n_17841),
.B(n_17739),
.Y(n_17889)
);

NOR3x2_ASAP7_75t_L g17890 ( 
.A(n_17868),
.B(n_17822),
.C(n_17828),
.Y(n_17890)
);

CKINVDCx5p33_ASAP7_75t_R g17891 ( 
.A(n_17821),
.Y(n_17891)
);

NAND2xp33_ASAP7_75t_L g17892 ( 
.A(n_17840),
.B(n_17736),
.Y(n_17892)
);

INVx1_ASAP7_75t_L g17893 ( 
.A(n_17850),
.Y(n_17893)
);

OAI222xp33_ASAP7_75t_L g17894 ( 
.A1(n_17879),
.A2(n_17779),
.B1(n_3808),
.B2(n_3810),
.C1(n_3811),
.C2(n_3806),
.Y(n_17894)
);

NOR4xp75_ASAP7_75t_L g17895 ( 
.A(n_17817),
.B(n_3808),
.C(n_3805),
.D(n_3806),
.Y(n_17895)
);

AOI22xp33_ASAP7_75t_L g17896 ( 
.A1(n_17834),
.A2(n_3810),
.B1(n_3805),
.B2(n_3809),
.Y(n_17896)
);

INVx1_ASAP7_75t_L g17897 ( 
.A(n_17830),
.Y(n_17897)
);

NAND3xp33_ASAP7_75t_L g17898 ( 
.A(n_17877),
.B(n_17818),
.C(n_17867),
.Y(n_17898)
);

INVx2_ASAP7_75t_L g17899 ( 
.A(n_17878),
.Y(n_17899)
);

NOR2x1_ASAP7_75t_L g17900 ( 
.A(n_17825),
.B(n_3809),
.Y(n_17900)
);

OR2x2_ASAP7_75t_L g17901 ( 
.A(n_17881),
.B(n_3811),
.Y(n_17901)
);

AOI22xp5_ASAP7_75t_L g17902 ( 
.A1(n_17869),
.A2(n_3820),
.B1(n_3828),
.B2(n_3812),
.Y(n_17902)
);

AND2x4_ASAP7_75t_L g17903 ( 
.A(n_17831),
.B(n_3812),
.Y(n_17903)
);

INVx1_ASAP7_75t_L g17904 ( 
.A(n_17858),
.Y(n_17904)
);

NOR2x1_ASAP7_75t_SL g17905 ( 
.A(n_17827),
.B(n_3813),
.Y(n_17905)
);

NOR2x1_ASAP7_75t_L g17906 ( 
.A(n_17826),
.B(n_3813),
.Y(n_17906)
);

INVx1_ASAP7_75t_L g17907 ( 
.A(n_17845),
.Y(n_17907)
);

OAI221xp5_ASAP7_75t_L g17908 ( 
.A1(n_17843),
.A2(n_17836),
.B1(n_17861),
.B2(n_17866),
.C(n_17876),
.Y(n_17908)
);

NAND2x1p5_ASAP7_75t_L g17909 ( 
.A(n_17838),
.B(n_3814),
.Y(n_17909)
);

NAND3xp33_ASAP7_75t_SL g17910 ( 
.A(n_17814),
.B(n_3815),
.C(n_3816),
.Y(n_17910)
);

NAND2xp5_ASAP7_75t_L g17911 ( 
.A(n_17832),
.B(n_3816),
.Y(n_17911)
);

AOI22xp5_ASAP7_75t_L g17912 ( 
.A1(n_17859),
.A2(n_3824),
.B1(n_3833),
.B2(n_3815),
.Y(n_17912)
);

NAND2x1p5_ASAP7_75t_L g17913 ( 
.A(n_17833),
.B(n_3817),
.Y(n_17913)
);

INVx2_ASAP7_75t_L g17914 ( 
.A(n_17873),
.Y(n_17914)
);

INVx3_ASAP7_75t_L g17915 ( 
.A(n_17819),
.Y(n_17915)
);

INVx1_ASAP7_75t_L g17916 ( 
.A(n_17835),
.Y(n_17916)
);

NOR4xp25_ASAP7_75t_L g17917 ( 
.A(n_17820),
.B(n_3819),
.C(n_3817),
.D(n_3818),
.Y(n_17917)
);

NOR2x1_ASAP7_75t_L g17918 ( 
.A(n_17862),
.B(n_3818),
.Y(n_17918)
);

NAND2xp5_ASAP7_75t_L g17919 ( 
.A(n_17856),
.B(n_3821),
.Y(n_17919)
);

INVx2_ASAP7_75t_L g17920 ( 
.A(n_17864),
.Y(n_17920)
);

NOR3xp33_ASAP7_75t_L g17921 ( 
.A(n_17846),
.B(n_3820),
.C(n_3821),
.Y(n_17921)
);

INVx1_ASAP7_75t_SL g17922 ( 
.A(n_17863),
.Y(n_17922)
);

AOI221x1_ASAP7_75t_L g17923 ( 
.A1(n_17874),
.A2(n_3824),
.B1(n_3822),
.B2(n_3823),
.C(n_3825),
.Y(n_17923)
);

AND2x4_ASAP7_75t_L g17924 ( 
.A(n_17816),
.B(n_3822),
.Y(n_17924)
);

INVxp67_ASAP7_75t_L g17925 ( 
.A(n_17823),
.Y(n_17925)
);

AND2x4_ASAP7_75t_L g17926 ( 
.A(n_17852),
.B(n_3823),
.Y(n_17926)
);

BUFx4f_ASAP7_75t_SL g17927 ( 
.A(n_17839),
.Y(n_17927)
);

AND2x2_ASAP7_75t_SL g17928 ( 
.A(n_17875),
.B(n_3825),
.Y(n_17928)
);

AND2x2_ASAP7_75t_L g17929 ( 
.A(n_17854),
.B(n_3826),
.Y(n_17929)
);

INVx1_ASAP7_75t_L g17930 ( 
.A(n_17872),
.Y(n_17930)
);

NOR3xp33_ASAP7_75t_L g17931 ( 
.A(n_17870),
.B(n_17860),
.C(n_17857),
.Y(n_17931)
);

AOI21x1_ASAP7_75t_L g17932 ( 
.A1(n_17864),
.A2(n_3826),
.B(n_3827),
.Y(n_17932)
);

INVx2_ASAP7_75t_L g17933 ( 
.A(n_17853),
.Y(n_17933)
);

AND2x4_ASAP7_75t_L g17934 ( 
.A(n_17847),
.B(n_3829),
.Y(n_17934)
);

INVx4_ASAP7_75t_L g17935 ( 
.A(n_17865),
.Y(n_17935)
);

OR2x2_ASAP7_75t_L g17936 ( 
.A(n_17842),
.B(n_17851),
.Y(n_17936)
);

INVx1_ASAP7_75t_L g17937 ( 
.A(n_17871),
.Y(n_17937)
);

AND2x4_ASAP7_75t_L g17938 ( 
.A(n_17837),
.B(n_3830),
.Y(n_17938)
);

NOR3xp33_ASAP7_75t_L g17939 ( 
.A(n_17844),
.B(n_3830),
.C(n_3831),
.Y(n_17939)
);

NAND2x1p5_ASAP7_75t_L g17940 ( 
.A(n_17822),
.B(n_3831),
.Y(n_17940)
);

NOR3xp33_ASAP7_75t_L g17941 ( 
.A(n_17844),
.B(n_3832),
.C(n_3833),
.Y(n_17941)
);

AND2x4_ASAP7_75t_L g17942 ( 
.A(n_17815),
.B(n_3832),
.Y(n_17942)
);

AND4x1_ASAP7_75t_L g17943 ( 
.A(n_17824),
.B(n_3836),
.C(n_3834),
.D(n_3835),
.Y(n_17943)
);

AOI221x1_ASAP7_75t_L g17944 ( 
.A1(n_17877),
.A2(n_3836),
.B1(n_3834),
.B2(n_3835),
.C(n_3837),
.Y(n_17944)
);

NAND3x2_ASAP7_75t_L g17945 ( 
.A(n_17855),
.B(n_3837),
.C(n_3838),
.Y(n_17945)
);

AND2x4_ASAP7_75t_L g17946 ( 
.A(n_17815),
.B(n_3839),
.Y(n_17946)
);

NOR2x1_ASAP7_75t_L g17947 ( 
.A(n_17822),
.B(n_3840),
.Y(n_17947)
);

OAI21xp33_ASAP7_75t_L g17948 ( 
.A1(n_17855),
.A2(n_3840),
.B(n_3841),
.Y(n_17948)
);

HB1xp67_ASAP7_75t_L g17949 ( 
.A(n_17880),
.Y(n_17949)
);

AND2x2_ASAP7_75t_L g17950 ( 
.A(n_17855),
.B(n_3841),
.Y(n_17950)
);

NOR4xp75_ASAP7_75t_SL g17951 ( 
.A(n_17826),
.B(n_3844),
.C(n_3842),
.D(n_3843),
.Y(n_17951)
);

AOI211x1_ASAP7_75t_SL g17952 ( 
.A1(n_17844),
.A2(n_3845),
.B(n_3846),
.C(n_3844),
.Y(n_17952)
);

AND2x4_ASAP7_75t_L g17953 ( 
.A(n_17815),
.B(n_3843),
.Y(n_17953)
);

NAND2xp5_ASAP7_75t_SL g17954 ( 
.A(n_17829),
.B(n_4304),
.Y(n_17954)
);

INVx1_ASAP7_75t_L g17955 ( 
.A(n_17840),
.Y(n_17955)
);

AND2x2_ASAP7_75t_L g17956 ( 
.A(n_17855),
.B(n_3845),
.Y(n_17956)
);

AO22x2_ASAP7_75t_L g17957 ( 
.A1(n_17831),
.A2(n_3848),
.B1(n_3846),
.B2(n_3847),
.Y(n_17957)
);

AOI21xp5_ASAP7_75t_L g17958 ( 
.A1(n_17892),
.A2(n_3849),
.B(n_3850),
.Y(n_17958)
);

INVx2_ASAP7_75t_L g17959 ( 
.A(n_17909),
.Y(n_17959)
);

OAI22xp5_ASAP7_75t_SL g17960 ( 
.A1(n_17907),
.A2(n_3851),
.B1(n_3849),
.B2(n_3850),
.Y(n_17960)
);

AOI21xp5_ASAP7_75t_L g17961 ( 
.A1(n_17884),
.A2(n_17898),
.B(n_17883),
.Y(n_17961)
);

AND2x4_ASAP7_75t_L g17962 ( 
.A(n_17895),
.B(n_3852),
.Y(n_17962)
);

O2A1O1Ixp33_ASAP7_75t_L g17963 ( 
.A1(n_17925),
.A2(n_3855),
.B(n_3853),
.C(n_3854),
.Y(n_17963)
);

AND2x4_ASAP7_75t_L g17964 ( 
.A(n_17905),
.B(n_4318),
.Y(n_17964)
);

AOI22xp33_ASAP7_75t_L g17965 ( 
.A1(n_17945),
.A2(n_17948),
.B1(n_17956),
.B2(n_17950),
.Y(n_17965)
);

O2A1O1Ixp33_ASAP7_75t_L g17966 ( 
.A1(n_17915),
.A2(n_3856),
.B(n_3853),
.C(n_3854),
.Y(n_17966)
);

AOI322xp5_ASAP7_75t_L g17967 ( 
.A1(n_17954),
.A2(n_3861),
.A3(n_3860),
.B1(n_3858),
.B2(n_3856),
.C1(n_3857),
.C2(n_3859),
.Y(n_17967)
);

NOR3xp33_ASAP7_75t_L g17968 ( 
.A(n_17886),
.B(n_3859),
.C(n_3860),
.Y(n_17968)
);

NAND2xp5_ASAP7_75t_L g17969 ( 
.A(n_17939),
.B(n_3861),
.Y(n_17969)
);

OAI221xp5_ASAP7_75t_L g17970 ( 
.A1(n_17896),
.A2(n_3864),
.B1(n_3862),
.B2(n_3863),
.C(n_3865),
.Y(n_17970)
);

NAND2x1_ASAP7_75t_L g17971 ( 
.A(n_17947),
.B(n_3863),
.Y(n_17971)
);

INVx1_ASAP7_75t_L g17972 ( 
.A(n_17932),
.Y(n_17972)
);

NAND3xp33_ASAP7_75t_L g17973 ( 
.A(n_17891),
.B(n_17887),
.C(n_17941),
.Y(n_17973)
);

OAI21xp33_ASAP7_75t_SL g17974 ( 
.A1(n_17919),
.A2(n_3864),
.B(n_3865),
.Y(n_17974)
);

AOI21xp33_ASAP7_75t_SL g17975 ( 
.A1(n_17882),
.A2(n_3866),
.B(n_3867),
.Y(n_17975)
);

XNOR2xp5_ASAP7_75t_SL g17976 ( 
.A(n_17885),
.B(n_3867),
.Y(n_17976)
);

INVx5_ASAP7_75t_L g17977 ( 
.A(n_17889),
.Y(n_17977)
);

AOI21xp5_ASAP7_75t_L g17978 ( 
.A1(n_17920),
.A2(n_3866),
.B(n_3868),
.Y(n_17978)
);

INVx1_ASAP7_75t_L g17979 ( 
.A(n_17900),
.Y(n_17979)
);

AOI222xp33_ASAP7_75t_L g17980 ( 
.A1(n_17934),
.A2(n_3870),
.B1(n_3872),
.B2(n_3868),
.C1(n_3869),
.C2(n_3871),
.Y(n_17980)
);

AOI21xp5_ASAP7_75t_L g17981 ( 
.A1(n_17893),
.A2(n_3869),
.B(n_3871),
.Y(n_17981)
);

INVxp67_ASAP7_75t_L g17982 ( 
.A(n_17906),
.Y(n_17982)
);

OAI21xp5_ASAP7_75t_SL g17983 ( 
.A1(n_17952),
.A2(n_3872),
.B(n_3873),
.Y(n_17983)
);

OAI221xp5_ASAP7_75t_L g17984 ( 
.A1(n_17912),
.A2(n_3875),
.B1(n_3873),
.B2(n_3874),
.C(n_3876),
.Y(n_17984)
);

INVx1_ASAP7_75t_L g17985 ( 
.A(n_17940),
.Y(n_17985)
);

AOI221xp5_ASAP7_75t_L g17986 ( 
.A1(n_17917),
.A2(n_3876),
.B1(n_3874),
.B2(n_3875),
.C(n_3877),
.Y(n_17986)
);

OR2x2_ASAP7_75t_L g17987 ( 
.A(n_17910),
.B(n_17913),
.Y(n_17987)
);

OAI221xp5_ASAP7_75t_L g17988 ( 
.A1(n_17918),
.A2(n_3879),
.B1(n_3877),
.B2(n_3878),
.C(n_3880),
.Y(n_17988)
);

OAI21xp5_ASAP7_75t_L g17989 ( 
.A1(n_17938),
.A2(n_3878),
.B(n_3879),
.Y(n_17989)
);

NOR4xp75_ASAP7_75t_L g17990 ( 
.A(n_17888),
.B(n_3882),
.C(n_3880),
.D(n_3881),
.Y(n_17990)
);

INVx1_ASAP7_75t_L g17991 ( 
.A(n_17943),
.Y(n_17991)
);

NAND3x1_ASAP7_75t_L g17992 ( 
.A(n_17897),
.B(n_3883),
.C(n_3884),
.Y(n_17992)
);

INVx1_ASAP7_75t_L g17993 ( 
.A(n_17928),
.Y(n_17993)
);

NOR3xp33_ASAP7_75t_L g17994 ( 
.A(n_17949),
.B(n_3883),
.C(n_3884),
.Y(n_17994)
);

NOR2x1_ASAP7_75t_L g17995 ( 
.A(n_17955),
.B(n_3885),
.Y(n_17995)
);

AOI21xp5_ASAP7_75t_L g17996 ( 
.A1(n_17899),
.A2(n_3886),
.B(n_3887),
.Y(n_17996)
);

AOI22xp5_ASAP7_75t_L g17997 ( 
.A1(n_17927),
.A2(n_3888),
.B1(n_3886),
.B2(n_3887),
.Y(n_17997)
);

NAND2xp5_ASAP7_75t_L g17998 ( 
.A(n_17921),
.B(n_3889),
.Y(n_17998)
);

INVx1_ASAP7_75t_L g17999 ( 
.A(n_17901),
.Y(n_17999)
);

OAI21xp5_ASAP7_75t_L g18000 ( 
.A1(n_17904),
.A2(n_17937),
.B(n_17931),
.Y(n_18000)
);

NAND2xp5_ASAP7_75t_SL g18001 ( 
.A(n_17951),
.B(n_3889),
.Y(n_18001)
);

OAI21xp5_ASAP7_75t_SL g18002 ( 
.A1(n_17894),
.A2(n_3890),
.B(n_3891),
.Y(n_18002)
);

A2O1A1Ixp33_ASAP7_75t_L g18003 ( 
.A1(n_17914),
.A2(n_3892),
.B(n_3890),
.C(n_3891),
.Y(n_18003)
);

AOI221xp5_ASAP7_75t_L g18004 ( 
.A1(n_17908),
.A2(n_3895),
.B1(n_3893),
.B2(n_3894),
.C(n_3896),
.Y(n_18004)
);

INVx1_ASAP7_75t_L g18005 ( 
.A(n_17911),
.Y(n_18005)
);

AOI21xp5_ASAP7_75t_L g18006 ( 
.A1(n_17930),
.A2(n_17922),
.B(n_17933),
.Y(n_18006)
);

HB1xp67_ASAP7_75t_L g18007 ( 
.A(n_17924),
.Y(n_18007)
);

NAND4xp75_ASAP7_75t_L g18008 ( 
.A(n_17916),
.B(n_3895),
.C(n_3893),
.D(n_3894),
.Y(n_18008)
);

HB1xp67_ASAP7_75t_L g18009 ( 
.A(n_17944),
.Y(n_18009)
);

INVx2_ASAP7_75t_L g18010 ( 
.A(n_17926),
.Y(n_18010)
);

NAND2x1p5_ASAP7_75t_L g18011 ( 
.A(n_17935),
.B(n_3898),
.Y(n_18011)
);

AOI22xp5_ASAP7_75t_L g18012 ( 
.A1(n_17936),
.A2(n_3899),
.B1(n_3897),
.B2(n_3898),
.Y(n_18012)
);

INVx1_ASAP7_75t_L g18013 ( 
.A(n_17890),
.Y(n_18013)
);

OAI22xp5_ASAP7_75t_L g18014 ( 
.A1(n_17902),
.A2(n_3901),
.B1(n_3897),
.B2(n_3900),
.Y(n_18014)
);

A2O1A1Ixp33_ASAP7_75t_L g18015 ( 
.A1(n_17903),
.A2(n_3902),
.B(n_3900),
.C(n_3901),
.Y(n_18015)
);

XOR2x2_ASAP7_75t_L g18016 ( 
.A(n_17942),
.B(n_3902),
.Y(n_18016)
);

AND4x1_ASAP7_75t_L g18017 ( 
.A(n_17923),
.B(n_3905),
.C(n_3906),
.D(n_3904),
.Y(n_18017)
);

NOR3xp33_ASAP7_75t_SL g18018 ( 
.A(n_17957),
.B(n_3903),
.C(n_3905),
.Y(n_18018)
);

OR2x2_ASAP7_75t_L g18019 ( 
.A(n_17946),
.B(n_3903),
.Y(n_18019)
);

A2O1A1Ixp33_ASAP7_75t_SL g18020 ( 
.A1(n_17929),
.A2(n_3908),
.B(n_3906),
.C(n_3907),
.Y(n_18020)
);

OAI21xp5_ASAP7_75t_SL g18021 ( 
.A1(n_17953),
.A2(n_3907),
.B(n_3909),
.Y(n_18021)
);

OR2x2_ASAP7_75t_L g18022 ( 
.A(n_17957),
.B(n_3910),
.Y(n_18022)
);

AOI22xp33_ASAP7_75t_SL g18023 ( 
.A1(n_17884),
.A2(n_3914),
.B1(n_3912),
.B2(n_3913),
.Y(n_18023)
);

NAND4xp75_ASAP7_75t_L g18024 ( 
.A(n_17889),
.B(n_3916),
.C(n_3914),
.D(n_3915),
.Y(n_18024)
);

OAI322xp33_ASAP7_75t_L g18025 ( 
.A1(n_17884),
.A2(n_3922),
.A3(n_3921),
.B1(n_3918),
.B2(n_3915),
.C1(n_3917),
.C2(n_3919),
.Y(n_18025)
);

AND4x1_ASAP7_75t_L g18026 ( 
.A(n_17884),
.B(n_3919),
.C(n_3921),
.D(n_3918),
.Y(n_18026)
);

O2A1O1Ixp33_ASAP7_75t_L g18027 ( 
.A1(n_17892),
.A2(n_3923),
.B(n_3917),
.C(n_3922),
.Y(n_18027)
);

NOR3xp33_ASAP7_75t_L g18028 ( 
.A(n_17898),
.B(n_3923),
.C(n_3924),
.Y(n_18028)
);

NAND2x1p5_ASAP7_75t_L g18029 ( 
.A(n_17907),
.B(n_3925),
.Y(n_18029)
);

NOR2x1p5_ASAP7_75t_L g18030 ( 
.A(n_17915),
.B(n_3924),
.Y(n_18030)
);

INVx2_ASAP7_75t_L g18031 ( 
.A(n_17909),
.Y(n_18031)
);

NOR2x1_ASAP7_75t_L g18032 ( 
.A(n_17893),
.B(n_3925),
.Y(n_18032)
);

OAI221xp5_ASAP7_75t_L g18033 ( 
.A1(n_17948),
.A2(n_3928),
.B1(n_3926),
.B2(n_3927),
.C(n_3929),
.Y(n_18033)
);

NAND4xp75_ASAP7_75t_L g18034 ( 
.A(n_17889),
.B(n_3929),
.C(n_3926),
.D(n_3927),
.Y(n_18034)
);

OAI22xp33_ASAP7_75t_SL g18035 ( 
.A1(n_17884),
.A2(n_3932),
.B1(n_3930),
.B2(n_3931),
.Y(n_18035)
);

NAND3xp33_ASAP7_75t_L g18036 ( 
.A(n_17884),
.B(n_3930),
.C(n_3931),
.Y(n_18036)
);

OAI31xp33_ASAP7_75t_L g18037 ( 
.A1(n_17948),
.A2(n_3935),
.A3(n_3933),
.B(n_3934),
.Y(n_18037)
);

OR2x6_ASAP7_75t_L g18038 ( 
.A(n_17885),
.B(n_3933),
.Y(n_18038)
);

NAND3x1_ASAP7_75t_L g18039 ( 
.A(n_17947),
.B(n_3934),
.C(n_3935),
.Y(n_18039)
);

AOI221xp5_ASAP7_75t_L g18040 ( 
.A1(n_17948),
.A2(n_3938),
.B1(n_3936),
.B2(n_3937),
.C(n_3939),
.Y(n_18040)
);

NAND2xp5_ASAP7_75t_L g18041 ( 
.A(n_17939),
.B(n_3936),
.Y(n_18041)
);

AOI22xp33_ASAP7_75t_L g18042 ( 
.A1(n_17945),
.A2(n_3939),
.B1(n_3937),
.B2(n_3938),
.Y(n_18042)
);

NOR2x1_ASAP7_75t_L g18043 ( 
.A(n_17893),
.B(n_3940),
.Y(n_18043)
);

CKINVDCx16_ASAP7_75t_R g18044 ( 
.A(n_17885),
.Y(n_18044)
);

OAI21xp33_ASAP7_75t_L g18045 ( 
.A1(n_17884),
.A2(n_3940),
.B(n_3941),
.Y(n_18045)
);

AOI222xp33_ASAP7_75t_L g18046 ( 
.A1(n_17948),
.A2(n_3943),
.B1(n_3945),
.B2(n_3941),
.C1(n_3942),
.C2(n_3944),
.Y(n_18046)
);

BUFx2_ASAP7_75t_L g18047 ( 
.A(n_18039),
.Y(n_18047)
);

INVx2_ASAP7_75t_L g18048 ( 
.A(n_18029),
.Y(n_18048)
);

CKINVDCx16_ASAP7_75t_R g18049 ( 
.A(n_18044),
.Y(n_18049)
);

BUFx2_ASAP7_75t_L g18050 ( 
.A(n_17976),
.Y(n_18050)
);

INVx2_ASAP7_75t_L g18051 ( 
.A(n_18011),
.Y(n_18051)
);

HB1xp67_ASAP7_75t_L g18052 ( 
.A(n_17995),
.Y(n_18052)
);

INVx2_ASAP7_75t_SL g18053 ( 
.A(n_17964),
.Y(n_18053)
);

HB1xp67_ASAP7_75t_L g18054 ( 
.A(n_18032),
.Y(n_18054)
);

HB1xp67_ASAP7_75t_L g18055 ( 
.A(n_18043),
.Y(n_18055)
);

NAND2xp5_ASAP7_75t_L g18056 ( 
.A(n_17964),
.B(n_4306),
.Y(n_18056)
);

CKINVDCx5p33_ASAP7_75t_R g18057 ( 
.A(n_18013),
.Y(n_18057)
);

AOI221x1_ASAP7_75t_L g18058 ( 
.A1(n_17961),
.A2(n_3946),
.B1(n_3943),
.B2(n_3944),
.C(n_3947),
.Y(n_18058)
);

BUFx6f_ASAP7_75t_L g18059 ( 
.A(n_17977),
.Y(n_18059)
);

BUFx2_ASAP7_75t_L g18060 ( 
.A(n_17974),
.Y(n_18060)
);

INVx1_ASAP7_75t_L g18061 ( 
.A(n_18022),
.Y(n_18061)
);

CKINVDCx5p33_ASAP7_75t_R g18062 ( 
.A(n_18007),
.Y(n_18062)
);

INVxp67_ASAP7_75t_L g18063 ( 
.A(n_18030),
.Y(n_18063)
);

OR2x2_ASAP7_75t_L g18064 ( 
.A(n_17971),
.B(n_3946),
.Y(n_18064)
);

CKINVDCx20_ASAP7_75t_R g18065 ( 
.A(n_18000),
.Y(n_18065)
);

INVx1_ASAP7_75t_SL g18066 ( 
.A(n_18016),
.Y(n_18066)
);

INVx3_ASAP7_75t_SL g18067 ( 
.A(n_17977),
.Y(n_18067)
);

CKINVDCx6p67_ASAP7_75t_R g18068 ( 
.A(n_17977),
.Y(n_18068)
);

NAND5xp2_ASAP7_75t_L g18069 ( 
.A(n_17983),
.B(n_3949),
.C(n_3947),
.D(n_3948),
.E(n_3950),
.Y(n_18069)
);

BUFx2_ASAP7_75t_L g18070 ( 
.A(n_17989),
.Y(n_18070)
);

BUFx2_ASAP7_75t_L g18071 ( 
.A(n_18018),
.Y(n_18071)
);

CKINVDCx5p33_ASAP7_75t_R g18072 ( 
.A(n_18010),
.Y(n_18072)
);

BUFx12f_ASAP7_75t_L g18073 ( 
.A(n_17987),
.Y(n_18073)
);

CKINVDCx5p33_ASAP7_75t_R g18074 ( 
.A(n_17959),
.Y(n_18074)
);

INVx2_ASAP7_75t_L g18075 ( 
.A(n_17992),
.Y(n_18075)
);

INVx1_ASAP7_75t_SL g18076 ( 
.A(n_18019),
.Y(n_18076)
);

INVx1_ASAP7_75t_L g18077 ( 
.A(n_18001),
.Y(n_18077)
);

INVx1_ASAP7_75t_L g18078 ( 
.A(n_17969),
.Y(n_18078)
);

CKINVDCx5p33_ASAP7_75t_R g18079 ( 
.A(n_18031),
.Y(n_18079)
);

NOR2xp33_ASAP7_75t_L g18080 ( 
.A(n_17991),
.B(n_18002),
.Y(n_18080)
);

INVx1_ASAP7_75t_L g18081 ( 
.A(n_18041),
.Y(n_18081)
);

BUFx2_ASAP7_75t_L g18082 ( 
.A(n_17962),
.Y(n_18082)
);

BUFx2_ASAP7_75t_L g18083 ( 
.A(n_18009),
.Y(n_18083)
);

CKINVDCx5p33_ASAP7_75t_R g18084 ( 
.A(n_17985),
.Y(n_18084)
);

HB1xp67_ASAP7_75t_L g18085 ( 
.A(n_17990),
.Y(n_18085)
);

BUFx12f_ASAP7_75t_L g18086 ( 
.A(n_18006),
.Y(n_18086)
);

AOI22xp33_ASAP7_75t_SL g18087 ( 
.A1(n_17970),
.A2(n_3950),
.B1(n_3948),
.B2(n_3949),
.Y(n_18087)
);

INVx1_ASAP7_75t_L g18088 ( 
.A(n_17998),
.Y(n_18088)
);

INVx1_ASAP7_75t_L g18089 ( 
.A(n_18017),
.Y(n_18089)
);

CKINVDCx20_ASAP7_75t_R g18090 ( 
.A(n_17973),
.Y(n_18090)
);

HB1xp67_ASAP7_75t_L g18091 ( 
.A(n_17972),
.Y(n_18091)
);

INVx1_ASAP7_75t_L g18092 ( 
.A(n_17966),
.Y(n_18092)
);

BUFx2_ASAP7_75t_L g18093 ( 
.A(n_17982),
.Y(n_18093)
);

AOI221xp5_ASAP7_75t_SL g18094 ( 
.A1(n_17965),
.A2(n_3953),
.B1(n_3951),
.B2(n_3952),
.C(n_3954),
.Y(n_18094)
);

BUFx2_ASAP7_75t_L g18095 ( 
.A(n_17979),
.Y(n_18095)
);

INVx1_ASAP7_75t_L g18096 ( 
.A(n_18028),
.Y(n_18096)
);

NAND2x1_ASAP7_75t_SL g18097 ( 
.A(n_17993),
.B(n_3951),
.Y(n_18097)
);

INVx2_ASAP7_75t_L g18098 ( 
.A(n_18024),
.Y(n_18098)
);

XNOR2xp5_ASAP7_75t_L g18099 ( 
.A(n_18042),
.B(n_3952),
.Y(n_18099)
);

INVx1_ASAP7_75t_SL g18100 ( 
.A(n_17999),
.Y(n_18100)
);

HB1xp67_ASAP7_75t_L g18101 ( 
.A(n_18026),
.Y(n_18101)
);

INVx1_ASAP7_75t_L g18102 ( 
.A(n_17988),
.Y(n_18102)
);

HB1xp67_ASAP7_75t_L g18103 ( 
.A(n_18036),
.Y(n_18103)
);

CKINVDCx16_ASAP7_75t_R g18104 ( 
.A(n_18005),
.Y(n_18104)
);

BUFx12f_ASAP7_75t_L g18105 ( 
.A(n_18038),
.Y(n_18105)
);

INVx1_ASAP7_75t_L g18106 ( 
.A(n_18021),
.Y(n_18106)
);

OA21x2_ASAP7_75t_L g18107 ( 
.A1(n_17986),
.A2(n_3955),
.B(n_3956),
.Y(n_18107)
);

CKINVDCx20_ASAP7_75t_R g18108 ( 
.A(n_18014),
.Y(n_18108)
);

BUFx2_ASAP7_75t_L g18109 ( 
.A(n_18040),
.Y(n_18109)
);

AND2x4_ASAP7_75t_L g18110 ( 
.A(n_17968),
.B(n_3955),
.Y(n_18110)
);

CKINVDCx14_ASAP7_75t_R g18111 ( 
.A(n_18038),
.Y(n_18111)
);

CKINVDCx5p33_ASAP7_75t_R g18112 ( 
.A(n_18035),
.Y(n_18112)
);

AND2x2_ASAP7_75t_L g18113 ( 
.A(n_18037),
.B(n_3956),
.Y(n_18113)
);

A2O1A1Ixp33_ASAP7_75t_L g18114 ( 
.A1(n_18027),
.A2(n_3959),
.B(n_3957),
.C(n_3958),
.Y(n_18114)
);

INVx1_ASAP7_75t_SL g18115 ( 
.A(n_18034),
.Y(n_18115)
);

NAND2xp33_ASAP7_75t_L g18116 ( 
.A(n_17994),
.B(n_3959),
.Y(n_18116)
);

AND2x2_ASAP7_75t_L g18117 ( 
.A(n_18046),
.B(n_3960),
.Y(n_18117)
);

OR2x2_ASAP7_75t_L g18118 ( 
.A(n_17984),
.B(n_3960),
.Y(n_18118)
);

HB1xp67_ASAP7_75t_L g18119 ( 
.A(n_18033),
.Y(n_18119)
);

CKINVDCx5p33_ASAP7_75t_R g18120 ( 
.A(n_18023),
.Y(n_18120)
);

INVx1_ASAP7_75t_L g18121 ( 
.A(n_18045),
.Y(n_18121)
);

HB1xp67_ASAP7_75t_L g18122 ( 
.A(n_17978),
.Y(n_18122)
);

INVx2_ASAP7_75t_L g18123 ( 
.A(n_18008),
.Y(n_18123)
);

NOR3xp33_ASAP7_75t_L g18124 ( 
.A(n_18049),
.B(n_18020),
.C(n_17963),
.Y(n_18124)
);

HB1xp67_ASAP7_75t_L g18125 ( 
.A(n_18064),
.Y(n_18125)
);

CKINVDCx20_ASAP7_75t_R g18126 ( 
.A(n_18090),
.Y(n_18126)
);

O2A1O1Ixp5_ASAP7_75t_L g18127 ( 
.A1(n_18075),
.A2(n_17958),
.B(n_17996),
.C(n_17981),
.Y(n_18127)
);

INVx1_ASAP7_75t_L g18128 ( 
.A(n_18056),
.Y(n_18128)
);

INVx2_ASAP7_75t_L g18129 ( 
.A(n_18097),
.Y(n_18129)
);

INVx2_ASAP7_75t_L g18130 ( 
.A(n_18107),
.Y(n_18130)
);

OAI22xp5_ASAP7_75t_L g18131 ( 
.A1(n_18087),
.A2(n_17975),
.B1(n_18015),
.B2(n_18003),
.Y(n_18131)
);

NAND5xp2_ASAP7_75t_L g18132 ( 
.A(n_18080),
.B(n_17980),
.C(n_18004),
.D(n_17967),
.E(n_18012),
.Y(n_18132)
);

OAI22xp5_ASAP7_75t_SL g18133 ( 
.A1(n_18111),
.A2(n_17960),
.B1(n_17997),
.B2(n_18025),
.Y(n_18133)
);

INVx2_ASAP7_75t_L g18134 ( 
.A(n_18107),
.Y(n_18134)
);

NAND2xp5_ASAP7_75t_L g18135 ( 
.A(n_18110),
.B(n_3961),
.Y(n_18135)
);

AOI32xp33_ASAP7_75t_L g18136 ( 
.A1(n_18116),
.A2(n_3963),
.A3(n_3961),
.B1(n_3962),
.B2(n_3964),
.Y(n_18136)
);

INVxp67_ASAP7_75t_L g18137 ( 
.A(n_18083),
.Y(n_18137)
);

NOR3xp33_ASAP7_75t_L g18138 ( 
.A(n_18104),
.B(n_3962),
.C(n_3964),
.Y(n_18138)
);

INVx1_ASAP7_75t_L g18139 ( 
.A(n_18099),
.Y(n_18139)
);

NAND2xp5_ASAP7_75t_L g18140 ( 
.A(n_18110),
.B(n_3965),
.Y(n_18140)
);

INVx1_ASAP7_75t_L g18141 ( 
.A(n_18068),
.Y(n_18141)
);

BUFx2_ASAP7_75t_SL g18142 ( 
.A(n_18051),
.Y(n_18142)
);

XNOR2x1_ASAP7_75t_L g18143 ( 
.A(n_18062),
.B(n_3965),
.Y(n_18143)
);

NAND3xp33_ASAP7_75t_L g18144 ( 
.A(n_18057),
.B(n_3966),
.C(n_3967),
.Y(n_18144)
);

INVx1_ASAP7_75t_L g18145 ( 
.A(n_18113),
.Y(n_18145)
);

INVx1_ASAP7_75t_SL g18146 ( 
.A(n_18067),
.Y(n_18146)
);

OAI21xp5_ASAP7_75t_SL g18147 ( 
.A1(n_18100),
.A2(n_3966),
.B(n_3968),
.Y(n_18147)
);

OAI211xp5_ASAP7_75t_L g18148 ( 
.A1(n_18091),
.A2(n_3970),
.B(n_3968),
.C(n_3969),
.Y(n_18148)
);

INVxp67_ASAP7_75t_L g18149 ( 
.A(n_18085),
.Y(n_18149)
);

INVx2_ASAP7_75t_L g18150 ( 
.A(n_18059),
.Y(n_18150)
);

XNOR2xp5_ASAP7_75t_L g18151 ( 
.A(n_18065),
.B(n_3969),
.Y(n_18151)
);

INVx2_ASAP7_75t_L g18152 ( 
.A(n_18059),
.Y(n_18152)
);

AND2x4_ASAP7_75t_L g18153 ( 
.A(n_18089),
.B(n_3970),
.Y(n_18153)
);

NAND2xp5_ASAP7_75t_L g18154 ( 
.A(n_18114),
.B(n_3971),
.Y(n_18154)
);

INVx1_ASAP7_75t_L g18155 ( 
.A(n_18117),
.Y(n_18155)
);

OAI211xp5_ASAP7_75t_SL g18156 ( 
.A1(n_18063),
.A2(n_3974),
.B(n_3975),
.C(n_3973),
.Y(n_18156)
);

NAND4xp25_ASAP7_75t_L g18157 ( 
.A(n_18095),
.B(n_18093),
.C(n_18069),
.D(n_18082),
.Y(n_18157)
);

XNOR2xp5_ASAP7_75t_L g18158 ( 
.A(n_18074),
.B(n_3972),
.Y(n_18158)
);

OR2x2_ASAP7_75t_L g18159 ( 
.A(n_18118),
.B(n_3972),
.Y(n_18159)
);

AOI211xp5_ASAP7_75t_L g18160 ( 
.A1(n_18077),
.A2(n_3977),
.B(n_3974),
.C(n_3976),
.Y(n_18160)
);

AOI22xp33_ASAP7_75t_R g18161 ( 
.A1(n_18101),
.A2(n_3978),
.B1(n_3976),
.B2(n_3977),
.Y(n_18161)
);

INVxp67_ASAP7_75t_L g18162 ( 
.A(n_18052),
.Y(n_18162)
);

OAI211xp5_ASAP7_75t_SL g18163 ( 
.A1(n_18061),
.A2(n_3980),
.B(n_3981),
.C(n_3979),
.Y(n_18163)
);

INVx2_ASAP7_75t_L g18164 ( 
.A(n_18059),
.Y(n_18164)
);

NAND2xp5_ASAP7_75t_L g18165 ( 
.A(n_18053),
.B(n_3978),
.Y(n_18165)
);

OAI22x1_ASAP7_75t_L g18166 ( 
.A1(n_18079),
.A2(n_3982),
.B1(n_3983),
.B2(n_3981),
.Y(n_18166)
);

AOI221xp5_ASAP7_75t_L g18167 ( 
.A1(n_18115),
.A2(n_3983),
.B1(n_3980),
.B2(n_3982),
.C(n_3984),
.Y(n_18167)
);

OA21x2_ASAP7_75t_L g18168 ( 
.A1(n_18047),
.A2(n_3984),
.B(n_3985),
.Y(n_18168)
);

OAI22x1_ASAP7_75t_L g18169 ( 
.A1(n_18112),
.A2(n_18123),
.B1(n_18098),
.B2(n_18072),
.Y(n_18169)
);

XNOR2xp5_ASAP7_75t_L g18170 ( 
.A(n_18084),
.B(n_3985),
.Y(n_18170)
);

OR2x2_ASAP7_75t_L g18171 ( 
.A(n_18071),
.B(n_3986),
.Y(n_18171)
);

AOI322xp5_ASAP7_75t_L g18172 ( 
.A1(n_18066),
.A2(n_3991),
.A3(n_3990),
.B1(n_3988),
.B2(n_3986),
.C1(n_3987),
.C2(n_3989),
.Y(n_18172)
);

NOR2xp33_ASAP7_75t_L g18173 ( 
.A(n_18086),
.B(n_3987),
.Y(n_18173)
);

NAND2xp5_ASAP7_75t_L g18174 ( 
.A(n_18076),
.B(n_3989),
.Y(n_18174)
);

INVx1_ASAP7_75t_L g18175 ( 
.A(n_18159),
.Y(n_18175)
);

AND2x2_ASAP7_75t_L g18176 ( 
.A(n_18137),
.B(n_18060),
.Y(n_18176)
);

NAND4xp75_ASAP7_75t_L g18177 ( 
.A(n_18141),
.B(n_18088),
.C(n_18078),
.D(n_18081),
.Y(n_18177)
);

AOI21xp33_ASAP7_75t_SL g18178 ( 
.A1(n_18124),
.A2(n_18092),
.B(n_18106),
.Y(n_18178)
);

OAI321xp33_ASAP7_75t_L g18179 ( 
.A1(n_18157),
.A2(n_18096),
.A3(n_18121),
.B1(n_18102),
.B2(n_18050),
.C(n_18109),
.Y(n_18179)
);

AOI221x1_ASAP7_75t_L g18180 ( 
.A1(n_18169),
.A2(n_18048),
.B1(n_18073),
.B2(n_18105),
.C(n_18055),
.Y(n_18180)
);

AOI22xp33_ASAP7_75t_L g18181 ( 
.A1(n_18150),
.A2(n_18070),
.B1(n_18122),
.B2(n_18103),
.Y(n_18181)
);

OR2x2_ASAP7_75t_L g18182 ( 
.A(n_18154),
.B(n_18054),
.Y(n_18182)
);

NAND4xp75_ASAP7_75t_L g18183 ( 
.A(n_18152),
.B(n_18094),
.C(n_18058),
.D(n_18120),
.Y(n_18183)
);

NOR3xp33_ASAP7_75t_L g18184 ( 
.A(n_18162),
.B(n_18119),
.C(n_18108),
.Y(n_18184)
);

AOI222xp33_ASAP7_75t_L g18185 ( 
.A1(n_18146),
.A2(n_3992),
.B1(n_3994),
.B2(n_3990),
.C1(n_3991),
.C2(n_3993),
.Y(n_18185)
);

INVx2_ASAP7_75t_L g18186 ( 
.A(n_18143),
.Y(n_18186)
);

NAND4xp75_ASAP7_75t_L g18187 ( 
.A(n_18164),
.B(n_18155),
.C(n_18145),
.D(n_18139),
.Y(n_18187)
);

OAI221xp5_ASAP7_75t_L g18188 ( 
.A1(n_18149),
.A2(n_3994),
.B1(n_3992),
.B2(n_3993),
.C(n_3995),
.Y(n_18188)
);

INVx1_ASAP7_75t_L g18189 ( 
.A(n_18135),
.Y(n_18189)
);

OA21x2_ASAP7_75t_L g18190 ( 
.A1(n_18130),
.A2(n_18134),
.B(n_18129),
.Y(n_18190)
);

AND2x4_ASAP7_75t_L g18191 ( 
.A(n_18125),
.B(n_3995),
.Y(n_18191)
);

NAND4xp75_ASAP7_75t_L g18192 ( 
.A(n_18128),
.B(n_3998),
.C(n_3996),
.D(n_3997),
.Y(n_18192)
);

AOI211xp5_ASAP7_75t_SL g18193 ( 
.A1(n_18126),
.A2(n_3998),
.B(n_3996),
.C(n_3997),
.Y(n_18193)
);

INVx2_ASAP7_75t_L g18194 ( 
.A(n_18140),
.Y(n_18194)
);

OAI221xp5_ASAP7_75t_L g18195 ( 
.A1(n_18136),
.A2(n_4002),
.B1(n_4000),
.B2(n_4001),
.C(n_4003),
.Y(n_18195)
);

INVx1_ASAP7_75t_L g18196 ( 
.A(n_18142),
.Y(n_18196)
);

AOI221xp5_ASAP7_75t_L g18197 ( 
.A1(n_18131),
.A2(n_4002),
.B1(n_4000),
.B2(n_4001),
.C(n_4003),
.Y(n_18197)
);

OAI21xp5_ASAP7_75t_L g18198 ( 
.A1(n_18127),
.A2(n_4004),
.B(n_4005),
.Y(n_18198)
);

NOR2x1p5_ASAP7_75t_L g18199 ( 
.A(n_18133),
.B(n_4005),
.Y(n_18199)
);

OAI22xp5_ASAP7_75t_L g18200 ( 
.A1(n_18147),
.A2(n_4007),
.B1(n_4004),
.B2(n_4006),
.Y(n_18200)
);

O2A1O1Ixp33_ASAP7_75t_L g18201 ( 
.A1(n_18132),
.A2(n_4008),
.B(n_4009),
.C(n_4007),
.Y(n_18201)
);

AOI221xp5_ASAP7_75t_L g18202 ( 
.A1(n_18156),
.A2(n_18163),
.B1(n_18138),
.B2(n_18148),
.C(n_18167),
.Y(n_18202)
);

NOR2xp67_ASAP7_75t_SL g18203 ( 
.A(n_18144),
.B(n_4006),
.Y(n_18203)
);

NAND2x1p5_ASAP7_75t_L g18204 ( 
.A(n_18168),
.B(n_4008),
.Y(n_18204)
);

AOI22xp5_ASAP7_75t_L g18205 ( 
.A1(n_18173),
.A2(n_4017),
.B1(n_4027),
.B2(n_4009),
.Y(n_18205)
);

OAI21xp5_ASAP7_75t_L g18206 ( 
.A1(n_18158),
.A2(n_4010),
.B(n_4011),
.Y(n_18206)
);

NAND4xp75_ASAP7_75t_L g18207 ( 
.A(n_18168),
.B(n_4012),
.C(n_4010),
.D(n_4011),
.Y(n_18207)
);

OR2x2_ASAP7_75t_L g18208 ( 
.A(n_18174),
.B(n_4014),
.Y(n_18208)
);

OAI22xp33_ASAP7_75t_L g18209 ( 
.A1(n_18171),
.A2(n_18166),
.B1(n_18165),
.B2(n_18161),
.Y(n_18209)
);

NOR2x1p5_ASAP7_75t_L g18210 ( 
.A(n_18153),
.B(n_4014),
.Y(n_18210)
);

AOI22xp5_ASAP7_75t_L g18211 ( 
.A1(n_18151),
.A2(n_4023),
.B1(n_4032),
.B2(n_4013),
.Y(n_18211)
);

AOI221x1_ASAP7_75t_L g18212 ( 
.A1(n_18153),
.A2(n_4016),
.B1(n_4013),
.B2(n_4015),
.C(n_4017),
.Y(n_18212)
);

NAND2xp5_ASAP7_75t_L g18213 ( 
.A(n_18203),
.B(n_18160),
.Y(n_18213)
);

OAI22xp33_ASAP7_75t_L g18214 ( 
.A1(n_18195),
.A2(n_18170),
.B1(n_18172),
.B2(n_4018),
.Y(n_18214)
);

NOR3xp33_ASAP7_75t_SL g18215 ( 
.A(n_18179),
.B(n_4015),
.C(n_4016),
.Y(n_18215)
);

HB1xp67_ASAP7_75t_L g18216 ( 
.A(n_18199),
.Y(n_18216)
);

INVx1_ASAP7_75t_L g18217 ( 
.A(n_18204),
.Y(n_18217)
);

HB1xp67_ASAP7_75t_L g18218 ( 
.A(n_18190),
.Y(n_18218)
);

OA21x2_ASAP7_75t_L g18219 ( 
.A1(n_18180),
.A2(n_4018),
.B(n_4019),
.Y(n_18219)
);

AOI22xp5_ASAP7_75t_L g18220 ( 
.A1(n_18196),
.A2(n_18184),
.B1(n_18176),
.B2(n_18200),
.Y(n_18220)
);

INVx2_ASAP7_75t_L g18221 ( 
.A(n_18210),
.Y(n_18221)
);

INVx1_ASAP7_75t_L g18222 ( 
.A(n_18190),
.Y(n_18222)
);

AOI22xp5_ASAP7_75t_L g18223 ( 
.A1(n_18187),
.A2(n_4021),
.B1(n_4023),
.B2(n_4020),
.Y(n_18223)
);

NOR2x1_ASAP7_75t_L g18224 ( 
.A(n_18183),
.B(n_4019),
.Y(n_18224)
);

AO22x2_ASAP7_75t_L g18225 ( 
.A1(n_18177),
.A2(n_4025),
.B1(n_4020),
.B2(n_4024),
.Y(n_18225)
);

INVx1_ASAP7_75t_L g18226 ( 
.A(n_18175),
.Y(n_18226)
);

OAI22xp5_ASAP7_75t_L g18227 ( 
.A1(n_18181),
.A2(n_4027),
.B1(n_4024),
.B2(n_4025),
.Y(n_18227)
);

NOR3xp33_ASAP7_75t_L g18228 ( 
.A(n_18178),
.B(n_18186),
.C(n_18189),
.Y(n_18228)
);

INVx1_ASAP7_75t_L g18229 ( 
.A(n_18194),
.Y(n_18229)
);

BUFx2_ASAP7_75t_L g18230 ( 
.A(n_18206),
.Y(n_18230)
);

INVx2_ASAP7_75t_L g18231 ( 
.A(n_18208),
.Y(n_18231)
);

INVx1_ASAP7_75t_L g18232 ( 
.A(n_18209),
.Y(n_18232)
);

NOR2x1_ASAP7_75t_L g18233 ( 
.A(n_18182),
.B(n_4028),
.Y(n_18233)
);

NOR2xp67_ASAP7_75t_L g18234 ( 
.A(n_18198),
.B(n_4028),
.Y(n_18234)
);

INVx1_ASAP7_75t_L g18235 ( 
.A(n_18202),
.Y(n_18235)
);

BUFx3_ASAP7_75t_L g18236 ( 
.A(n_18211),
.Y(n_18236)
);

AOI22xp33_ASAP7_75t_L g18237 ( 
.A1(n_18185),
.A2(n_4031),
.B1(n_4029),
.B2(n_4030),
.Y(n_18237)
);

HB1xp67_ASAP7_75t_L g18238 ( 
.A(n_18207),
.Y(n_18238)
);

AO22x2_ASAP7_75t_L g18239 ( 
.A1(n_18192),
.A2(n_4032),
.B1(n_4029),
.B2(n_4031),
.Y(n_18239)
);

AND2x2_ASAP7_75t_L g18240 ( 
.A(n_18201),
.B(n_4033),
.Y(n_18240)
);

INVx1_ASAP7_75t_L g18241 ( 
.A(n_18205),
.Y(n_18241)
);

OAI22x1_ASAP7_75t_L g18242 ( 
.A1(n_18191),
.A2(n_4035),
.B1(n_4033),
.B2(n_4034),
.Y(n_18242)
);

AND2x4_ASAP7_75t_L g18243 ( 
.A(n_18212),
.B(n_4035),
.Y(n_18243)
);

INVx1_ASAP7_75t_SL g18244 ( 
.A(n_18191),
.Y(n_18244)
);

OR2x2_ASAP7_75t_L g18245 ( 
.A(n_18188),
.B(n_4320),
.Y(n_18245)
);

HB1xp67_ASAP7_75t_L g18246 ( 
.A(n_18193),
.Y(n_18246)
);

AO22x2_ASAP7_75t_L g18247 ( 
.A1(n_18244),
.A2(n_18197),
.B1(n_4323),
.B2(n_4324),
.Y(n_18247)
);

INVx2_ASAP7_75t_L g18248 ( 
.A(n_18219),
.Y(n_18248)
);

AOI21xp5_ASAP7_75t_L g18249 ( 
.A1(n_18218),
.A2(n_4034),
.B(n_4036),
.Y(n_18249)
);

INVx1_ASAP7_75t_L g18250 ( 
.A(n_18222),
.Y(n_18250)
);

AOI22xp33_ASAP7_75t_L g18251 ( 
.A1(n_18224),
.A2(n_4038),
.B1(n_4036),
.B2(n_4037),
.Y(n_18251)
);

INVx2_ASAP7_75t_L g18252 ( 
.A(n_18233),
.Y(n_18252)
);

AOI22x1_ASAP7_75t_SL g18253 ( 
.A1(n_18217),
.A2(n_4039),
.B1(n_4037),
.B2(n_4038),
.Y(n_18253)
);

OAI22xp5_ASAP7_75t_SL g18254 ( 
.A1(n_18238),
.A2(n_4041),
.B1(n_4039),
.B2(n_4040),
.Y(n_18254)
);

OAI22x1_ASAP7_75t_L g18255 ( 
.A1(n_18220),
.A2(n_4042),
.B1(n_4040),
.B2(n_4041),
.Y(n_18255)
);

INVx1_ASAP7_75t_L g18256 ( 
.A(n_18234),
.Y(n_18256)
);

INVx2_ASAP7_75t_L g18257 ( 
.A(n_18239),
.Y(n_18257)
);

NAND2xp5_ASAP7_75t_L g18258 ( 
.A(n_18240),
.B(n_4042),
.Y(n_18258)
);

HB1xp67_ASAP7_75t_L g18259 ( 
.A(n_18246),
.Y(n_18259)
);

AO22x2_ASAP7_75t_L g18260 ( 
.A1(n_18232),
.A2(n_4045),
.B1(n_4043),
.B2(n_4044),
.Y(n_18260)
);

AOI22xp5_ASAP7_75t_L g18261 ( 
.A1(n_18228),
.A2(n_4046),
.B1(n_4043),
.B2(n_4045),
.Y(n_18261)
);

INVx2_ASAP7_75t_L g18262 ( 
.A(n_18239),
.Y(n_18262)
);

OAI22xp5_ASAP7_75t_L g18263 ( 
.A1(n_18237),
.A2(n_4048),
.B1(n_4046),
.B2(n_4047),
.Y(n_18263)
);

AOI221x1_ASAP7_75t_L g18264 ( 
.A1(n_18226),
.A2(n_4051),
.B1(n_4047),
.B2(n_4050),
.C(n_4052),
.Y(n_18264)
);

INVx1_ASAP7_75t_L g18265 ( 
.A(n_18243),
.Y(n_18265)
);

INVx4_ASAP7_75t_L g18266 ( 
.A(n_18221),
.Y(n_18266)
);

AOI22x1_ASAP7_75t_L g18267 ( 
.A1(n_18216),
.A2(n_4058),
.B1(n_4067),
.B2(n_4050),
.Y(n_18267)
);

INVx2_ASAP7_75t_L g18268 ( 
.A(n_18245),
.Y(n_18268)
);

INVx1_ASAP7_75t_SL g18269 ( 
.A(n_18230),
.Y(n_18269)
);

INVx1_ASAP7_75t_L g18270 ( 
.A(n_18215),
.Y(n_18270)
);

OAI22xp5_ASAP7_75t_L g18271 ( 
.A1(n_18229),
.A2(n_4053),
.B1(n_4051),
.B2(n_4052),
.Y(n_18271)
);

A2O1A1Ixp33_ASAP7_75t_L g18272 ( 
.A1(n_18235),
.A2(n_18236),
.B(n_18231),
.C(n_18241),
.Y(n_18272)
);

OAI22xp5_ASAP7_75t_L g18273 ( 
.A1(n_18213),
.A2(n_4055),
.B1(n_4053),
.B2(n_4054),
.Y(n_18273)
);

XNOR2x1_ASAP7_75t_L g18274 ( 
.A(n_18214),
.B(n_4055),
.Y(n_18274)
);

INVx1_ASAP7_75t_L g18275 ( 
.A(n_18227),
.Y(n_18275)
);

OAI22xp5_ASAP7_75t_L g18276 ( 
.A1(n_18274),
.A2(n_18223),
.B1(n_18225),
.B2(n_18242),
.Y(n_18276)
);

XNOR2xp5_ASAP7_75t_L g18277 ( 
.A(n_18269),
.B(n_18225),
.Y(n_18277)
);

AOI221xp5_ASAP7_75t_L g18278 ( 
.A1(n_18250),
.A2(n_4058),
.B1(n_4056),
.B2(n_4057),
.C(n_4059),
.Y(n_18278)
);

OR2x2_ASAP7_75t_L g18279 ( 
.A(n_18248),
.B(n_4303),
.Y(n_18279)
);

NAND3xp33_ASAP7_75t_L g18280 ( 
.A(n_18272),
.B(n_4056),
.C(n_4057),
.Y(n_18280)
);

NOR2xp33_ASAP7_75t_L g18281 ( 
.A(n_18266),
.B(n_4059),
.Y(n_18281)
);

AOI22xp5_ASAP7_75t_L g18282 ( 
.A1(n_18259),
.A2(n_18270),
.B1(n_18265),
.B2(n_18258),
.Y(n_18282)
);

OAI22xp5_ASAP7_75t_L g18283 ( 
.A1(n_18247),
.A2(n_18275),
.B1(n_18262),
.B2(n_18257),
.Y(n_18283)
);

AOI22xp5_ASAP7_75t_L g18284 ( 
.A1(n_18263),
.A2(n_4063),
.B1(n_4060),
.B2(n_4062),
.Y(n_18284)
);

AOI22xp5_ASAP7_75t_L g18285 ( 
.A1(n_18256),
.A2(n_4063),
.B1(n_4060),
.B2(n_4062),
.Y(n_18285)
);

XOR2xp5_ASAP7_75t_L g18286 ( 
.A(n_18268),
.B(n_4064),
.Y(n_18286)
);

NAND4xp25_ASAP7_75t_L g18287 ( 
.A(n_18252),
.B(n_4067),
.C(n_4065),
.D(n_4066),
.Y(n_18287)
);

AOI22xp5_ASAP7_75t_L g18288 ( 
.A1(n_18251),
.A2(n_4069),
.B1(n_4066),
.B2(n_4068),
.Y(n_18288)
);

OAI22xp5_ASAP7_75t_L g18289 ( 
.A1(n_18249),
.A2(n_4071),
.B1(n_4069),
.B2(n_4070),
.Y(n_18289)
);

OAI211xp5_ASAP7_75t_SL g18290 ( 
.A1(n_18261),
.A2(n_4073),
.B(n_4070),
.C(n_4072),
.Y(n_18290)
);

INVx1_ASAP7_75t_L g18291 ( 
.A(n_18267),
.Y(n_18291)
);

AOI22xp5_ASAP7_75t_L g18292 ( 
.A1(n_18283),
.A2(n_18254),
.B1(n_18271),
.B2(n_18255),
.Y(n_18292)
);

OAI22xp5_ASAP7_75t_L g18293 ( 
.A1(n_18282),
.A2(n_18273),
.B1(n_18260),
.B2(n_18253),
.Y(n_18293)
);

AOI22xp5_ASAP7_75t_L g18294 ( 
.A1(n_18277),
.A2(n_18260),
.B1(n_18264),
.B2(n_4074),
.Y(n_18294)
);

INVx2_ASAP7_75t_L g18295 ( 
.A(n_18291),
.Y(n_18295)
);

AOI21xp5_ASAP7_75t_L g18296 ( 
.A1(n_18276),
.A2(n_4072),
.B(n_4073),
.Y(n_18296)
);

INVx1_ASAP7_75t_L g18297 ( 
.A(n_18290),
.Y(n_18297)
);

AOI21xp5_ASAP7_75t_L g18298 ( 
.A1(n_18289),
.A2(n_4074),
.B(n_4075),
.Y(n_18298)
);

OAI22xp5_ASAP7_75t_L g18299 ( 
.A1(n_18284),
.A2(n_4077),
.B1(n_4075),
.B2(n_4076),
.Y(n_18299)
);

NAND2xp5_ASAP7_75t_L g18300 ( 
.A(n_18288),
.B(n_18280),
.Y(n_18300)
);

INVx1_ASAP7_75t_L g18301 ( 
.A(n_18286),
.Y(n_18301)
);

AOI22xp33_ASAP7_75t_L g18302 ( 
.A1(n_18278),
.A2(n_4078),
.B1(n_4076),
.B2(n_4077),
.Y(n_18302)
);

OAI22xp5_ASAP7_75t_L g18303 ( 
.A1(n_18285),
.A2(n_4080),
.B1(n_4078),
.B2(n_4079),
.Y(n_18303)
);

INVx1_ASAP7_75t_L g18304 ( 
.A(n_18297),
.Y(n_18304)
);

AOI21xp33_ASAP7_75t_L g18305 ( 
.A1(n_18295),
.A2(n_18281),
.B(n_18279),
.Y(n_18305)
);

AOI22xp5_ASAP7_75t_L g18306 ( 
.A1(n_18301),
.A2(n_18287),
.B1(n_4081),
.B2(n_4079),
.Y(n_18306)
);

AOI221xp5_ASAP7_75t_L g18307 ( 
.A1(n_18293),
.A2(n_4083),
.B1(n_4080),
.B2(n_4082),
.C(n_4084),
.Y(n_18307)
);

INVx1_ASAP7_75t_L g18308 ( 
.A(n_18300),
.Y(n_18308)
);

NAND2xp5_ASAP7_75t_L g18309 ( 
.A(n_18292),
.B(n_4082),
.Y(n_18309)
);

OAI21xp5_ASAP7_75t_L g18310 ( 
.A1(n_18294),
.A2(n_4083),
.B(n_4084),
.Y(n_18310)
);

NAND2xp5_ASAP7_75t_L g18311 ( 
.A(n_18304),
.B(n_18298),
.Y(n_18311)
);

OAI322xp33_ASAP7_75t_L g18312 ( 
.A1(n_18308),
.A2(n_18303),
.A3(n_18299),
.B1(n_18296),
.B2(n_18302),
.C1(n_4087),
.C2(n_4090),
.Y(n_18312)
);

OAI322xp33_ASAP7_75t_L g18313 ( 
.A1(n_18306),
.A2(n_4090),
.A3(n_4089),
.B1(n_4087),
.B2(n_4085),
.C1(n_4086),
.C2(n_4088),
.Y(n_18313)
);

OAI322xp33_ASAP7_75t_L g18314 ( 
.A1(n_18305),
.A2(n_4093),
.A3(n_4092),
.B1(n_4089),
.B2(n_4085),
.C1(n_4088),
.C2(n_4091),
.Y(n_18314)
);

AOI22xp5_ASAP7_75t_L g18315 ( 
.A1(n_18311),
.A2(n_18310),
.B1(n_18307),
.B2(n_18309),
.Y(n_18315)
);

OR2x2_ASAP7_75t_L g18316 ( 
.A(n_18312),
.B(n_4092),
.Y(n_18316)
);

AOI21xp33_ASAP7_75t_L g18317 ( 
.A1(n_18313),
.A2(n_4093),
.B(n_4094),
.Y(n_18317)
);

INVxp67_ASAP7_75t_SL g18318 ( 
.A(n_18314),
.Y(n_18318)
);

AOI22xp33_ASAP7_75t_L g18319 ( 
.A1(n_18316),
.A2(n_4096),
.B1(n_4094),
.B2(n_4095),
.Y(n_18319)
);

AOI21xp5_ASAP7_75t_L g18320 ( 
.A1(n_18318),
.A2(n_4095),
.B(n_4096),
.Y(n_18320)
);

AOI222xp33_ASAP7_75t_L g18321 ( 
.A1(n_18315),
.A2(n_4099),
.B1(n_4102),
.B2(n_4097),
.C1(n_4098),
.C2(n_4101),
.Y(n_18321)
);

AOI21xp33_ASAP7_75t_L g18322 ( 
.A1(n_18319),
.A2(n_18317),
.B(n_4320),
.Y(n_18322)
);

HB1xp67_ASAP7_75t_L g18323 ( 
.A(n_18320),
.Y(n_18323)
);

HB1xp67_ASAP7_75t_L g18324 ( 
.A(n_18321),
.Y(n_18324)
);

INVx1_ASAP7_75t_L g18325 ( 
.A(n_18320),
.Y(n_18325)
);

AOI322xp5_ASAP7_75t_L g18326 ( 
.A1(n_18324),
.A2(n_4106),
.A3(n_4105),
.B1(n_4103),
.B2(n_4099),
.C1(n_4102),
.C2(n_4104),
.Y(n_18326)
);

AOI322xp5_ASAP7_75t_L g18327 ( 
.A1(n_18323),
.A2(n_4109),
.A3(n_4108),
.B1(n_4106),
.B2(n_4103),
.C1(n_4104),
.C2(n_4107),
.Y(n_18327)
);

AOI322xp5_ASAP7_75t_L g18328 ( 
.A1(n_18325),
.A2(n_4113),
.A3(n_4112),
.B1(n_4110),
.B2(n_4107),
.C1(n_4109),
.C2(n_4111),
.Y(n_18328)
);

OR2x6_ASAP7_75t_L g18329 ( 
.A(n_18326),
.B(n_18322),
.Y(n_18329)
);

AOI22xp33_ASAP7_75t_SL g18330 ( 
.A1(n_18329),
.A2(n_18327),
.B1(n_18328),
.B2(n_4114),
.Y(n_18330)
);

AOI21xp5_ASAP7_75t_L g18331 ( 
.A1(n_18330),
.A2(n_4110),
.B(n_4112),
.Y(n_18331)
);

AOI211xp5_ASAP7_75t_L g18332 ( 
.A1(n_18331),
.A2(n_4116),
.B(n_4114),
.C(n_4115),
.Y(n_18332)
);


endmodule