module real_aes_15630_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1648;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_1740;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_1699;
wire n_419;
wire n_1023;
wire n_730;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_1689;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_1102;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_1749;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1015;
wire n_1375;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1176;
wire n_640;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_0), .A2(n_61), .B1(n_587), .B2(n_588), .Y(n_586) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_0), .Y(n_618) );
INVx1_ASAP7_75t_L g795 ( .A(n_1), .Y(n_795) );
XNOR2xp5_ASAP7_75t_L g1132 ( .A(n_2), .B(n_1133), .Y(n_1132) );
OAI22xp33_ASAP7_75t_L g1394 ( .A1(n_3), .A2(n_309), .B1(n_378), .B2(n_685), .Y(n_1394) );
OAI22xp33_ASAP7_75t_SL g1404 ( .A1(n_3), .A2(n_309), .B1(n_459), .B2(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1295 ( .A(n_4), .Y(n_1295) );
INVx1_ASAP7_75t_L g358 ( .A(n_5), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_5), .B(n_368), .Y(n_480) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_5), .B(n_381), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_5), .B(n_253), .Y(n_1733) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_6), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g1668 ( .A1(n_7), .A2(n_257), .B1(n_975), .B2(n_1669), .Y(n_1668) );
AOI22xp33_ASAP7_75t_L g1686 ( .A1(n_7), .A2(n_199), .B1(n_951), .B2(n_965), .Y(n_1686) );
INVx1_ASAP7_75t_L g482 ( .A(n_8), .Y(n_482) );
INVx1_ASAP7_75t_L g1342 ( .A(n_9), .Y(n_1342) );
OAI22xp5_ASAP7_75t_SL g1357 ( .A1(n_10), .A2(n_223), .B1(n_405), .B2(n_1124), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g1360 ( .A1(n_10), .A2(n_223), .B1(n_777), .B2(n_1178), .Y(n_1360) );
OAI22xp33_ASAP7_75t_SL g684 ( .A1(n_11), .A2(n_330), .B1(n_597), .B2(n_685), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_11), .A2(n_181), .B1(n_459), .B2(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g1330 ( .A(n_12), .Y(n_1330) );
AOI22xp5_ASAP7_75t_L g1438 ( .A1(n_13), .A2(n_57), .B1(n_1421), .B2(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g1661 ( .A(n_14), .Y(n_1661) );
AOI22xp33_ASAP7_75t_L g1690 ( .A1(n_14), .A2(n_257), .B1(n_965), .B2(n_1185), .Y(n_1690) );
INVx1_ASAP7_75t_L g805 ( .A(n_15), .Y(n_805) );
INVx1_ASAP7_75t_L g558 ( .A(n_16), .Y(n_558) );
OAI22xp33_ASAP7_75t_L g1358 ( .A1(n_17), .A2(n_152), .B1(n_360), .B2(n_378), .Y(n_1358) );
OAI22xp33_ASAP7_75t_L g1366 ( .A1(n_17), .A2(n_152), .B1(n_457), .B2(n_789), .Y(n_1366) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_18), .A2(n_45), .B1(n_787), .B2(n_789), .Y(n_879) );
OAI22xp33_ASAP7_75t_L g896 ( .A1(n_18), .A2(n_45), .B1(n_360), .B2(n_378), .Y(n_896) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_19), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g1401 ( .A1(n_20), .A2(n_291), .B1(n_745), .B2(n_1402), .Y(n_1401) );
OAI22xp33_ASAP7_75t_L g1409 ( .A1(n_20), .A2(n_291), .B1(n_422), .B2(n_432), .Y(n_1409) );
INVx2_ASAP7_75t_L g425 ( .A(n_21), .Y(n_425) );
INVx1_ASAP7_75t_L g1201 ( .A(n_22), .Y(n_1201) );
INVx1_ASAP7_75t_L g1199 ( .A(n_23), .Y(n_1199) );
XNOR2xp5_ASAP7_75t_L g545 ( .A(n_24), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g1259 ( .A(n_25), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_26), .A2(n_180), .B1(n_957), .B2(n_960), .Y(n_956) );
AOI22xp33_ASAP7_75t_SL g984 ( .A1(n_26), .A2(n_137), .B1(n_985), .B2(n_986), .Y(n_984) );
AOI221xp5_ASAP7_75t_L g1187 ( .A1(n_27), .A2(n_91), .B1(n_820), .B2(n_968), .C(n_1188), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_27), .A2(n_44), .B1(n_986), .B2(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g847 ( .A(n_28), .Y(n_847) );
INVx1_ASAP7_75t_L g1090 ( .A(n_29), .Y(n_1090) );
INVx1_ASAP7_75t_L g998 ( .A(n_30), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g1448 ( .A1(n_30), .A2(n_218), .B1(n_1428), .B2(n_1431), .Y(n_1448) );
OAI221xp5_ASAP7_75t_L g1306 ( .A1(n_31), .A2(n_90), .B1(n_422), .B2(n_702), .C(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1320 ( .A(n_31), .Y(n_1320) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_32), .Y(n_353) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_32), .B(n_351), .Y(n_1422) );
AOI22xp5_ASAP7_75t_L g1437 ( .A1(n_33), .A2(n_195), .B1(n_1428), .B2(n_1431), .Y(n_1437) );
INVx1_ASAP7_75t_L g1146 ( .A(n_34), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1717 ( .A1(n_35), .A2(n_312), .B1(n_592), .B2(n_609), .Y(n_1717) );
INVxp67_ASAP7_75t_SL g1737 ( .A(n_35), .Y(n_1737) );
OAI22xp33_ASAP7_75t_SL g404 ( .A1(n_36), .A2(n_168), .B1(n_405), .B2(n_407), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_36), .A2(n_168), .B1(n_421), .B2(n_430), .Y(n_420) );
OAI222xp33_ASAP7_75t_L g941 ( .A1(n_37), .A2(n_205), .B1(n_328), .B2(n_621), .C1(n_622), .C2(n_942), .Y(n_941) );
OAI222xp33_ASAP7_75t_L g992 ( .A1(n_37), .A2(n_205), .B1(n_328), .B2(n_496), .C1(n_587), .C2(n_588), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g1473 ( .A1(n_38), .A2(n_272), .B1(n_1428), .B2(n_1431), .Y(n_1473) );
CKINVDCx5p33_ASAP7_75t_R g1050 ( .A(n_39), .Y(n_1050) );
INVx1_ASAP7_75t_L g1355 ( .A(n_40), .Y(n_1355) );
AOI22xp5_ASAP7_75t_L g1444 ( .A1(n_41), .A2(n_117), .B1(n_1428), .B2(n_1431), .Y(n_1444) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_42), .A2(n_185), .B1(n_856), .B2(n_857), .Y(n_855) );
OAI22xp33_ASAP7_75t_L g867 ( .A1(n_42), .A2(n_185), .B1(n_360), .B2(n_868), .Y(n_867) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_43), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_43), .A2(n_61), .B1(n_621), .B2(n_622), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g1189 ( .A1(n_44), .A2(n_75), .B1(n_820), .B2(n_968), .C(n_1190), .Y(n_1189) );
AOI22xp5_ASAP7_75t_L g1442 ( .A1(n_46), .A2(n_169), .B1(n_1421), .B2(n_1443), .Y(n_1442) );
INVx1_ASAP7_75t_L g1116 ( .A(n_47), .Y(n_1116) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_47), .A2(n_335), .B1(n_771), .B2(n_1124), .Y(n_1123) );
AOI22xp33_ASAP7_75t_SL g1722 ( .A1(n_48), .A2(n_263), .B1(n_592), .B2(n_986), .Y(n_1722) );
AOI22xp33_ASAP7_75t_L g1738 ( .A1(n_48), .A2(n_235), .B1(n_1739), .B2(n_1740), .Y(n_1738) );
INVx1_ASAP7_75t_L g902 ( .A(n_49), .Y(n_902) );
INVx1_ASAP7_75t_L g864 ( .A(n_50), .Y(n_864) );
OAI211xp5_ASAP7_75t_L g869 ( .A1(n_50), .A2(n_390), .B(n_762), .C(n_870), .Y(n_869) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_51), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g1659 ( .A(n_52), .Y(n_1659) );
INVx1_ASAP7_75t_L g1149 ( .A(n_53), .Y(n_1149) );
INVx1_ASAP7_75t_L g1382 ( .A(n_54), .Y(n_1382) );
OAI22xp33_ASAP7_75t_SL g1710 ( .A1(n_55), .A2(n_245), .B1(n_500), .B2(n_502), .Y(n_1710) );
INVx1_ASAP7_75t_L g1753 ( .A(n_55), .Y(n_1753) );
INVx1_ASAP7_75t_L g1193 ( .A(n_56), .Y(n_1193) );
AOI22xp33_ASAP7_75t_SL g1223 ( .A1(n_56), .A2(n_261), .B1(n_975), .B2(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1298 ( .A(n_58), .Y(n_1298) );
INVx1_ASAP7_75t_L g1083 ( .A(n_59), .Y(n_1083) );
XNOR2xp5_ASAP7_75t_L g758 ( .A(n_60), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g1266 ( .A(n_62), .Y(n_1266) );
INVx1_ASAP7_75t_L g1341 ( .A(n_63), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_64), .B(n_451), .Y(n_1309) );
INVxp67_ASAP7_75t_SL g1317 ( .A(n_64), .Y(n_1317) );
OAI211xp5_ASAP7_75t_SL g880 ( .A1(n_65), .A2(n_700), .B(n_780), .C(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g892 ( .A(n_65), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1552 ( .A1(n_66), .A2(n_233), .B1(n_1421), .B2(n_1439), .Y(n_1552) );
OAI211xp5_ASAP7_75t_L g672 ( .A1(n_67), .A2(n_673), .B(n_674), .C(n_678), .Y(n_672) );
INVx1_ASAP7_75t_L g699 ( .A(n_67), .Y(n_699) );
INVx1_ASAP7_75t_L g845 ( .A(n_68), .Y(n_845) );
OAI22xp33_ASAP7_75t_L g884 ( .A1(n_69), .A2(n_175), .B1(n_421), .B2(n_885), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_69), .A2(n_175), .B1(n_405), .B2(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g1339 ( .A(n_70), .Y(n_1339) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_71), .Y(n_641) );
INVx1_ASAP7_75t_L g590 ( .A(n_72), .Y(n_590) );
OAI222xp33_ASAP7_75t_L g1648 ( .A1(n_73), .A2(n_182), .B1(n_683), .B2(n_686), .C1(n_1649), .C2(n_1650), .Y(n_1648) );
OAI222xp33_ASAP7_75t_L g1675 ( .A1(n_73), .A2(n_182), .B1(n_224), .B2(n_1286), .C1(n_1676), .C2(n_1677), .Y(n_1675) );
OAI22xp33_ASAP7_75t_L g1312 ( .A1(n_74), .A2(n_187), .B1(n_459), .B2(n_940), .Y(n_1312) );
INVxp67_ASAP7_75t_SL g1319 ( .A(n_74), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_75), .A2(n_91), .B1(n_1226), .B2(n_1228), .Y(n_1225) );
INVx1_ASAP7_75t_L g1381 ( .A(n_76), .Y(n_1381) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_77), .Y(n_725) );
OAI22xp33_ASAP7_75t_L g865 ( .A1(n_78), .A2(n_172), .B1(n_421), .B2(n_430), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_78), .A2(n_172), .B1(n_407), .B2(n_771), .Y(n_872) );
INVx1_ASAP7_75t_L g595 ( .A(n_79), .Y(n_595) );
INVx1_ASAP7_75t_L g912 ( .A(n_80), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_81), .Y(n_1012) );
INVx1_ASAP7_75t_L g580 ( .A(n_82), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_83), .A2(n_171), .B1(n_1421), .B2(n_1428), .Y(n_1457) );
INVx1_ASAP7_75t_L g769 ( .A(n_84), .Y(n_769) );
OAI211xp5_ASAP7_75t_L g779 ( .A1(n_84), .A2(n_700), .B(n_780), .C(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g1297 ( .A(n_85), .Y(n_1297) );
INVx1_ASAP7_75t_L g515 ( .A(n_86), .Y(n_515) );
INVx1_ASAP7_75t_L g1143 ( .A(n_87), .Y(n_1143) );
XNOR2xp5_ASAP7_75t_L g1038 ( .A(n_88), .B(n_1039), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_89), .A2(n_290), .B1(n_1431), .B2(n_1439), .Y(n_1456) );
OAI22xp33_ASAP7_75t_L g1322 ( .A1(n_90), .A2(n_187), .B1(n_685), .B2(n_746), .Y(n_1322) );
OAI22xp5_ASAP7_75t_L g1196 ( .A1(n_92), .A2(n_196), .B1(n_422), .B2(n_459), .Y(n_1196) );
INVx1_ASAP7_75t_L g1207 ( .A(n_92), .Y(n_1207) );
AOI22xp5_ASAP7_75t_L g1420 ( .A1(n_93), .A2(n_158), .B1(n_1421), .B2(n_1425), .Y(n_1420) );
INVx1_ASAP7_75t_L g1029 ( .A(n_94), .Y(n_1029) );
OAI211xp5_ASAP7_75t_L g1034 ( .A1(n_94), .A2(n_444), .B(n_524), .C(n_1035), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_95), .A2(n_267), .B1(n_685), .B2(n_738), .Y(n_737) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_95), .A2(n_131), .B1(n_432), .B2(n_459), .Y(n_749) );
INVx1_ASAP7_75t_L g911 ( .A(n_96), .Y(n_911) );
INVx1_ASAP7_75t_L g1311 ( .A(n_97), .Y(n_1311) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_98), .Y(n_741) );
CKINVDCx5p33_ASAP7_75t_R g710 ( .A(n_99), .Y(n_710) );
CKINVDCx5p33_ASAP7_75t_R g639 ( .A(n_100), .Y(n_639) );
INVx1_ASAP7_75t_L g1202 ( .A(n_101), .Y(n_1202) );
XOR2xp5_ASAP7_75t_L g634 ( .A(n_102), .B(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g1553 ( .A1(n_103), .A2(n_321), .B1(n_1428), .B2(n_1431), .Y(n_1553) );
INVx1_ASAP7_75t_L g1374 ( .A(n_104), .Y(n_1374) );
INVx1_ASAP7_75t_L g1147 ( .A(n_105), .Y(n_1147) );
INVx1_ASAP7_75t_L g560 ( .A(n_106), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_106), .A2(n_283), .B1(n_608), .B2(n_615), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_107), .Y(n_1054) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_108), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g1170 ( .A1(n_109), .A2(n_142), .B1(n_378), .B2(n_685), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_109), .A2(n_129), .B1(n_421), .B2(n_459), .Y(n_1172) );
INVx1_ASAP7_75t_L g1139 ( .A(n_110), .Y(n_1139) );
INVx1_ASAP7_75t_L g1151 ( .A(n_111), .Y(n_1151) );
OAI211xp5_ASAP7_75t_L g1025 ( .A1(n_112), .A2(n_674), .B(n_927), .C(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1036 ( .A(n_112), .Y(n_1036) );
INVx1_ASAP7_75t_L g351 ( .A(n_113), .Y(n_351) );
INVx1_ASAP7_75t_L g1333 ( .A(n_114), .Y(n_1333) );
INVx1_ASAP7_75t_L g576 ( .A(n_115), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g1031 ( .A1(n_116), .A2(n_287), .B1(n_378), .B2(n_406), .Y(n_1031) );
OAI22xp33_ASAP7_75t_L g1037 ( .A1(n_116), .A2(n_160), .B1(n_422), .B2(n_432), .Y(n_1037) );
INVx1_ASAP7_75t_L g800 ( .A(n_118), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g1709 ( .A1(n_119), .A2(n_154), .B1(n_728), .B2(n_729), .Y(n_1709) );
NOR2xp33_ASAP7_75t_L g1757 ( .A(n_119), .B(n_939), .Y(n_1757) );
INVx1_ASAP7_75t_L g399 ( .A(n_120), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g1166 ( .A(n_121), .Y(n_1166) );
XOR2xp5_ASAP7_75t_L g1641 ( .A(n_122), .B(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g555 ( .A(n_123), .Y(n_555) );
INVx1_ASAP7_75t_L g489 ( .A(n_124), .Y(n_489) );
INVx1_ASAP7_75t_L g1385 ( .A(n_125), .Y(n_1385) );
AOI22xp33_ASAP7_75t_SL g1472 ( .A1(n_126), .A2(n_211), .B1(n_1421), .B2(n_1439), .Y(n_1472) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_127), .A2(n_255), .B1(n_939), .B2(n_940), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_127), .A2(n_255), .B1(n_597), .B2(n_771), .Y(n_991) );
INVx1_ASAP7_75t_L g1262 ( .A(n_128), .Y(n_1262) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_129), .A2(n_219), .B1(n_771), .B2(n_1169), .Y(n_1168) );
OAI22xp33_ASAP7_75t_SL g744 ( .A1(n_130), .A2(n_131), .B1(n_745), .B2(n_746), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_130), .A2(n_135), .B1(n_696), .B2(n_697), .Y(n_753) );
INVx1_ASAP7_75t_L g915 ( .A(n_132), .Y(n_915) );
INVx1_ASAP7_75t_L g1265 ( .A(n_133), .Y(n_1265) );
INVx1_ASAP7_75t_L g1397 ( .A(n_134), .Y(n_1397) );
INVx1_ASAP7_75t_L g742 ( .A(n_135), .Y(n_742) );
INVx1_ASAP7_75t_L g843 ( .A(n_136), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_137), .A2(n_281), .B1(n_967), .B2(n_968), .Y(n_966) );
INVx1_ASAP7_75t_L g1263 ( .A(n_138), .Y(n_1263) );
AOI31xp33_ASAP7_75t_L g1182 ( .A1(n_139), .A2(n_1183), .A3(n_1195), .B(n_1205), .Y(n_1182) );
NAND2xp33_ASAP7_75t_SL g1221 ( .A(n_139), .B(n_1222), .Y(n_1221) );
INVxp67_ASAP7_75t_SL g1234 ( .A(n_139), .Y(n_1234) );
OAI22xp33_ASAP7_75t_L g1067 ( .A1(n_140), .A2(n_188), .B1(n_378), .B2(n_745), .Y(n_1067) );
OAI22xp33_ASAP7_75t_L g1073 ( .A1(n_140), .A2(n_179), .B1(n_422), .B2(n_432), .Y(n_1073) );
CKINVDCx5p33_ASAP7_75t_R g1052 ( .A(n_141), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1177 ( .A1(n_142), .A2(n_219), .B1(n_789), .B2(n_1178), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_143), .Y(n_717) );
CKINVDCx5p33_ASAP7_75t_R g1043 ( .A(n_144), .Y(n_1043) );
OAI211xp5_ASAP7_75t_L g384 ( .A1(n_145), .A2(n_385), .B(n_390), .C(n_395), .Y(n_384) );
INVx1_ASAP7_75t_L g453 ( .A(n_145), .Y(n_453) );
OAI221xp5_ASAP7_75t_L g1725 ( .A1(n_146), .A2(n_316), .B1(n_1051), .B2(n_1726), .C(n_1729), .Y(n_1725) );
INVx1_ASAP7_75t_L g1749 ( .A(n_146), .Y(n_1749) );
INVx1_ASAP7_75t_L g403 ( .A(n_147), .Y(n_403) );
OAI211xp5_ASAP7_75t_L g436 ( .A1(n_147), .A2(n_437), .B(n_444), .C(n_448), .Y(n_436) );
INVx1_ASAP7_75t_L g906 ( .A(n_148), .Y(n_906) );
INVx1_ASAP7_75t_L g1714 ( .A(n_149), .Y(n_1714) );
AOI22xp33_ASAP7_75t_L g1743 ( .A1(n_149), .A2(n_263), .B1(n_1308), .B2(n_1739), .Y(n_1743) );
INVx1_ASAP7_75t_L g1376 ( .A(n_150), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g1719 ( .A(n_151), .Y(n_1719) );
INVx1_ASAP7_75t_L g882 ( .A(n_153), .Y(n_882) );
INVx1_ASAP7_75t_L g1751 ( .A(n_154), .Y(n_1751) );
INVx1_ASAP7_75t_L g484 ( .A(n_155), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_156), .Y(n_643) );
INVx1_ASAP7_75t_L g1141 ( .A(n_157), .Y(n_1141) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_159), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_160), .A2(n_269), .B1(n_685), .B2(n_773), .Y(n_1030) );
INVx1_ASAP7_75t_L g1065 ( .A(n_161), .Y(n_1065) );
OAI211xp5_ASAP7_75t_L g1070 ( .A1(n_161), .A2(n_444), .B(n_524), .C(n_1071), .Y(n_1070) );
CKINVDCx5p33_ASAP7_75t_R g1003 ( .A(n_162), .Y(n_1003) );
INVx1_ASAP7_75t_L g1294 ( .A(n_163), .Y(n_1294) );
OAI211xp5_ASAP7_75t_SL g1353 ( .A1(n_164), .A2(n_390), .B(n_762), .C(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g1365 ( .A(n_164), .Y(n_1365) );
INVx1_ASAP7_75t_L g1260 ( .A(n_165), .Y(n_1260) );
INVx1_ASAP7_75t_L g768 ( .A(n_166), .Y(n_768) );
OAI211xp5_ASAP7_75t_L g1062 ( .A1(n_167), .A2(n_674), .B(n_927), .C(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1072 ( .A(n_167), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1695 ( .A1(n_169), .A2(n_1696), .B1(n_1699), .B2(n_1758), .Y(n_1695) );
INVx1_ASAP7_75t_L g1702 ( .A(n_169), .Y(n_1702) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_170), .Y(n_649) );
INVx1_ASAP7_75t_L g514 ( .A(n_173), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_174), .A2(n_254), .B1(n_771), .B2(n_772), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_174), .A2(n_254), .B1(n_777), .B2(n_778), .Y(n_776) );
OAI22xp33_ASAP7_75t_L g1066 ( .A1(n_176), .A2(n_179), .B1(n_685), .B2(n_773), .Y(n_1066) );
OAI22xp33_ASAP7_75t_L g1069 ( .A1(n_176), .A2(n_188), .B1(n_459), .B2(n_702), .Y(n_1069) );
INVx1_ASAP7_75t_L g883 ( .A(n_177), .Y(n_883) );
OAI211xp5_ASAP7_75t_L g889 ( .A1(n_177), .A2(n_385), .B(n_390), .C(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g809 ( .A(n_178), .Y(n_809) );
AOI22xp33_ASAP7_75t_SL g976 ( .A1(n_180), .A2(n_281), .B1(n_977), .B2(n_981), .Y(n_976) );
OAI22xp33_ASAP7_75t_SL g687 ( .A1(n_181), .A2(n_294), .B1(n_378), .B2(n_406), .Y(n_687) );
INVx1_ASAP7_75t_L g1256 ( .A(n_183), .Y(n_1256) );
INVx2_ASAP7_75t_L g1424 ( .A(n_184), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_184), .B(n_289), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_184), .B(n_1430), .Y(n_1432) );
AO22x2_ASAP7_75t_L g1368 ( .A1(n_186), .A2(n_1369), .B1(n_1410), .B2(n_1411), .Y(n_1368) );
INVx1_ASAP7_75t_L g1410 ( .A(n_186), .Y(n_1410) );
CKINVDCx5p33_ASAP7_75t_R g1048 ( .A(n_189), .Y(n_1048) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_190), .Y(n_720) );
INVx1_ASAP7_75t_L g804 ( .A(n_191), .Y(n_804) );
INVx1_ASAP7_75t_L g903 ( .A(n_192), .Y(n_903) );
INVx1_ASAP7_75t_L g837 ( .A(n_193), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g1450 ( .A1(n_194), .A2(n_247), .B1(n_1421), .B2(n_1431), .Y(n_1450) );
XNOR2xp5_ASAP7_75t_L g1324 ( .A(n_195), .B(n_1325), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_196), .A2(n_275), .B1(n_738), .B2(n_745), .Y(n_1211) );
INVx1_ASAP7_75t_L g1167 ( .A(n_197), .Y(n_1167) );
OAI211xp5_ASAP7_75t_L g1173 ( .A1(n_197), .A2(n_444), .B(n_1174), .C(n_1175), .Y(n_1173) );
XOR2xp5_ASAP7_75t_L g1280 ( .A(n_198), .B(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1662 ( .A(n_199), .Y(n_1662) );
INVx1_ASAP7_75t_L g1118 ( .A(n_200), .Y(n_1118) );
OAI22xp33_ASAP7_75t_L g1128 ( .A1(n_200), .A2(n_230), .B1(n_378), .B2(n_685), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_201), .A2(n_319), .B1(n_948), .B2(n_964), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_201), .A2(n_246), .B1(n_977), .B2(n_981), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1451 ( .A1(n_202), .A2(n_207), .B1(n_1425), .B2(n_1428), .Y(n_1451) );
INVx1_ASAP7_75t_L g1287 ( .A(n_203), .Y(n_1287) );
INVx1_ASAP7_75t_L g1243 ( .A(n_204), .Y(n_1243) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_206), .Y(n_1009) );
INVx1_ASAP7_75t_L g1337 ( .A(n_208), .Y(n_1337) );
INVx1_ASAP7_75t_L g834 ( .A(n_209), .Y(n_834) );
OAI211xp5_ASAP7_75t_L g1645 ( .A1(n_210), .A2(n_868), .B(n_1646), .C(n_1654), .Y(n_1645) );
INVx1_ASAP7_75t_L g1680 ( .A(n_210), .Y(n_1680) );
INVx1_ASAP7_75t_L g1291 ( .A(n_212), .Y(n_1291) );
OAI22xp33_ASAP7_75t_L g377 ( .A1(n_213), .A2(n_282), .B1(n_360), .B2(n_378), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g456 ( .A1(n_213), .A2(n_282), .B1(n_457), .B2(n_460), .Y(n_456) );
INVx2_ASAP7_75t_L g469 ( .A(n_214), .Y(n_469) );
INVx1_ASAP7_75t_L g543 ( .A(n_214), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g1004 ( .A(n_215), .Y(n_1004) );
XOR2xp5_ASAP7_75t_L g828 ( .A(n_216), .B(n_829), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g1427 ( .A1(n_216), .A2(n_327), .B1(n_1428), .B2(n_1431), .Y(n_1427) );
OAI22xp33_ASAP7_75t_L g1239 ( .A1(n_217), .A2(n_274), .B1(n_738), .B2(n_745), .Y(n_1239) );
OAI22xp5_ASAP7_75t_SL g1246 ( .A1(n_217), .A2(n_244), .B1(n_422), .B2(n_459), .Y(n_1246) );
INVx1_ASAP7_75t_L g1093 ( .A(n_220), .Y(n_1093) );
XOR2xp5_ASAP7_75t_L g931 ( .A(n_221), .B(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g1653 ( .A(n_222), .Y(n_1653) );
OAI22xp5_ASAP7_75t_L g1678 ( .A1(n_222), .A2(n_252), .B1(n_422), .B2(n_432), .Y(n_1678) );
INVx1_ASAP7_75t_L g1647 ( .A(n_224), .Y(n_1647) );
INVx1_ASAP7_75t_L g1111 ( .A(n_225), .Y(n_1111) );
OA211x2_ASAP7_75t_L g1125 ( .A1(n_225), .A2(n_496), .B(n_765), .C(n_1126), .Y(n_1125) );
BUFx3_ASAP7_75t_L g427 ( .A(n_226), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g1014 ( .A(n_227), .Y(n_1014) );
CKINVDCx5p33_ASAP7_75t_R g1055 ( .A(n_228), .Y(n_1055) );
OAI22xp5_ASAP7_75t_SL g1077 ( .A1(n_229), .A2(n_1078), .B1(n_1121), .B2(n_1130), .Y(n_1077) );
NAND4xp25_ASAP7_75t_L g1078 ( .A(n_229), .B(n_1079), .C(n_1095), .D(n_1105), .Y(n_1078) );
INVx1_ASAP7_75t_L g1115 ( .A(n_230), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_231), .A2(n_246), .B1(n_948), .B2(n_954), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_231), .A2(n_319), .B1(n_973), .B2(n_974), .Y(n_972) );
INVx1_ASAP7_75t_L g565 ( .A(n_232), .Y(n_565) );
INVx1_ASAP7_75t_L g1658 ( .A(n_234), .Y(n_1658) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_234), .B(n_1688), .Y(n_1687) );
AOI21xp33_ASAP7_75t_L g1715 ( .A1(n_235), .A2(n_1226), .B(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1398 ( .A(n_236), .Y(n_1398) );
CKINVDCx5p33_ASAP7_75t_R g1047 ( .A(n_237), .Y(n_1047) );
INVx1_ASAP7_75t_L g1085 ( .A(n_238), .Y(n_1085) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_239), .Y(n_1006) );
INVx1_ASAP7_75t_L g841 ( .A(n_240), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g774 ( .A1(n_241), .A2(n_307), .B1(n_360), .B2(n_378), .Y(n_774) );
OAI22xp33_ASAP7_75t_L g786 ( .A1(n_241), .A2(n_307), .B1(n_787), .B2(n_789), .Y(n_786) );
INVx1_ASAP7_75t_L g495 ( .A(n_242), .Y(n_495) );
INVx1_ASAP7_75t_L g1242 ( .A(n_243), .Y(n_1242) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_244), .A2(n_277), .B1(n_685), .B2(n_746), .Y(n_1244) );
INVx1_ASAP7_75t_L g1756 ( .A(n_245), .Y(n_1756) );
INVx1_ASAP7_75t_L g573 ( .A(n_248), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_248), .A2(n_292), .B1(n_606), .B2(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g1373 ( .A(n_249), .Y(n_1373) );
XOR2xp5_ASAP7_75t_L g705 ( .A(n_250), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g801 ( .A(n_251), .Y(n_801) );
INVx1_ASAP7_75t_L g1655 ( .A(n_252), .Y(n_1655) );
BUFx3_ASAP7_75t_L g368 ( .A(n_253), .Y(n_368) );
INVx1_ASAP7_75t_L g381 ( .A(n_253), .Y(n_381) );
XOR2x2_ASAP7_75t_L g876 ( .A(n_256), .B(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g1110 ( .A(n_258), .Y(n_1110) );
INVx1_ASAP7_75t_L g1285 ( .A(n_259), .Y(n_1285) );
INVx1_ASAP7_75t_L g1094 ( .A(n_260), .Y(n_1094) );
AOI22xp5_ASAP7_75t_L g1184 ( .A1(n_261), .A2(n_278), .B1(n_1113), .B2(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g936 ( .A(n_262), .Y(n_936) );
INVx1_ASAP7_75t_L g833 ( .A(n_264), .Y(n_833) );
OAI211xp5_ASAP7_75t_L g1240 ( .A1(n_265), .A2(n_496), .B(n_674), .C(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1251 ( .A(n_265), .Y(n_1251) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_266), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_267), .B(n_422), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g724 ( .A(n_268), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g1033 ( .A1(n_269), .A2(n_287), .B1(n_459), .B2(n_702), .Y(n_1033) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_270), .Y(n_650) );
INVx1_ASAP7_75t_L g1089 ( .A(n_271), .Y(n_1089) );
XOR2x2_ASAP7_75t_L g374 ( .A(n_272), .B(n_375), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g1045 ( .A(n_273), .Y(n_1045) );
OAI22xp33_ASAP7_75t_L g1252 ( .A1(n_274), .A2(n_277), .B1(n_432), .B2(n_702), .Y(n_1252) );
OAI22xp5_ASAP7_75t_L g1203 ( .A1(n_275), .A2(n_310), .B1(n_432), .B2(n_702), .Y(n_1203) );
INVx1_ASAP7_75t_L g429 ( .A(n_276), .Y(n_429) );
INVx1_ASAP7_75t_L g435 ( .A(n_276), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_278), .A2(n_311), .B1(n_1226), .B2(n_1228), .Y(n_1229) );
INVx1_ASAP7_75t_L g1086 ( .A(n_279), .Y(n_1086) );
OAI211xp5_ASAP7_75t_L g858 ( .A1(n_280), .A2(n_700), .B(n_859), .C(n_861), .Y(n_858) );
INVx1_ASAP7_75t_L g871 ( .A(n_280), .Y(n_871) );
INVx1_ASAP7_75t_L g568 ( .A(n_283), .Y(n_568) );
INVx1_ASAP7_75t_L g679 ( .A(n_284), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g691 ( .A1(n_284), .A2(n_621), .B(n_692), .C(n_700), .Y(n_691) );
INVx1_ASAP7_75t_L g907 ( .A(n_285), .Y(n_907) );
AOI22xp5_ASAP7_75t_SL g1447 ( .A1(n_286), .A2(n_336), .B1(n_1421), .B2(n_1425), .Y(n_1447) );
INVx1_ASAP7_75t_L g1289 ( .A(n_288), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_289), .B(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1430 ( .A(n_289), .Y(n_1430) );
INVx1_ASAP7_75t_L g551 ( .A(n_292), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g1007 ( .A(n_293), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_294), .A2(n_330), .B1(n_422), .B2(n_432), .Y(n_690) );
INVx1_ASAP7_75t_L g935 ( .A(n_295), .Y(n_935) );
INVx1_ASAP7_75t_L g1724 ( .A(n_296), .Y(n_1724) );
INVx1_ASAP7_75t_L g579 ( .A(n_297), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g1064 ( .A(n_298), .Y(n_1064) );
INVx1_ASAP7_75t_L g1384 ( .A(n_299), .Y(n_1384) );
CKINVDCx5p33_ASAP7_75t_R g1664 ( .A(n_300), .Y(n_1664) );
OAI211xp5_ASAP7_75t_SL g739 ( .A1(n_301), .A2(n_673), .B(n_674), .C(n_740), .Y(n_739) );
OAI211xp5_ASAP7_75t_SL g750 ( .A1(n_301), .A2(n_700), .B(n_751), .C(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g1257 ( .A(n_302), .Y(n_1257) );
INVx1_ASAP7_75t_L g1356 ( .A(n_303), .Y(n_1356) );
OAI211xp5_ASAP7_75t_SL g1361 ( .A1(n_303), .A2(n_700), .B(n_1362), .C(n_1364), .Y(n_1361) );
INVx1_ASAP7_75t_L g1310 ( .A(n_304), .Y(n_1310) );
XOR2x2_ASAP7_75t_L g1236 ( .A(n_305), .B(n_1237), .Y(n_1236) );
AOI21xp5_ASAP7_75t_SL g1720 ( .A1(n_306), .A2(n_1226), .B(n_1721), .Y(n_1720) );
INVx1_ASAP7_75t_L g1736 ( .A(n_306), .Y(n_1736) );
OAI211xp5_ASAP7_75t_L g1164 ( .A1(n_308), .A2(n_734), .B(n_765), .C(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1176 ( .A(n_308), .Y(n_1176) );
INVxp67_ASAP7_75t_SL g1209 ( .A(n_310), .Y(n_1209) );
INVx1_ASAP7_75t_L g1192 ( .A(n_311), .Y(n_1192) );
INVxp67_ASAP7_75t_L g1742 ( .A(n_312), .Y(n_1742) );
OAI211xp5_ASAP7_75t_SL g761 ( .A1(n_313), .A2(n_762), .B(n_765), .C(n_766), .Y(n_761) );
INVx1_ASAP7_75t_L g784 ( .A(n_313), .Y(n_784) );
INVx1_ASAP7_75t_L g797 ( .A(n_314), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_315), .Y(n_653) );
INVxp67_ASAP7_75t_SL g1755 ( .A(n_316), .Y(n_1755) );
INVx1_ASAP7_75t_L g1082 ( .A(n_317), .Y(n_1082) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_318), .Y(n_364) );
INVx1_ASAP7_75t_L g501 ( .A(n_320), .Y(n_501) );
INVx1_ASAP7_75t_L g1377 ( .A(n_322), .Y(n_1377) );
INVx1_ASAP7_75t_L g839 ( .A(n_323), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_324), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_325), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_326), .Y(n_715) );
INVx1_ASAP7_75t_L g1400 ( .A(n_329), .Y(n_1400) );
INVx1_ASAP7_75t_L g418 ( .A(n_331), .Y(n_418) );
INVx2_ASAP7_75t_L g479 ( .A(n_331), .Y(n_479) );
INVx1_ASAP7_75t_L g542 ( .A(n_331), .Y(n_542) );
INVx1_ASAP7_75t_L g863 ( .A(n_332), .Y(n_863) );
INVx1_ASAP7_75t_L g1137 ( .A(n_333), .Y(n_1137) );
INVx1_ASAP7_75t_L g1329 ( .A(n_334), .Y(n_1329) );
INVx1_ASAP7_75t_L g1120 ( .A(n_335), .Y(n_1120) );
INVx1_ASAP7_75t_L g1332 ( .A(n_337), .Y(n_1332) );
INVx1_ASAP7_75t_L g504 ( .A(n_338), .Y(n_504) );
AOI21xp33_ASAP7_75t_L g1665 ( .A1(n_339), .A2(n_1226), .B(n_1666), .Y(n_1665) );
INVx1_ASAP7_75t_L g1683 ( .A(n_339), .Y(n_1683) );
INVx1_ASAP7_75t_L g914 ( .A(n_340), .Y(n_914) );
INVx1_ASAP7_75t_L g1112 ( .A(n_341), .Y(n_1112) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_342), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1651 ( .A(n_343), .Y(n_1651) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_369), .B(n_1413), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_354), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g1698 ( .A(n_348), .B(n_357), .Y(n_1698) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g1694 ( .A(n_350), .B(n_353), .Y(n_1694) );
INVx1_ASAP7_75t_L g1761 ( .A(n_350), .Y(n_1761) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g1763 ( .A(n_353), .B(n_1761), .Y(n_1763) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_359), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g414 ( .A(n_357), .B(n_415), .Y(n_414) );
AOI21xp5_ASAP7_75t_SL g1644 ( .A1(n_357), .A2(n_1645), .B(n_1656), .Y(n_1644) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g507 ( .A(n_358), .B(n_368), .Y(n_507) );
AND2x4_ASAP7_75t_L g1667 ( .A(n_358), .B(n_367), .Y(n_1667) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_359), .A2(n_379), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_359), .A2(n_379), .B1(n_935), .B2(n_936), .Y(n_989) );
AND2x4_ASAP7_75t_SL g1697 ( .A(n_359), .B(n_1698), .Y(n_1697) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_361), .B(n_366), .Y(n_360) );
OR2x6_ASAP7_75t_L g406 ( .A(n_361), .B(n_380), .Y(n_406) );
BUFx4f_ASAP7_75t_L g483 ( .A(n_361), .Y(n_483) );
INVx1_ASAP7_75t_L g668 ( .A(n_361), .Y(n_668) );
OR2x2_ASAP7_75t_L g745 ( .A(n_361), .B(n_380), .Y(n_745) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx4f_ASAP7_75t_L g513 ( .A(n_362), .Y(n_513) );
INVx3_ASAP7_75t_L g686 ( .A(n_362), .Y(n_686) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AND2x2_ASAP7_75t_L g382 ( .A(n_364), .B(n_383), .Y(n_382) );
NAND2x1_ASAP7_75t_L g389 ( .A(n_364), .B(n_365), .Y(n_389) );
AND2x2_ASAP7_75t_L g394 ( .A(n_364), .B(n_365), .Y(n_394) );
INVx1_ASAP7_75t_L g402 ( .A(n_364), .Y(n_402) );
INVx2_ASAP7_75t_L g412 ( .A(n_364), .Y(n_412) );
INVx2_ASAP7_75t_L g494 ( .A(n_364), .Y(n_494) );
INVx2_ASAP7_75t_L g383 ( .A(n_365), .Y(n_383) );
BUFx2_ASAP7_75t_L g398 ( .A(n_365), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_365), .B(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g493 ( .A(n_365), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g594 ( .A(n_365), .Y(n_594) );
AND2x2_ASAP7_75t_L g610 ( .A(n_365), .B(n_412), .Y(n_610) );
OR2x6_ASAP7_75t_L g685 ( .A(n_366), .B(n_686), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g1650 ( .A1(n_366), .A2(n_1651), .B1(n_1652), .B2(n_1653), .Y(n_1650) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g392 ( .A(n_367), .Y(n_392) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
AND2x4_ASAP7_75t_L g400 ( .A(n_368), .B(n_401), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_1275), .B1(n_1276), .B2(n_1412), .Y(n_369) );
INVx1_ASAP7_75t_L g1412 ( .A(n_370), .Y(n_1412) );
AO22x1_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_873), .B1(n_1273), .B2(n_1274), .Y(n_370) );
INVx1_ASAP7_75t_L g1274 ( .A(n_371), .Y(n_1274) );
XNOR2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_755), .Y(n_371) );
XOR2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_632), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_545), .B1(n_630), .B2(n_631), .Y(n_373) );
INVx2_ASAP7_75t_L g630 ( .A(n_374), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_419), .C(n_473), .Y(n_375) );
OAI31xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_384), .A3(n_404), .B(n_413), .Y(n_376) );
CKINVDCx16_ASAP7_75t_R g378 ( .A(n_379), .Y(n_378) );
INVx4_ASAP7_75t_L g746 ( .A(n_379), .Y(n_746) );
INVx3_ASAP7_75t_SL g868 ( .A(n_379), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g1206 ( .A1(n_379), .A2(n_1207), .B1(n_1208), .B2(n_1209), .Y(n_1206) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g980 ( .A(n_382), .Y(n_980) );
BUFx6f_ASAP7_75t_L g1227 ( .A(n_382), .Y(n_1227) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI221xp5_ASAP7_75t_L g602 ( .A1(n_387), .A2(n_558), .B1(n_565), .B2(n_603), .C(n_605), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_387), .A2(n_555), .B1(n_576), .B2(n_612), .C(n_614), .Y(n_611) );
BUFx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_SL g497 ( .A(n_388), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_388), .A2(n_803), .B1(n_804), .B2(n_805), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_388), .A2(n_803), .B1(n_834), .B2(n_847), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_388), .A2(n_1004), .B1(n_1015), .B2(n_1021), .Y(n_1020) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_388), .A2(n_1019), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
BUFx2_ASAP7_75t_SL g1338 ( .A(n_388), .Y(n_1338) );
BUFx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_389), .Y(n_503) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI211xp5_ASAP7_75t_L g581 ( .A1(n_391), .A2(n_582), .B(n_585), .C(n_586), .Y(n_581) );
INVx3_ASAP7_75t_L g765 ( .A(n_391), .Y(n_765) );
NOR3xp33_ASAP7_75t_L g990 ( .A(n_391), .B(n_991), .C(n_992), .Y(n_990) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
AND2x2_ASAP7_75t_L g675 ( .A(n_392), .B(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g738 ( .A(n_392), .B(n_410), .Y(n_738) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_392), .B(n_398), .Y(n_1027) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_393), .Y(n_584) );
BUFx3_ASAP7_75t_L g1228 ( .A(n_393), .Y(n_1228) );
BUFx3_ASAP7_75t_L g1316 ( .A(n_393), .Y(n_1316) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g677 ( .A(n_394), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .B1(n_400), .B2(n_403), .Y(n_395) );
INVx1_ASAP7_75t_L g587 ( .A(n_396), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_396), .A2(n_741), .B1(n_742), .B2(n_743), .Y(n_740) );
BUFx3_ASAP7_75t_L g767 ( .A(n_396), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g870 ( .A1(n_396), .A2(n_400), .B1(n_863), .B2(n_871), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_396), .A2(n_891), .B1(n_1110), .B2(n_1112), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_396), .A2(n_682), .B1(n_1166), .B2(n_1167), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_396), .A2(n_743), .B1(n_1242), .B2(n_1243), .Y(n_1241) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
OR2x2_ASAP7_75t_L g409 ( .A(n_397), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g591 ( .A(n_397), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g680 ( .A(n_397), .B(n_398), .Y(n_680) );
O2A1O1Ixp33_ASAP7_75t_L g1646 ( .A1(n_397), .A2(n_1316), .B(n_1647), .C(n_1648), .Y(n_1646) );
INVx1_ASAP7_75t_L g1652 ( .A(n_397), .Y(n_1652) );
INVx1_ASAP7_75t_L g1728 ( .A(n_398), .Y(n_1728) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_399), .A2(n_449), .B1(n_453), .B2(n_454), .Y(n_448) );
INVx2_ASAP7_75t_L g588 ( .A(n_400), .Y(n_588) );
INVx2_ASAP7_75t_L g683 ( .A(n_400), .Y(n_683) );
BUFx3_ASAP7_75t_L g743 ( .A(n_400), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_400), .A2(n_1027), .B1(n_1199), .B2(n_1201), .Y(n_1213) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_406), .Y(n_771) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g1124 ( .A(n_408), .Y(n_1124) );
INVxp67_ASAP7_75t_SL g1169 ( .A(n_408), .Y(n_1169) );
INVx1_ASAP7_75t_L g1402 ( .A(n_408), .Y(n_1402) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g598 ( .A(n_409), .Y(n_598) );
BUFx2_ASAP7_75t_L g773 ( .A(n_409), .Y(n_773) );
INVx8_ASAP7_75t_L g487 ( .A(n_410), .Y(n_487) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_410), .Y(n_1100) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI31xp33_ASAP7_75t_L g866 ( .A1(n_413), .A2(n_867), .A3(n_869), .B(n_872), .Y(n_866) );
BUFx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g599 ( .A(n_414), .Y(n_599) );
BUFx2_ASAP7_75t_L g688 ( .A(n_414), .Y(n_688) );
OAI31xp33_ASAP7_75t_L g736 ( .A1(n_414), .A2(n_737), .A3(n_739), .B(n_744), .Y(n_736) );
BUFx3_ASAP7_75t_L g897 ( .A(n_414), .Y(n_897) );
OAI31xp33_ASAP7_75t_L g1238 ( .A1(n_414), .A2(n_1239), .A3(n_1240), .B(n_1244), .Y(n_1238) );
OAI21xp5_ASAP7_75t_L g1313 ( .A1(n_414), .A2(n_1314), .B(n_1322), .Y(n_1313) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g472 ( .A(n_417), .Y(n_472) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI31xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_436), .A3(n_456), .B(n_466), .Y(n_419) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_SL g626 ( .A(n_422), .Y(n_626) );
BUFx2_ASAP7_75t_L g777 ( .A(n_422), .Y(n_777) );
BUFx2_ASAP7_75t_L g939 ( .A(n_422), .Y(n_939) );
OR2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_426), .Y(n_422) );
AND2x4_ASAP7_75t_L g461 ( .A(n_423), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g703 ( .A(n_423), .B(n_462), .Y(n_703) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x6_ASAP7_75t_L g432 ( .A(n_424), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g445 ( .A(n_424), .B(n_446), .Y(n_445) );
OR2x4_ASAP7_75t_L g459 ( .A(n_424), .B(n_426), .Y(n_459) );
NAND3x1_ASAP7_75t_L g540 ( .A(n_424), .B(n_541), .C(n_543), .Y(n_540) );
NAND2x1p5_ASAP7_75t_L g655 ( .A(n_424), .B(n_543), .Y(n_655) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx3_ASAP7_75t_L g451 ( .A(n_425), .Y(n_451) );
NAND2xp33_ASAP7_75t_SL g519 ( .A(n_425), .B(n_469), .Y(n_519) );
INVx2_ASAP7_75t_L g523 ( .A(n_426), .Y(n_523) );
BUFx4f_ASAP7_75t_L g640 ( .A(n_426), .Y(n_640) );
BUFx3_ASAP7_75t_L g816 ( .A(n_426), .Y(n_816) );
BUFx3_ASAP7_75t_L g826 ( .A(n_426), .Y(n_826) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_427), .B(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_427), .Y(n_443) );
AND2x4_ASAP7_75t_L g446 ( .A(n_427), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
INVx1_ASAP7_75t_L g953 ( .A(n_428), .Y(n_953) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g464 ( .A(n_429), .Y(n_464) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g627 ( .A(n_432), .Y(n_627) );
INVx1_ASAP7_75t_L g886 ( .A(n_432), .Y(n_886) );
BUFx3_ASAP7_75t_L g1178 ( .A(n_432), .Y(n_1178) );
INVx1_ASAP7_75t_L g532 ( .A(n_433), .Y(n_532) );
BUFx3_ASAP7_75t_L g821 ( .A(n_433), .Y(n_821) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g537 ( .A(n_434), .Y(n_537) );
INVx1_ASAP7_75t_L g442 ( .A(n_435), .Y(n_442) );
INVx2_ASAP7_75t_L g447 ( .A(n_435), .Y(n_447) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI22xp33_ASAP7_75t_L g544 ( .A1(n_438), .A2(n_484), .B1(n_504), .B2(n_521), .Y(n_544) );
OAI22xp33_ASAP7_75t_L g1153 ( .A1(n_438), .A2(n_1137), .B1(n_1146), .B2(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g780 ( .A(n_439), .Y(n_780) );
INVx1_ASAP7_75t_L g846 ( .A(n_439), .Y(n_846) );
INVx1_ASAP7_75t_L g942 ( .A(n_439), .Y(n_942) );
INVx1_ASAP7_75t_L g1174 ( .A(n_439), .Y(n_1174) );
INVx2_ASAP7_75t_L g1286 ( .A(n_439), .Y(n_1286) );
INVx4_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_440), .Y(n_556) );
INVx3_ASAP7_75t_L g712 ( .A(n_440), .Y(n_712) );
HB1xp67_ASAP7_75t_L g1345 ( .A(n_440), .Y(n_1345) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g526 ( .A(n_441), .Y(n_526) );
BUFx3_ASAP7_75t_L g575 ( .A(n_441), .Y(n_575) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
BUFx2_ASAP7_75t_L g455 ( .A(n_442), .Y(n_455) );
BUFx2_ASAP7_75t_L g452 ( .A(n_443), .Y(n_452) );
INVx2_ASAP7_75t_L g697 ( .A(n_443), .Y(n_697) );
AND2x4_ASAP7_75t_L g962 ( .A(n_443), .B(n_695), .Y(n_962) );
NAND3xp33_ASAP7_75t_SL g1197 ( .A(n_444), .B(n_1198), .C(n_1200), .Y(n_1197) );
NAND3xp33_ASAP7_75t_SL g1247 ( .A(n_444), .B(n_1248), .C(n_1250), .Y(n_1247) );
CKINVDCx8_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
AOI211xp5_ASAP7_75t_L g617 ( .A1(n_445), .A2(n_618), .B(n_619), .C(n_620), .Y(n_617) );
CKINVDCx8_ASAP7_75t_R g700 ( .A(n_445), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g937 ( .A(n_445), .B(n_938), .C(n_941), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_445), .B(n_1108), .Y(n_1107) );
NOR3xp33_ASAP7_75t_L g1674 ( .A(n_445), .B(n_1675), .C(n_1678), .Y(n_1674) );
OAI31xp33_ASAP7_75t_L g1745 ( .A1(n_445), .A2(n_704), .A3(n_1746), .B(n_1757), .Y(n_1745) );
BUFx3_ASAP7_75t_L g619 ( .A(n_446), .Y(n_619) );
INVx2_ASAP7_75t_L g955 ( .A(n_446), .Y(n_955) );
BUFx2_ASAP7_75t_L g965 ( .A(n_446), .Y(n_965) );
BUFx2_ASAP7_75t_L g1113 ( .A(n_446), .Y(n_1113) );
BUFx2_ASAP7_75t_L g1249 ( .A(n_446), .Y(n_1249) );
BUFx2_ASAP7_75t_L g1308 ( .A(n_446), .Y(n_1308) );
INVx1_ASAP7_75t_L g695 ( .A(n_447), .Y(n_695) );
INVx1_ASAP7_75t_L g621 ( .A(n_449), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_449), .A2(n_454), .B1(n_1166), .B2(n_1176), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1407 ( .A1(n_449), .A2(n_454), .B1(n_1397), .B2(n_1400), .Y(n_1407) );
AOI22xp5_ASAP7_75t_L g1754 ( .A1(n_449), .A2(n_454), .B1(n_1755), .B2(n_1756), .Y(n_1754) );
AND2x4_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
AND2x4_ASAP7_75t_L g454 ( .A(n_450), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g698 ( .A(n_450), .B(n_455), .Y(n_698) );
AND2x4_ASAP7_75t_L g754 ( .A(n_450), .B(n_452), .Y(n_754) );
AND2x2_ASAP7_75t_L g783 ( .A(n_450), .B(n_452), .Y(n_783) );
A2O1A1Ixp33_ASAP7_75t_L g1746 ( .A1(n_450), .A2(n_1747), .B(n_1750), .C(n_1754), .Y(n_1746) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g693 ( .A(n_451), .B(n_694), .Y(n_693) );
AND3x4_ASAP7_75t_L g945 ( .A(n_451), .B(n_469), .C(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g622 ( .A(n_454), .Y(n_622) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_454), .Y(n_785) );
AOI222xp33_ASAP7_75t_L g1109 ( .A1(n_454), .A2(n_754), .B1(n_1110), .B2(n_1111), .C1(n_1112), .C2(n_1113), .Y(n_1109) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g1679 ( .A1(n_458), .A2(n_703), .B1(n_1651), .B2(n_1680), .Y(n_1679) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_SL g624 ( .A(n_459), .Y(n_624) );
INVx2_ASAP7_75t_SL g788 ( .A(n_459), .Y(n_788) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_459), .Y(n_856) );
INVx1_ASAP7_75t_L g1119 ( .A(n_459), .Y(n_1119) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_461), .A2(n_579), .B1(n_580), .B2(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g789 ( .A(n_461), .Y(n_789) );
INVx1_ASAP7_75t_L g857 ( .A(n_461), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_461), .A2(n_624), .B1(n_935), .B2(n_936), .Y(n_934) );
INVx1_ASAP7_75t_L g1405 ( .A(n_461), .Y(n_1405) );
INVx2_ASAP7_75t_L g716 ( .A(n_462), .Y(n_716) );
BUFx6f_ASAP7_75t_L g820 ( .A(n_462), .Y(n_820) );
INVx1_ASAP7_75t_L g842 ( .A(n_462), .Y(n_842) );
INVx2_ASAP7_75t_L g1159 ( .A(n_462), .Y(n_1159) );
INVx2_ASAP7_75t_L g1349 ( .A(n_462), .Y(n_1349) );
BUFx6f_ASAP7_75t_L g1685 ( .A(n_462), .Y(n_1685) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_463), .Y(n_529) );
BUFx8_ASAP7_75t_L g564 ( .A(n_463), .Y(n_564) );
INVx2_ASAP7_75t_L g959 ( .A(n_463), .Y(n_959) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
AND2x4_ASAP7_75t_L g952 ( .A(n_465), .B(n_953), .Y(n_952) );
OAI31xp33_ASAP7_75t_L g854 ( .A1(n_466), .A2(n_855), .A3(n_858), .B(n_865), .Y(n_854) );
OAI31xp33_ASAP7_75t_L g1171 ( .A1(n_466), .A2(n_1172), .A3(n_1173), .B(n_1177), .Y(n_1171) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .Y(n_466) );
AND2x4_ASAP7_75t_L g629 ( .A(n_467), .B(n_470), .Y(n_629) );
AND2x2_ASAP7_75t_L g704 ( .A(n_467), .B(n_470), .Y(n_704) );
AND2x2_ASAP7_75t_SL g790 ( .A(n_467), .B(n_470), .Y(n_790) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_467), .B(n_470), .Y(n_1204) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g509 ( .A(n_472), .Y(n_509) );
OR2x2_ASAP7_75t_L g518 ( .A(n_472), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_SL g670 ( .A(n_472), .B(n_507), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_516), .Y(n_473) );
OAI33xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_481), .A3(n_488), .B1(n_498), .B2(n_505), .B3(n_510), .Y(n_474) );
OAI33xp33_ASAP7_75t_L g848 ( .A1(n_475), .A2(n_806), .A3(n_849), .B1(n_851), .B2(n_852), .B3(n_853), .Y(n_848) );
INVx1_ASAP7_75t_L g971 ( .A(n_475), .Y(n_971) );
OAI33xp33_ASAP7_75t_L g1327 ( .A1(n_475), .A2(n_806), .A3(n_1328), .B1(n_1331), .B2(n_1334), .B3(n_1340), .Y(n_1327) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI33xp33_ASAP7_75t_L g726 ( .A1(n_476), .A2(n_669), .A3(n_727), .B1(n_731), .B2(n_733), .B3(n_735), .Y(n_726) );
OAI33xp33_ASAP7_75t_L g1041 ( .A1(n_476), .A2(n_1023), .A3(n_1042), .B1(n_1046), .B2(n_1049), .B3(n_1053), .Y(n_1041) );
OAI33xp33_ASAP7_75t_L g1254 ( .A1(n_476), .A2(n_1023), .A3(n_1255), .B1(n_1258), .B2(n_1261), .B3(n_1264), .Y(n_1254) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g601 ( .A(n_477), .Y(n_601) );
INVx4_ASAP7_75t_L g793 ( .A(n_477), .Y(n_793) );
INVx2_ASAP7_75t_L g917 ( .A(n_477), .Y(n_917) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
OR2x2_ASAP7_75t_L g654 ( .A(n_478), .B(n_655), .Y(n_654) );
OR2x6_ASAP7_75t_L g1091 ( .A(n_478), .B(n_655), .Y(n_1091) );
INVx1_ASAP7_75t_L g1671 ( .A(n_478), .Y(n_1671) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g946 ( .A(n_479), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B1(n_484), .B2(n_485), .Y(n_481) );
OAI22xp33_ASAP7_75t_L g520 ( .A1(n_482), .A2(n_501), .B1(n_521), .B2(n_524), .Y(n_520) );
OAI22xp33_ASAP7_75t_L g1099 ( .A1(n_483), .A2(n_1082), .B1(n_1093), .B2(n_1100), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_483), .A2(n_1044), .B1(n_1086), .B2(n_1090), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1657 ( .A1(n_483), .A2(n_485), .B1(n_1658), .B2(n_1659), .Y(n_1657) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_485), .A2(n_511), .B1(n_514), .B2(n_515), .Y(n_510) );
INVx5_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx6_ASAP7_75t_L g798 ( .A(n_486), .Y(n_798) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx4_ASAP7_75t_L g659 ( .A(n_487), .Y(n_659) );
INVx2_ASAP7_75t_L g730 ( .A(n_487), .Y(n_730) );
INVx1_ASAP7_75t_L g811 ( .A(n_487), .Y(n_811) );
INVx1_ASAP7_75t_L g850 ( .A(n_487), .Y(n_850) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_487), .Y(n_1044) );
INVx2_ASAP7_75t_L g1150 ( .A(n_487), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B1(n_495), .B2(n_496), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_489), .A2(n_514), .B1(n_528), .B2(n_530), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_490), .A2(n_732), .B1(n_837), .B2(n_841), .Y(n_851) );
INVx4_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g803 ( .A(n_491), .Y(n_803) );
INVx2_ASAP7_75t_L g1142 ( .A(n_491), .Y(n_1142) );
INVx4_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx3_ASAP7_75t_L g500 ( .A(n_493), .Y(n_500) );
INVx2_ASAP7_75t_L g604 ( .A(n_493), .Y(n_604) );
INVx1_ASAP7_75t_L g662 ( .A(n_493), .Y(n_662) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_493), .Y(n_1021) );
AND2x2_ASAP7_75t_L g593 ( .A(n_494), .B(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g1731 ( .A(n_494), .Y(n_1731) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_495), .A2(n_515), .B1(n_534), .B2(n_535), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_496), .A2(n_603), .B1(n_800), .B2(n_801), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g1144 ( .A1(n_496), .A2(n_1145), .B1(n_1146), .B2(n_1147), .Y(n_1144) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_496), .A2(n_803), .B1(n_1332), .B2(n_1333), .Y(n_1331) );
INVx5_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI22xp33_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_501), .B1(n_502), .B2(n_504), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g613 ( .A(n_500), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_500), .A2(n_713), .B1(n_725), .B2(n_734), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g1301 ( .A1(n_500), .A2(n_673), .B1(n_1289), .B2(n_1294), .Y(n_1301) );
OAI22xp5_ASAP7_75t_L g1383 ( .A1(n_500), .A2(n_732), .B1(n_1384), .B2(n_1385), .Y(n_1383) );
OAI211xp5_ASAP7_75t_SL g1663 ( .A1(n_502), .A2(n_1664), .B(n_1665), .C(n_1668), .Y(n_1663) );
OAI211xp5_ASAP7_75t_SL g1713 ( .A1(n_502), .A2(n_1714), .B(n_1715), .C(n_1717), .Y(n_1713) );
OAI211xp5_ASAP7_75t_SL g1718 ( .A1(n_502), .A2(n_1719), .B(n_1720), .C(n_1722), .Y(n_1718) );
BUFx4f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx4_ASAP7_75t_L g664 ( .A(n_503), .Y(n_664) );
BUFx4f_ASAP7_75t_L g673 ( .A(n_503), .Y(n_673) );
BUFx4f_ASAP7_75t_L g732 ( .A(n_503), .Y(n_732) );
BUFx4f_ASAP7_75t_L g764 ( .A(n_503), .Y(n_764) );
BUFx6f_ASAP7_75t_L g1051 ( .A(n_503), .Y(n_1051) );
OAI22xp5_ASAP7_75t_SL g600 ( .A1(n_505), .A2(n_601), .B1(n_602), .B2(n_611), .Y(n_600) );
OAI33xp33_ASAP7_75t_L g916 ( .A1(n_505), .A2(n_917), .A3(n_918), .B1(n_922), .B2(n_926), .B3(n_928), .Y(n_916) );
OAI33xp33_ASAP7_75t_L g1135 ( .A1(n_505), .A2(n_793), .A3(n_1136), .B1(n_1140), .B2(n_1144), .B3(n_1148), .Y(n_1135) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g806 ( .A(n_506), .Y(n_806) );
AOI33xp33_ASAP7_75t_L g970 ( .A1(n_506), .A2(n_971), .A3(n_972), .B1(n_976), .B2(n_983), .B3(n_984), .Y(n_970) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
OAI221xp5_ASAP7_75t_L g1660 ( .A1(n_507), .A2(n_923), .B1(n_1102), .B2(n_1661), .C(n_1662), .Y(n_1660) );
INVx4_ASAP7_75t_L g1716 ( .A(n_507), .Y(n_1716) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g849 ( .A1(n_511), .A2(n_833), .B1(n_845), .B2(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g808 ( .A(n_512), .Y(n_808) );
INVx3_ASAP7_75t_L g1138 ( .A(n_512), .Y(n_1138) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g658 ( .A(n_513), .Y(n_658) );
INVx3_ASAP7_75t_L g921 ( .A(n_513), .Y(n_921) );
OAI33xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_520), .A3(n_527), .B1(n_533), .B2(n_538), .B3(n_544), .Y(n_516) );
BUFx4f_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx4f_ASAP7_75t_L g549 ( .A(n_518), .Y(n_549) );
BUFx8_ASAP7_75t_L g814 ( .A(n_518), .Y(n_814) );
BUFx2_ASAP7_75t_L g900 ( .A(n_518), .Y(n_900) );
BUFx4f_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g1081 ( .A1(n_522), .A2(n_711), .B1(n_1082), .B2(n_1083), .Y(n_1081) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_SL g554 ( .A(n_523), .Y(n_554) );
OAI22xp33_ASAP7_75t_L g913 ( .A1(n_524), .A2(n_816), .B1(n_914), .B2(n_915), .Y(n_913) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g860 ( .A(n_526), .Y(n_860) );
INVx1_ASAP7_75t_L g1363 ( .A(n_526), .Y(n_1363) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_528), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_528), .A2(n_561), .B1(n_1048), .B2(n_1055), .Y(n_1059) );
INVx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx5_ASAP7_75t_L g534 ( .A(n_529), .Y(n_534) );
INVx2_ASAP7_75t_SL g559 ( .A(n_529), .Y(n_559) );
INVx3_ASAP7_75t_L g648 ( .A(n_529), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g1750 ( .A1(n_529), .A2(n_1751), .B1(n_1752), .B2(n_1753), .Y(n_1750) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_530), .A2(n_837), .B1(n_838), .B2(n_839), .Y(n_836) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g645 ( .A(n_532), .Y(n_645) );
BUFx3_ASAP7_75t_L g838 ( .A(n_534), .Y(n_838) );
OAI22xp33_ASAP7_75t_SL g1388 ( .A1(n_534), .A2(n_645), .B1(n_1373), .B2(n_1381), .Y(n_1388) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_535), .A2(n_841), .B1(n_842), .B2(n_843), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_535), .A2(n_838), .B1(n_906), .B2(n_907), .Y(n_905) );
OAI22xp33_ASAP7_75t_SL g1158 ( .A1(n_535), .A2(n_1143), .B1(n_1151), .B2(n_1159), .Y(n_1158) );
OAI221xp5_ASAP7_75t_L g1689 ( .A1(n_535), .A2(n_1290), .B1(n_1659), .B2(n_1664), .C(n_1690), .Y(n_1689) );
OAI221xp5_ASAP7_75t_L g1735 ( .A1(n_535), .A2(n_1684), .B1(n_1736), .B2(n_1737), .C(n_1738), .Y(n_1735) );
OAI221xp5_ASAP7_75t_L g1741 ( .A1(n_535), .A2(n_1157), .B1(n_1719), .B2(n_1742), .C(n_1743), .Y(n_1741) );
CKINVDCx8_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
INVx3_ASAP7_75t_L g561 ( .A(n_536), .Y(n_561) );
INVx3_ASAP7_75t_L g718 ( .A(n_536), .Y(n_718) );
INVx3_ASAP7_75t_L g722 ( .A(n_536), .Y(n_722) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g567 ( .A(n_537), .Y(n_567) );
OAI33xp33_ASAP7_75t_L g813 ( .A1(n_538), .A2(n_814), .A3(n_815), .B1(n_818), .B2(n_822), .B3(n_823), .Y(n_813) );
OAI33xp33_ASAP7_75t_L g831 ( .A1(n_538), .A2(n_814), .A3(n_832), .B1(n_836), .B2(n_840), .B3(n_844), .Y(n_831) );
OAI33xp33_ASAP7_75t_L g899 ( .A1(n_538), .A2(n_900), .A3(n_901), .B1(n_905), .B2(n_908), .B3(n_913), .Y(n_899) );
INVx1_ASAP7_75t_L g969 ( .A(n_538), .Y(n_969) );
OAI33xp33_ASAP7_75t_L g1343 ( .A1(n_538), .A2(n_900), .A3(n_1344), .B1(n_1346), .B2(n_1348), .B3(n_1350), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g1681 ( .A1(n_538), .A2(n_900), .B1(n_1682), .B2(n_1689), .Y(n_1681) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g1160 ( .A(n_539), .Y(n_1160) );
INVx2_ASAP7_75t_L g1744 ( .A(n_539), .Y(n_1744) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx3_ASAP7_75t_L g571 ( .A(n_540), .Y(n_571) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g631 ( .A(n_545), .Y(n_631) );
NOR4xp25_ASAP7_75t_L g546 ( .A(n_547), .B(n_577), .C(n_600), .D(n_616), .Y(n_546) );
OAI33xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_550), .A3(n_557), .B1(n_562), .B2(n_569), .B3(n_572), .Y(n_547) );
OAI22xp33_ASAP7_75t_L g1734 ( .A1(n_548), .A2(n_1735), .B1(n_1741), .B2(n_1744), .Y(n_1734) );
BUFx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI33xp33_ASAP7_75t_L g637 ( .A1(n_549), .A2(n_638), .A3(n_642), .B1(n_647), .B2(n_651), .B3(n_654), .Y(n_637) );
OAI33xp33_ASAP7_75t_L g708 ( .A1(n_549), .A2(n_654), .A3(n_709), .B1(n_714), .B2(n_719), .B3(n_723), .Y(n_708) );
OAI33xp33_ASAP7_75t_L g1001 ( .A1(n_549), .A2(n_654), .A3(n_1002), .B1(n_1005), .B2(n_1008), .B3(n_1013), .Y(n_1001) );
OAI33xp33_ASAP7_75t_L g1056 ( .A1(n_549), .A2(n_654), .A3(n_1057), .B1(n_1058), .B2(n_1059), .B3(n_1060), .Y(n_1056) );
OAI33xp33_ASAP7_75t_L g1267 ( .A1(n_549), .A2(n_654), .A3(n_1268), .B1(n_1269), .B2(n_1270), .B3(n_1271), .Y(n_1267) );
OAI22xp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B1(n_555), .B2(n_556), .Y(n_550) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_554), .A2(n_573), .B1(n_574), .B2(n_576), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g1013 ( .A1(n_554), .A2(n_575), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
OAI22xp33_ASAP7_75t_L g1057 ( .A1(n_554), .A2(n_556), .B1(n_1043), .B2(n_1050), .Y(n_1057) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_554), .A2(n_575), .B1(n_1045), .B2(n_1052), .Y(n_1060) );
OAI22xp33_ASAP7_75t_L g1268 ( .A1(n_554), .A2(n_575), .B1(n_1256), .B2(n_1262), .Y(n_1268) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_556), .A2(n_639), .B1(n_640), .B2(n_641), .Y(n_638) );
OAI22xp33_ASAP7_75t_L g1092 ( .A1(n_556), .A2(n_816), .B1(n_1093), .B2(n_1094), .Y(n_1092) );
OAI22xp33_ASAP7_75t_L g1296 ( .A1(n_556), .A2(n_640), .B1(n_1297), .B2(n_1298), .Y(n_1296) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_560), .B2(n_561), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g1292 ( .A1(n_561), .A2(n_1293), .B1(n_1294), .B2(n_1295), .Y(n_1292) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .B1(n_566), .B2(n_568), .Y(n_562) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_SL g644 ( .A(n_564), .Y(n_644) );
INVx3_ASAP7_75t_L g1088 ( .A(n_564), .Y(n_1088) );
INVx3_ASAP7_75t_L g1293 ( .A(n_564), .Y(n_1293) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_566), .A2(n_648), .B1(n_649), .B2(n_650), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_566), .A2(n_958), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_566), .A2(n_1088), .B1(n_1089), .B2(n_1090), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1288 ( .A1(n_566), .A2(n_1289), .B1(n_1290), .B2(n_1291), .Y(n_1288) );
BUFx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g1391 ( .A(n_567), .Y(n_1391) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g651 ( .A1(n_575), .A2(n_640), .B1(n_652), .B2(n_653), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_575), .A2(n_640), .B1(n_724), .B2(n_725), .Y(n_723) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_575), .Y(n_817) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_575), .Y(n_835) );
OAI22xp33_ASAP7_75t_L g1392 ( .A1(n_575), .A2(n_640), .B1(n_1377), .B2(n_1385), .Y(n_1392) );
AOI31xp33_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_581), .A3(n_589), .B(n_599), .Y(n_577) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g891 ( .A(n_588), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_595), .B2(n_596), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_590), .A2(n_595), .B1(n_626), .B2(n_627), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_591), .A2(n_1319), .B1(n_1320), .B2(n_1321), .Y(n_1318) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_592), .Y(n_615) );
INVx3_ASAP7_75t_L g1232 ( .A(n_592), .Y(n_1232) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx3_ASAP7_75t_L g607 ( .A(n_593), .Y(n_607) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g1654 ( .A(n_598), .B(n_1655), .Y(n_1654) );
AO21x1_ASAP7_75t_L g988 ( .A1(n_599), .A2(n_989), .B(n_990), .Y(n_988) );
AO21x1_ASAP7_75t_L g1205 ( .A1(n_599), .A2(n_1206), .B(n_1210), .Y(n_1205) );
OAI33xp33_ASAP7_75t_L g656 ( .A1(n_601), .A2(n_657), .A3(n_660), .B1(n_665), .B2(n_666), .B3(n_669), .Y(n_656) );
OAI33xp33_ASAP7_75t_L g1016 ( .A1(n_601), .A2(n_1017), .A3(n_1018), .B1(n_1020), .B2(n_1022), .B3(n_1023), .Y(n_1016) );
OAI33xp33_ASAP7_75t_L g1299 ( .A1(n_601), .A2(n_669), .A3(n_1300), .B1(n_1301), .B2(n_1302), .B3(n_1303), .Y(n_1299) );
INVx1_ASAP7_75t_L g1336 ( .A(n_603), .Y(n_1336) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx2_ASAP7_75t_L g924 ( .A(n_604), .Y(n_924) );
INVx2_ASAP7_75t_L g1019 ( .A(n_604), .Y(n_1019) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g973 ( .A(n_607), .Y(n_973) );
INVx2_ASAP7_75t_SL g985 ( .A(n_607), .Y(n_985) );
INVx2_ASAP7_75t_L g1224 ( .A(n_607), .Y(n_1224) );
INVx2_ASAP7_75t_L g1669 ( .A(n_607), .Y(n_1669) );
BUFx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx3_ASAP7_75t_L g975 ( .A(n_610), .Y(n_975) );
INVx2_ASAP7_75t_L g987 ( .A(n_610), .Y(n_987) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
A2O1A1Ixp33_ASAP7_75t_SL g1723 ( .A1(n_615), .A2(n_1724), .B(n_1725), .C(n_1732), .Y(n_1723) );
AOI31xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_623), .A3(n_625), .B(n_628), .Y(n_616) );
INVx1_ASAP7_75t_L g1191 ( .A(n_619), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1747 ( .A1(n_619), .A2(n_1724), .B1(n_1748), .B2(n_1749), .Y(n_1747) );
AOI22xp5_ASAP7_75t_L g1117 ( .A1(n_626), .A2(n_1118), .B1(n_1119), .B2(n_1120), .Y(n_1117) );
INVx1_ASAP7_75t_L g778 ( .A(n_627), .Y(n_778) );
INVx2_ASAP7_75t_L g940 ( .A(n_627), .Y(n_940) );
AO21x1_ASAP7_75t_L g933 ( .A1(n_628), .A2(n_934), .B(n_937), .Y(n_933) );
AOI31xp33_ASAP7_75t_L g1106 ( .A1(n_628), .A2(n_1107), .A3(n_1114), .B(n_1117), .Y(n_1106) );
CKINVDCx14_ASAP7_75t_R g628 ( .A(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
XNOR2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_705), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_671), .C(n_689), .Y(n_635) );
NOR2xp33_ASAP7_75t_SL g636 ( .A(n_637), .B(n_656), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_639), .A2(n_652), .B1(n_658), .B2(n_659), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_640), .A2(n_710), .B1(n_711), .B2(n_713), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_640), .A2(n_711), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1271 ( .A1(n_640), .A2(n_846), .B1(n_1257), .B2(n_1263), .Y(n_1271) );
OAI22xp33_ASAP7_75t_L g1284 ( .A1(n_640), .A2(n_1285), .B1(n_1286), .B2(n_1287), .Y(n_1284) );
OAI22xp33_ASAP7_75t_L g1387 ( .A1(n_640), .A2(n_711), .B1(n_1376), .B2(n_1384), .Y(n_1387) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_641), .A2(n_653), .B1(n_661), .B2(n_663), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B1(n_645), .B2(n_646), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_643), .A2(n_649), .B1(n_661), .B2(n_663), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_645), .A2(n_1009), .B1(n_1010), .B2(n_1012), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_646), .A2(n_650), .B1(n_659), .B2(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g910 ( .A(n_648), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_648), .A2(n_718), .B1(n_1259), .B2(n_1265), .Y(n_1269) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_658), .A2(n_729), .B1(n_1003), .B2(n_1014), .Y(n_1017) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_658), .A2(n_659), .B1(n_1007), .B2(n_1012), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_658), .A2(n_1043), .B1(n_1044), .B2(n_1045), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_658), .A2(n_729), .B1(n_1054), .B2(n_1055), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_658), .A2(n_729), .B1(n_1256), .B2(n_1257), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_658), .A2(n_1044), .B1(n_1265), .B2(n_1266), .Y(n_1264) );
OAI22xp33_ASAP7_75t_L g1375 ( .A1(n_658), .A2(n_811), .B1(n_1376), .B2(n_1377), .Y(n_1375) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_659), .A2(n_717), .B1(n_721), .B2(n_728), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g1300 ( .A1(n_659), .A2(n_728), .B1(n_1285), .B2(n_1297), .Y(n_1300) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_661), .A2(n_715), .B1(n_720), .B2(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g1372 ( .A1(n_661), .A2(n_1051), .B1(n_1373), .B2(n_1374), .Y(n_1372) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g1145 ( .A(n_662), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_663), .A2(n_1006), .B1(n_1009), .B2(n_1019), .Y(n_1018) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g734 ( .A(n_664), .Y(n_734) );
INVx2_ASAP7_75t_L g925 ( .A(n_664), .Y(n_925) );
INVx1_ASAP7_75t_L g927 ( .A(n_664), .Y(n_927) );
INVx1_ASAP7_75t_L g1102 ( .A(n_664), .Y(n_1102) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g1023 ( .A(n_670), .Y(n_1023) );
AOI33xp33_ASAP7_75t_L g1222 ( .A1(n_670), .A2(n_1098), .A3(n_1223), .B1(n_1225), .B2(n_1229), .B3(n_1230), .Y(n_1222) );
OAI31xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_684), .A3(n_687), .B(n_688), .Y(n_671) );
NAND3xp33_ASAP7_75t_SL g1314 ( .A(n_674), .B(n_1315), .C(n_1318), .Y(n_1314) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g1217 ( .A(n_675), .Y(n_1217) );
INVx1_ASAP7_75t_L g1216 ( .A(n_676), .Y(n_1216) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
BUFx2_ASAP7_75t_L g982 ( .A(n_677), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_681), .B2(n_682), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_680), .A2(n_882), .B1(n_891), .B2(n_892), .Y(n_890) );
AOI222xp33_ASAP7_75t_L g1315 ( .A1(n_680), .A2(n_743), .B1(n_1310), .B2(n_1311), .C1(n_1316), .C2(n_1317), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1396 ( .A1(n_680), .A2(n_743), .B1(n_1397), .B2(n_1398), .Y(n_1396) );
AOI32xp33_ASAP7_75t_L g692 ( .A1(n_681), .A2(n_693), .A3(n_696), .B1(n_698), .B2(n_699), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g1026 ( .A1(n_682), .A2(n_1027), .B1(n_1028), .B2(n_1029), .Y(n_1026) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g1208 ( .A(n_685), .Y(n_1208) );
BUFx3_ASAP7_75t_L g728 ( .A(n_686), .Y(n_728) );
BUFx3_ASAP7_75t_L g796 ( .A(n_686), .Y(n_796) );
BUFx6f_ASAP7_75t_L g1304 ( .A(n_686), .Y(n_1304) );
OAI31xp33_ASAP7_75t_L g760 ( .A1(n_688), .A2(n_761), .A3(n_770), .B(n_774), .Y(n_760) );
OAI31xp33_ASAP7_75t_L g1024 ( .A1(n_688), .A2(n_1025), .A3(n_1030), .B(n_1031), .Y(n_1024) );
OAI31xp33_ASAP7_75t_L g1061 ( .A1(n_688), .A2(n_1062), .A3(n_1066), .B(n_1067), .Y(n_1061) );
INVx1_ASAP7_75t_L g1129 ( .A(n_688), .Y(n_1129) );
OAI31xp33_ASAP7_75t_L g1163 ( .A1(n_688), .A2(n_1164), .A3(n_1168), .B(n_1170), .Y(n_1163) );
OAI31xp33_ASAP7_75t_L g1393 ( .A1(n_688), .A2(n_1394), .A3(n_1395), .B(n_1401), .Y(n_1393) );
OAI31xp33_ASAP7_75t_SL g689 ( .A1(n_690), .A2(n_691), .A3(n_701), .B(n_704), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_693), .A2(n_741), .B1(n_753), .B2(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_L g751 ( .A(n_698), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_698), .A2(n_754), .B1(n_1028), .B2(n_1036), .Y(n_1035) );
AOI22xp33_ASAP7_75t_SL g1071 ( .A1(n_698), .A2(n_754), .B1(n_1064), .B2(n_1072), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_698), .A2(n_754), .B1(n_1201), .B2(n_1202), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1250 ( .A1(n_698), .A2(n_754), .B1(n_1242), .B2(n_1251), .Y(n_1250) );
AOI222xp33_ASAP7_75t_L g1307 ( .A1(n_698), .A2(n_754), .B1(n_1308), .B2(n_1309), .C1(n_1310), .C2(n_1311), .Y(n_1307) );
INVxp67_ASAP7_75t_L g1677 ( .A(n_698), .Y(n_1677) );
NAND3xp33_ASAP7_75t_L g1406 ( .A(n_700), .B(n_1407), .C(n_1408), .Y(n_1406) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_703), .A2(n_886), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
OAI31xp33_ASAP7_75t_SL g747 ( .A1(n_704), .A2(n_748), .A3(n_749), .B(n_750), .Y(n_747) );
OAI31xp33_ASAP7_75t_SL g1032 ( .A1(n_704), .A2(n_1033), .A3(n_1034), .B(n_1037), .Y(n_1032) );
OAI31xp33_ASAP7_75t_SL g1068 ( .A1(n_704), .A2(n_1069), .A3(n_1070), .B(n_1073), .Y(n_1068) );
OAI21xp5_ASAP7_75t_L g1305 ( .A1(n_704), .A2(n_1306), .B(n_1312), .Y(n_1305) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_736), .C(n_747), .Y(n_706) );
NOR2xp33_ASAP7_75t_SL g707 ( .A(n_708), .B(n_726), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_710), .A2(n_724), .B1(n_728), .B2(n_729), .Y(n_727) );
INVx3_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g904 ( .A(n_712), .Y(n_904) );
INVx2_ASAP7_75t_L g1162 ( .A(n_712), .Y(n_1162) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_716), .A2(n_801), .B1(n_812), .B2(n_821), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_716), .A2(n_718), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_716), .A2(n_718), .B1(n_1047), .B2(n_1054), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g1270 ( .A1(n_716), .A2(n_722), .B1(n_1260), .B2(n_1266), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_728), .A2(n_729), .B1(n_1381), .B2(n_1382), .Y(n_1380) );
OAI22xp5_ASAP7_75t_L g1303 ( .A1(n_729), .A2(n_1291), .B1(n_1295), .B2(n_1304), .Y(n_1303) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g1261 ( .A1(n_732), .A2(n_1019), .B1(n_1262), .B2(n_1263), .Y(n_1261) );
INVx1_ASAP7_75t_L g1321 ( .A(n_738), .Y(n_1321) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_743), .A2(n_767), .B1(n_768), .B2(n_769), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_743), .A2(n_1027), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_743), .A2(n_767), .B1(n_1355), .B2(n_1356), .Y(n_1354) );
INVx1_ASAP7_75t_L g1676 ( .A(n_754), .Y(n_1676) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B1(n_827), .B2(n_828), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_775), .C(n_791), .Y(n_759) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_764), .A2(n_1141), .B1(n_1142), .B2(n_1143), .Y(n_1140) );
NAND3xp33_ASAP7_75t_L g1395 ( .A(n_765), .B(n_1396), .C(n_1399), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_768), .A2(n_782), .B1(n_784), .B2(n_785), .Y(n_781) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_SL g895 ( .A(n_773), .Y(n_895) );
OAI31xp33_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_779), .A3(n_786), .B(n_790), .Y(n_775) );
OAI22xp33_ASAP7_75t_L g823 ( .A1(n_780), .A2(n_797), .B1(n_805), .B2(n_824), .Y(n_823) );
BUFx3_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
BUFx3_ASAP7_75t_L g862 ( .A(n_783), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_785), .A2(n_862), .B1(n_863), .B2(n_864), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_785), .A2(n_862), .B1(n_882), .B2(n_883), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_785), .A2(n_862), .B1(n_1355), .B2(n_1365), .Y(n_1364) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
BUFx2_ASAP7_75t_L g887 ( .A(n_790), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g1672 ( .A1(n_790), .A2(n_1673), .B(n_1681), .Y(n_1672) );
NOR2xp33_ASAP7_75t_SL g791 ( .A(n_792), .B(n_813), .Y(n_791) );
OAI33xp33_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .A3(n_799), .B1(n_802), .B2(n_806), .B3(n_807), .Y(n_792) );
INVx2_ASAP7_75t_SL g1098 ( .A(n_793), .Y(n_1098) );
INVx2_ASAP7_75t_SL g1379 ( .A(n_793), .Y(n_1379) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_796), .B1(n_797), .B2(n_798), .Y(n_794) );
OAI22xp33_ASAP7_75t_L g815 ( .A1(n_795), .A2(n_804), .B1(n_816), .B2(n_817), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_796), .A2(n_798), .B1(n_839), .B2(n_843), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_796), .A2(n_1149), .B1(n_1150), .B2(n_1151), .Y(n_1148) );
OAI22xp33_ASAP7_75t_L g1328 ( .A1(n_796), .A2(n_798), .B1(n_1329), .B2(n_1330), .Y(n_1328) );
OAI22xp5_ASAP7_75t_L g1340 ( .A1(n_796), .A2(n_810), .B1(n_1341), .B2(n_1342), .Y(n_1340) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_798), .A2(n_902), .B1(n_914), .B2(n_919), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_798), .A2(n_907), .B1(n_912), .B2(n_919), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_800), .A2(n_809), .B1(n_819), .B2(n_821), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_809), .B1(n_810), .B2(n_812), .Y(n_807) );
BUFx3_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI33xp33_ASAP7_75t_L g1152 ( .A1(n_814), .A2(n_1153), .A3(n_1156), .B1(n_1158), .B2(n_1160), .B3(n_1161), .Y(n_1152) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_816), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g844 ( .A1(n_816), .A2(n_845), .B1(n_846), .B2(n_847), .Y(n_844) );
OAI22xp33_ASAP7_75t_L g901 ( .A1(n_816), .A2(n_902), .B1(n_903), .B2(n_904), .Y(n_901) );
OAI22xp33_ASAP7_75t_L g1344 ( .A1(n_816), .A2(n_1329), .B1(n_1337), .B2(n_1345), .Y(n_1344) );
OAI22xp33_ASAP7_75t_L g1350 ( .A1(n_816), .A2(n_1330), .B1(n_1339), .B2(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g1347 ( .A(n_820), .Y(n_1347) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_821), .A2(n_909), .B1(n_911), .B2(n_912), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_821), .A2(n_1141), .B1(n_1149), .B2(n_1157), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_821), .A2(n_1332), .B1(n_1341), .B2(n_1347), .Y(n_1346) );
OAI22xp5_ASAP7_75t_L g1348 ( .A1(n_821), .A2(n_1333), .B1(n_1342), .B2(n_1349), .Y(n_1348) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g1155 ( .A(n_826), .Y(n_1155) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
NAND3xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_854), .C(n_866), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_831), .B(n_848), .Y(n_830) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVxp67_ASAP7_75t_SL g1351 ( .A(n_860), .Y(n_1351) );
INVx1_ASAP7_75t_L g1273 ( .A(n_873), .Y(n_1273) );
XNOR2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_993), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_876), .B1(n_929), .B2(n_930), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g877 ( .A(n_878), .B(n_888), .C(n_898), .Y(n_877) );
OAI31xp33_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_880), .A3(n_884), .B(n_887), .Y(n_878) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
OAI31xp33_ASAP7_75t_L g1359 ( .A1(n_887), .A2(n_1360), .A3(n_1361), .B(n_1366), .Y(n_1359) );
OAI31xp33_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_893), .A3(n_896), .B(n_897), .Y(n_888) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
OAI31xp33_ASAP7_75t_L g1352 ( .A1(n_897), .A2(n_1353), .A3(n_1357), .B(n_1358), .Y(n_1352) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_916), .Y(n_898) );
OAI33xp33_ASAP7_75t_L g1080 ( .A1(n_900), .A2(n_1081), .A3(n_1084), .B1(n_1087), .B2(n_1091), .B3(n_1092), .Y(n_1080) );
OAI33xp33_ASAP7_75t_L g1283 ( .A1(n_900), .A2(n_1091), .A3(n_1284), .B1(n_1288), .B2(n_1292), .B3(n_1296), .Y(n_1283) );
OAI33xp33_ASAP7_75t_L g1386 ( .A1(n_900), .A2(n_1091), .A3(n_1387), .B1(n_1388), .B2(n_1389), .B3(n_1392), .Y(n_1386) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_903), .A2(n_915), .B1(n_923), .B2(n_927), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_906), .A2(n_911), .B1(n_923), .B2(n_925), .Y(n_922) );
INVx2_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx2_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_923), .A2(n_1083), .B1(n_1094), .B2(n_1102), .Y(n_1103) );
INVx4_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
NAND4xp25_ASAP7_75t_SL g932 ( .A(n_933), .B(n_943), .C(n_970), .D(n_988), .Y(n_932) );
AOI33xp33_ASAP7_75t_L g943 ( .A1(n_944), .A2(n_947), .A3(n_956), .B1(n_963), .B2(n_966), .B3(n_969), .Y(n_943) );
BUFx3_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g1188 ( .A(n_945), .Y(n_1188) );
INVx1_ASAP7_75t_L g1706 ( .A(n_946), .Y(n_1706) );
BUFx2_ASAP7_75t_SL g948 ( .A(n_949), .Y(n_948) );
INVx2_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
OAI221xp5_ASAP7_75t_L g1190 ( .A1(n_950), .A2(n_1191), .B1(n_1192), .B2(n_1193), .C(n_1194), .Y(n_1190) );
INVx2_ASAP7_75t_SL g950 ( .A(n_951), .Y(n_950) );
BUFx3_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx8_ASAP7_75t_L g1186 ( .A(n_952), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_954), .B(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx2_ASAP7_75t_L g1740 ( .A(n_955), .Y(n_1740) );
INVx2_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
BUFx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g967 ( .A(n_959), .Y(n_967) );
INVx3_ASAP7_75t_L g1011 ( .A(n_959), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1290 ( .A(n_959), .Y(n_1290) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx2_ASAP7_75t_L g968 ( .A(n_961), .Y(n_968) );
INVx5_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
BUFx2_ASAP7_75t_L g1688 ( .A(n_962), .Y(n_1688) );
BUFx12f_ASAP7_75t_L g1748 ( .A(n_962), .Y(n_1748) );
BUFx2_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
XOR2xp5_ASAP7_75t_L g993 ( .A(n_994), .B(n_1074), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
XNOR2x1_ASAP7_75t_L g996 ( .A(n_997), .B(n_1038), .Y(n_996) );
XNOR2xp5_ASAP7_75t_L g997 ( .A(n_998), .B(n_999), .Y(n_997) );
AND3x1_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1024), .C(n_1032), .Y(n_999) );
NOR2xp33_ASAP7_75t_SL g1000 ( .A(n_1001), .B(n_1016), .Y(n_1000) );
INVx2_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1011), .Y(n_1157) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_1019), .A2(n_1050), .B1(n_1051), .B2(n_1052), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1258 ( .A1(n_1019), .A2(n_1051), .B1(n_1259), .B2(n_1260), .Y(n_1258) );
OAI22xp5_ASAP7_75t_SL g1101 ( .A1(n_1021), .A2(n_1085), .B1(n_1089), .B2(n_1102), .Y(n_1101) );
OAI33xp33_ASAP7_75t_L g1096 ( .A1(n_1023), .A2(n_1097), .A3(n_1099), .B1(n_1101), .B2(n_1103), .B3(n_1104), .Y(n_1096) );
OAI33xp33_ASAP7_75t_L g1371 ( .A1(n_1023), .A2(n_1372), .A3(n_1375), .B1(n_1378), .B2(n_1380), .B3(n_1383), .Y(n_1371) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1027), .Y(n_1649) );
AND3x1_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1061), .C(n_1068), .Y(n_1039) );
NOR2xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1056), .Y(n_1040) );
OAI22xp33_ASAP7_75t_L g1136 ( .A1(n_1044), .A2(n_1137), .B1(n_1138), .B2(n_1139), .Y(n_1136) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_1051), .A2(n_1145), .B1(n_1287), .B2(n_1298), .Y(n_1302) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_1075), .A2(n_1076), .B1(n_1180), .B2(n_1272), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
AOI22xp5_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1131), .B1(n_1132), .B2(n_1179), .Y(n_1076) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1077), .Y(n_1179) );
INVxp67_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
NOR4xp25_ASAP7_75t_L g1130 ( .A(n_1080), .B(n_1096), .C(n_1106), .D(n_1121), .Y(n_1130) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1091), .Y(n_1194) );
INVxp67_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVxp67_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVxp67_ASAP7_75t_SL g1108 ( .A(n_1109), .Y(n_1108) );
AOI31xp67_ASAP7_75t_SL g1121 ( .A1(n_1122), .A2(n_1125), .A3(n_1127), .B(n_1129), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVxp67_ASAP7_75t_SL g1127 ( .A(n_1128), .Y(n_1127) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
NAND3xp33_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1163), .C(n_1171), .Y(n_1133) );
NOR2xp33_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1152), .Y(n_1134) );
OAI22xp33_ASAP7_75t_L g1161 ( .A1(n_1139), .A2(n_1147), .B1(n_1154), .B2(n_1162), .Y(n_1161) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1180), .Y(n_1272) );
XNOR2x1_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1236), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1218), .Y(n_1181) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1183), .Y(n_1220) );
AOI21xp5_ASAP7_75t_L g1183 ( .A1(n_1184), .A2(n_1187), .B(n_1189), .Y(n_1183) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
CKINVDCx5p33_ASAP7_75t_R g1739 ( .A(n_1186), .Y(n_1739) );
INVx8_ASAP7_75t_L g1752 ( .A(n_1186), .Y(n_1752) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1195), .B(n_1205), .Y(n_1219) );
OAI31xp33_ASAP7_75t_SL g1195 ( .A1(n_1196), .A2(n_1197), .A3(n_1203), .B(n_1204), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1202), .B(n_1215), .Y(n_1214) );
OAI31xp33_ASAP7_75t_SL g1245 ( .A1(n_1204), .A2(n_1246), .A3(n_1247), .B(n_1252), .Y(n_1245) );
OAI31xp33_ASAP7_75t_L g1403 ( .A1(n_1204), .A2(n_1404), .A3(n_1406), .B(n_1409), .Y(n_1403) );
NOR2xp33_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1212), .Y(n_1210) );
NAND3xp33_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1214), .C(n_1217), .Y(n_1212) );
INVx2_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
OAI31xp33_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1220), .A3(n_1221), .B(n_1233), .Y(n_1218) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1222), .Y(n_1235) );
BUFx6f_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1235), .Y(n_1233) );
NAND3xp33_ASAP7_75t_SL g1237 ( .A(n_1238), .B(n_1245), .C(n_1253), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1243), .B(n_1249), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1408 ( .A(n_1249), .B(n_1398), .Y(n_1408) );
NOR2xp33_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1267), .Y(n_1253) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
OAI22xp5_ASAP7_75t_L g1276 ( .A1(n_1277), .A2(n_1278), .B1(n_1367), .B2(n_1368), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
XNOR2xp5_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1323), .Y(n_1278) );
HB1xp67_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
NAND3xp33_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1305), .C(n_1313), .Y(n_1281) );
NOR2xp33_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1299), .Y(n_1282) );
OAI22xp5_ASAP7_75t_L g1389 ( .A1(n_1293), .A2(n_1374), .B1(n_1382), .B2(n_1390), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1316), .B(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
NAND3xp33_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1352), .C(n_1359), .Y(n_1325) );
NOR2xp33_ASAP7_75t_SL g1326 ( .A(n_1327), .B(n_1343), .Y(n_1326) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_1335), .A2(n_1337), .B1(n_1338), .B2(n_1339), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
INVxp67_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx3_ASAP7_75t_SL g1367 ( .A(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1369), .Y(n_1411) );
NAND3xp33_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1393), .C(n_1403), .Y(n_1369) );
NOR2xp33_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1386), .Y(n_1370) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
OAI221xp5_ASAP7_75t_SL g1413 ( .A1(n_1414), .A2(n_1639), .B1(n_1641), .B2(n_1691), .C(n_1695), .Y(n_1413) );
NOR5xp2_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1554), .C(n_1616), .D(n_1622), .E(n_1633), .Y(n_1414) );
AOI31xp33_ASAP7_75t_L g1415 ( .A1(n_1416), .A2(n_1498), .A3(n_1528), .B(n_1548), .Y(n_1415) );
AOI211xp5_ASAP7_75t_SL g1416 ( .A1(n_1417), .A2(n_1433), .B(n_1452), .C(n_1466), .Y(n_1416) );
A2O1A1Ixp33_ASAP7_75t_L g1555 ( .A1(n_1417), .A2(n_1556), .B(n_1558), .C(n_1570), .Y(n_1555) );
CKINVDCx6p67_ASAP7_75t_R g1417 ( .A(n_1418), .Y(n_1417) );
CKINVDCx6p67_ASAP7_75t_R g1418 ( .A(n_1419), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1419), .B(n_1494), .Y(n_1496) );
INVx2_ASAP7_75t_L g1506 ( .A(n_1419), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1419), .B(n_1566), .Y(n_1565) );
OAI22xp5_ASAP7_75t_L g1576 ( .A1(n_1419), .A2(n_1577), .B1(n_1579), .B2(n_1581), .Y(n_1576) );
AND2x4_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1427), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1420), .B(n_1427), .Y(n_1458) );
AND2x6_ASAP7_75t_L g1421 ( .A(n_1422), .B(n_1423), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1422), .B(n_1426), .Y(n_1425) );
AND2x4_ASAP7_75t_L g1428 ( .A(n_1422), .B(n_1429), .Y(n_1428) );
AND2x6_ASAP7_75t_L g1431 ( .A(n_1422), .B(n_1432), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1422), .B(n_1426), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1422), .B(n_1426), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1424), .B(n_1430), .Y(n_1429) );
OAI21xp5_ASAP7_75t_L g1760 ( .A1(n_1426), .A2(n_1761), .B(n_1762), .Y(n_1760) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1435), .B(n_1440), .Y(n_1434) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1435), .B(n_1481), .Y(n_1480) );
NAND2xp5_ASAP7_75t_SL g1502 ( .A(n_1435), .B(n_1503), .Y(n_1502) );
OR2x2_ASAP7_75t_L g1581 ( .A(n_1435), .B(n_1582), .Y(n_1581) );
INVx2_ASAP7_75t_L g1585 ( .A(n_1435), .Y(n_1585) );
INVx2_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx3_ASAP7_75t_L g1460 ( .A(n_1436), .Y(n_1460) );
NOR2xp33_ASAP7_75t_L g1478 ( .A(n_1436), .B(n_1441), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1436), .B(n_1511), .Y(n_1510) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1436), .B(n_1441), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_1436), .B(n_1475), .Y(n_1537) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1436), .B(n_1524), .Y(n_1567) );
NOR2xp33_ASAP7_75t_L g1575 ( .A(n_1436), .B(n_1486), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1438), .Y(n_1436) );
HB1xp67_ASAP7_75t_L g1640 ( .A(n_1439), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1620 ( .A(n_1440), .B(n_1470), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1445), .Y(n_1440) );
CKINVDCx5p33_ASAP7_75t_R g1501 ( .A(n_1441), .Y(n_1501) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_1441), .B(n_1513), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1441), .B(n_1464), .Y(n_1590) );
OR2x2_ASAP7_75t_L g1602 ( .A(n_1441), .B(n_1477), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1605 ( .A(n_1441), .B(n_1538), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1444), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1442), .B(n_1444), .Y(n_1462) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1445), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1445), .B(n_1533), .Y(n_1543) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1445), .B(n_1501), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1449), .Y(n_1445) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1446), .Y(n_1465) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1446), .Y(n_1538) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1448), .Y(n_1446) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1449), .Y(n_1464) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1449), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1449), .B(n_1465), .Y(n_1490) );
OR2x2_ASAP7_75t_L g1504 ( .A(n_1449), .B(n_1465), .Y(n_1504) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1451), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1453), .B(n_1459), .Y(n_1452) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
OR2x2_ASAP7_75t_L g1454 ( .A(n_1455), .B(n_1458), .Y(n_1454) );
INVx3_ASAP7_75t_L g1475 ( .A(n_1455), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1455), .B(n_1492), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1455), .B(n_1506), .Y(n_1505) );
OR2x2_ASAP7_75t_L g1508 ( .A(n_1455), .B(n_1493), .Y(n_1508) );
NOR2xp33_ASAP7_75t_L g1516 ( .A(n_1455), .B(n_1469), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1455), .B(n_1458), .Y(n_1530) );
AND2x2_ASAP7_75t_L g1544 ( .A(n_1455), .B(n_1469), .Y(n_1544) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1455), .B(n_1520), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1455), .B(n_1524), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1455), .B(n_1570), .Y(n_1588) );
INVx3_ASAP7_75t_L g1632 ( .A(n_1455), .Y(n_1632) );
AND2x4_ASAP7_75t_SL g1455 ( .A(n_1456), .B(n_1457), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1458), .B(n_1475), .Y(n_1474) );
OR2x2_ASAP7_75t_L g1482 ( .A(n_1458), .B(n_1471), .Y(n_1482) );
OR2x2_ASAP7_75t_L g1493 ( .A(n_1458), .B(n_1494), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1458), .B(n_1471), .Y(n_1520) );
NOR2xp33_ASAP7_75t_L g1603 ( .A(n_1458), .B(n_1551), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1461), .Y(n_1459) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1460), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1557 ( .A(n_1460), .B(n_1490), .Y(n_1557) );
NOR2xp33_ASAP7_75t_L g1560 ( .A(n_1460), .B(n_1504), .Y(n_1560) );
O2A1O1Ixp33_ASAP7_75t_L g1562 ( .A1(n_1460), .A2(n_1520), .B(n_1563), .C(n_1564), .Y(n_1562) );
NAND2xp5_ASAP7_75t_L g1592 ( .A(n_1460), .B(n_1494), .Y(n_1592) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1460), .B(n_1596), .Y(n_1595) );
NOR2xp33_ASAP7_75t_L g1601 ( .A(n_1460), .B(n_1602), .Y(n_1601) );
NOR2xp33_ASAP7_75t_L g1604 ( .A(n_1460), .B(n_1605), .Y(n_1604) );
NAND3xp33_ASAP7_75t_L g1608 ( .A(n_1460), .B(n_1570), .C(n_1609), .Y(n_1608) );
NAND2xp5_ASAP7_75t_L g1625 ( .A(n_1460), .B(n_1492), .Y(n_1625) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1461), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1462), .B(n_1463), .Y(n_1461) );
AOI32xp33_ASAP7_75t_L g1479 ( .A1(n_1462), .A2(n_1480), .A3(n_1483), .B1(n_1487), .B2(n_1491), .Y(n_1479) );
OR2x2_ASAP7_75t_L g1488 ( .A(n_1462), .B(n_1489), .Y(n_1488) );
OR2x2_ASAP7_75t_L g1526 ( .A(n_1462), .B(n_1527), .Y(n_1526) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1462), .B(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1463), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_1463), .B(n_1501), .Y(n_1540) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1463), .B(n_1478), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1546 ( .A(n_1463), .B(n_1547), .Y(n_1546) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1465), .Y(n_1463) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1465), .Y(n_1513) );
OAI211xp5_ASAP7_75t_L g1466 ( .A1(n_1467), .A2(n_1476), .B(n_1479), .C(n_1495), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1474), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1578 ( .A(n_1469), .B(n_1532), .Y(n_1578) );
O2A1O1Ixp33_ASAP7_75t_L g1626 ( .A1(n_1469), .A2(n_1557), .B(n_1563), .C(n_1627), .Y(n_1626) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1469), .Y(n_1629) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1470), .B(n_1532), .Y(n_1531) );
AOI322xp5_ASAP7_75t_L g1600 ( .A1(n_1470), .A2(n_1516), .A3(n_1542), .B1(n_1588), .B2(n_1601), .C1(n_1603), .C2(n_1604), .Y(n_1600) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1471), .Y(n_1494) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1471), .Y(n_1524) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1473), .Y(n_1471) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1474), .Y(n_1621) );
NAND2xp5_ASAP7_75t_L g1599 ( .A(n_1475), .B(n_1481), .Y(n_1599) );
OR2x2_ASAP7_75t_L g1611 ( .A(n_1475), .B(n_1482), .Y(n_1611) );
AOI32xp33_ASAP7_75t_L g1635 ( .A1(n_1475), .A2(n_1480), .A3(n_1569), .B1(n_1570), .B2(n_1636), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1478), .Y(n_1476) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1477), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1478), .B(n_1490), .Y(n_1497) );
AOI311xp33_ASAP7_75t_L g1583 ( .A1(n_1481), .A2(n_1584), .A3(n_1585), .B(n_1586), .C(n_1597), .Y(n_1583) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
OAI321xp33_ASAP7_75t_L g1534 ( .A1(n_1482), .A2(n_1535), .A3(n_1536), .B1(n_1538), .B2(n_1539), .C(n_1541), .Y(n_1534) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
NAND2xp5_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1486), .Y(n_1484) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
OR2x2_ASAP7_75t_L g1638 ( .A(n_1489), .B(n_1501), .Y(n_1638) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
NAND2xp5_ASAP7_75t_L g1527 ( .A(n_1490), .B(n_1519), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1490), .B(n_1533), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1492), .B(n_1519), .Y(n_1615) );
INVx2_ASAP7_75t_SL g1492 ( .A(n_1493), .Y(n_1492) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1497), .Y(n_1495) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1496), .Y(n_1535) );
AOI221xp5_ASAP7_75t_L g1498 ( .A1(n_1499), .A2(n_1505), .B1(n_1507), .B2(n_1509), .C(n_1514), .Y(n_1498) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
OR2x2_ASAP7_75t_L g1500 ( .A(n_1501), .B(n_1502), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1501), .B(n_1538), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_1501), .B(n_1560), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1501), .B(n_1513), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1598 ( .A(n_1503), .B(n_1533), .Y(n_1598) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1505), .Y(n_1561) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
INVxp67_ASAP7_75t_SL g1509 ( .A(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
A2O1A1Ixp33_ASAP7_75t_L g1514 ( .A1(n_1515), .A2(n_1517), .B(n_1521), .C(n_1522), .Y(n_1514) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1519), .B(n_1520), .Y(n_1518) );
CKINVDCx14_ASAP7_75t_R g1634 ( .A(n_1520), .Y(n_1634) );
NAND2xp5_ASAP7_75t_L g1584 ( .A(n_1521), .B(n_1582), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_1523), .B(n_1525), .Y(n_1522) );
NAND2xp5_ASAP7_75t_L g1617 ( .A(n_1523), .B(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_1526), .B(n_1574), .Y(n_1573) );
AOI211xp5_ASAP7_75t_L g1528 ( .A1(n_1529), .A2(n_1531), .B(n_1534), .C(n_1545), .Y(n_1528) );
NAND3xp33_ASAP7_75t_L g1593 ( .A(n_1529), .B(n_1550), .C(n_1594), .Y(n_1593) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
A2O1A1Ixp33_ASAP7_75t_L g1586 ( .A1(n_1530), .A2(n_1587), .B(n_1589), .C(n_1593), .Y(n_1586) );
NOR2xp33_ASAP7_75t_L g1564 ( .A(n_1535), .B(n_1539), .Y(n_1564) );
OAI221xp5_ASAP7_75t_SL g1597 ( .A1(n_1535), .A2(n_1539), .B1(n_1598), .B2(n_1599), .C(n_1600), .Y(n_1597) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1538), .Y(n_1609) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
OAI21xp5_ASAP7_75t_L g1541 ( .A1(n_1542), .A2(n_1543), .B(n_1544), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1628 ( .A(n_1543), .B(n_1629), .Y(n_1628) );
AOI221xp5_ASAP7_75t_L g1571 ( .A1(n_1544), .A2(n_1547), .B1(n_1572), .B2(n_1573), .C(n_1576), .Y(n_1571) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1544), .Y(n_1637) );
INVxp67_ASAP7_75t_SL g1545 ( .A(n_1546), .Y(n_1545) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1550), .B(n_1632), .Y(n_1631) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1551), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1553), .Y(n_1551) );
NAND4xp25_ASAP7_75t_L g1554 ( .A(n_1555), .B(n_1571), .C(n_1583), .D(n_1606), .Y(n_1554) );
CKINVDCx14_ASAP7_75t_R g1619 ( .A(n_1556), .Y(n_1619) );
OAI211xp5_ASAP7_75t_SL g1558 ( .A1(n_1559), .A2(n_1561), .B(n_1562), .C(n_1565), .Y(n_1558) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1563), .Y(n_1582) );
O2A1O1Ixp33_ASAP7_75t_L g1606 ( .A1(n_1563), .A2(n_1607), .B(n_1610), .C(n_1612), .Y(n_1606) );
NOR2xp33_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1568), .Y(n_1566) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1581), .Y(n_1618) );
O2A1O1Ixp33_ASAP7_75t_L g1612 ( .A1(n_1587), .A2(n_1598), .B(n_1613), .C(n_1614), .Y(n_1612) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1589 ( .A(n_1590), .B(n_1591), .Y(n_1589) );
O2A1O1Ixp33_ASAP7_75t_L g1622 ( .A1(n_1590), .A2(n_1623), .B(n_1626), .C(n_1630), .Y(n_1622) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVxp67_ASAP7_75t_SL g1607 ( .A(n_1608), .Y(n_1607) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
A2O1A1Ixp33_ASAP7_75t_L g1633 ( .A1(n_1611), .A2(n_1619), .B(n_1634), .C(n_1635), .Y(n_1633) );
INVxp67_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
AOI31xp33_ASAP7_75t_L g1616 ( .A1(n_1617), .A2(n_1619), .A3(n_1620), .B(n_1621), .Y(n_1616) );
INVxp67_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1628), .Y(n_1627) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
NOR2xp33_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1638), .Y(n_1636) );
INVx4_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
HB1xp67_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
OAI21xp5_ASAP7_75t_L g1643 ( .A1(n_1644), .A2(n_1670), .B(n_1672), .Y(n_1643) );
OAI21xp5_ASAP7_75t_L g1656 ( .A1(n_1657), .A2(n_1660), .B(n_1663), .Y(n_1656) );
INVx2_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1667), .Y(n_1721) );
BUFx2_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
NAND2xp5_ASAP7_75t_SL g1673 ( .A(n_1674), .B(n_1679), .Y(n_1673) );
OAI211xp5_ASAP7_75t_L g1682 ( .A1(n_1683), .A2(n_1684), .B(n_1686), .C(n_1687), .Y(n_1682) );
INVx2_ASAP7_75t_SL g1684 ( .A(n_1685), .Y(n_1684) );
CKINVDCx5p33_ASAP7_75t_R g1691 ( .A(n_1692), .Y(n_1691) );
BUFx2_ASAP7_75t_SL g1692 ( .A(n_1693), .Y(n_1692) );
BUFx3_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
BUFx3_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
HB1xp67_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
HB1xp67_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
XNOR2x1_ASAP7_75t_L g1701 ( .A(n_1702), .B(n_1703), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1745), .Y(n_1703) );
AOI21xp5_ASAP7_75t_L g1704 ( .A1(n_1705), .A2(n_1707), .B(n_1734), .Y(n_1704) );
HB1xp67_ASAP7_75t_L g1705 ( .A(n_1706), .Y(n_1705) );
NAND4xp25_ASAP7_75t_L g1707 ( .A(n_1708), .B(n_1713), .C(n_1718), .D(n_1723), .Y(n_1707) );
OAI21xp5_ASAP7_75t_L g1708 ( .A1(n_1709), .A2(n_1710), .B(n_1711), .Y(n_1708) );
BUFx2_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
HB1xp67_ASAP7_75t_L g1732 ( .A(n_1733), .Y(n_1732) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
endmodule