module fake_jpeg_5242_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_18),
.B(n_16),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_6),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_20),
.B(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_49),
.Y(n_58)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_28),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_7),
.B(n_13),
.Y(n_53)
);

HAxp5_ASAP7_75t_SL g95 ( 
.A(n_53),
.B(n_18),
.CON(n_95),
.SN(n_95)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_66),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_60),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_31),
.B1(n_20),
.B2(n_33),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_83),
.B1(n_36),
.B2(n_29),
.Y(n_106)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_72),
.Y(n_100)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_71),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_31),
.B1(n_35),
.B2(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_73),
.B1(n_36),
.B2(n_34),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_28),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_31),
.B1(n_35),
.B2(n_23),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_75),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_33),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_30),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_77),
.Y(n_121)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_32),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_32),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_19),
.B1(n_18),
.B2(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

BUFx16f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_19),
.B1(n_36),
.B2(n_29),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_95),
.B(n_34),
.C(n_27),
.Y(n_103)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_39),
.B(n_22),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_96),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_37),
.B(n_12),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_34),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_27),
.B1(n_22),
.B2(n_25),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_58),
.C(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_113),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_103),
.A2(n_120),
.B1(n_108),
.B2(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_73),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_69),
.B1(n_82),
.B2(n_59),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_34),
.C(n_27),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_63),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_94),
.B1(n_56),
.B2(n_24),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_25),
.B1(n_27),
.B2(n_17),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_126),
.B1(n_82),
.B2(n_69),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_55),
.A2(n_17),
.B1(n_24),
.B2(n_2),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_57),
.B(n_24),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_128),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_70),
.B(n_0),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_116),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_64),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_120),
.B(n_102),
.C(n_124),
.D(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_135),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_142),
.B1(n_147),
.B2(n_161),
.Y(n_163)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_136),
.B(n_139),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_64),
.C(n_88),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g179 ( 
.A(n_137),
.B(n_149),
.C(n_131),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_88),
.A3(n_55),
.B1(n_91),
.B2(n_68),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_141),
.Y(n_181)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_122),
.B1(n_123),
.B2(n_114),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_100),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_93),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_143),
.A2(n_157),
.B1(n_147),
.B2(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_145),
.C(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_103),
.B(n_74),
.C(n_66),
.Y(n_149)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_59),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_152),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_109),
.B(n_63),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_112),
.A2(n_75),
.B1(n_79),
.B2(n_98),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_62),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_108),
.B(n_11),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_166),
.B(n_1),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_121),
.B1(n_114),
.B2(n_122),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_168),
.B(n_184),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_136),
.B(n_130),
.C(n_139),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_172),
.B1(n_151),
.B2(n_148),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_123),
.B1(n_119),
.B2(n_111),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_121),
.B1(n_99),
.B2(n_111),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_173),
.A2(n_174),
.B(n_3),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_99),
.B(n_62),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_117),
.C(n_2),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_187),
.C(n_5),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_190),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_7),
.B1(n_15),
.B2(n_12),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_138),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_149),
.C(n_143),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_197),
.Y(n_225)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_194),
.B(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_191),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_145),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_208),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_192),
.A2(n_135),
.B1(n_132),
.B2(n_142),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_206),
.Y(n_224)
);

A2O1A1O1Ixp25_ASAP7_75t_L g201 ( 
.A1(n_181),
.A2(n_155),
.B(n_7),
.C(n_8),
.D(n_4),
.Y(n_201)
);

AOI221xp5_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_204),
.B1(n_213),
.B2(n_3),
.C(n_185),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_186),
.B(n_175),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_182),
.B(n_5),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_189),
.C(n_180),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_162),
.B(n_15),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_189),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_177),
.A2(n_2),
.B1(n_3),
.B2(n_15),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_212),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_169),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_173),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_220),
.C(n_234),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_226),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_170),
.C(n_163),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_205),
.A2(n_167),
.B(n_176),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_233),
.B(n_200),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_190),
.B1(n_167),
.B2(n_166),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_222),
.A2(n_197),
.B1(n_193),
.B2(n_203),
.Y(n_242)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_201),
.B(n_176),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_229),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_185),
.C(n_165),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

OA21x2_ASAP7_75t_SL g243 ( 
.A1(n_236),
.A2(n_207),
.B(n_208),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_194),
.B(n_204),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_225),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_213),
.C(n_199),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_217),
.C(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_224),
.A2(n_196),
.B1(n_203),
.B2(n_202),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_247),
.B1(n_196),
.B2(n_226),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_221),
.B1(n_218),
.B2(n_222),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_252),
.C(n_254),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_234),
.C(n_219),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_223),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_230),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_238),
.C(n_240),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_248),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_257),
.A2(n_246),
.B(n_249),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_245),
.B1(n_247),
.B2(n_246),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_253),
.B(n_250),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_260),
.A2(n_237),
.B(n_243),
.C(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_265),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_262),
.B(n_195),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_240),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_269),
.A2(n_263),
.B(n_244),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_271),
.B(n_241),
.Y(n_272)
);

AOI21x1_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_255),
.B(n_242),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_267),
.Y(n_273)
);


endmodule