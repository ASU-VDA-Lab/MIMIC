module fake_netlist_6_399_n_794 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_794);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_794;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_772;
wire n_656;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g151 ( 
.A(n_16),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_59),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_22),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_26),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_32),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_8),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_93),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_36),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_13),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_12),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_9),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_141),
.Y(n_172)
);

BUFx2_ASAP7_75t_SL g173 ( 
.A(n_21),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_97),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_123),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_77),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_51),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_134),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_19),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_18),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_128),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_35),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_81),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_42),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_21),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_10),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_4),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_39),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_48),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_80),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_110),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_124),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_10),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_129),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_61),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_22),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_43),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_92),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_12),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_72),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_54),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_14),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_58),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_0),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_0),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_1),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_1),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_153),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_198),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_157),
.B(n_2),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_165),
.Y(n_235)
);

BUFx8_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_157),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_155),
.B(n_2),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_158),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_158),
.B(n_3),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_176),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_3),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_178),
.B(n_4),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_173),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_205),
.B1(n_195),
.B2(n_167),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g251 ( 
.A(n_209),
.B(n_179),
.Y(n_251)
);

OA22x2_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_166),
.B1(n_180),
.B2(n_189),
.Y(n_252)
);

NAND3x1_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_5),
.C(n_6),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_179),
.B1(n_204),
.B2(n_200),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_182),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_217),
.B(n_197),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

OR2x6_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_197),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_200),
.B1(n_204),
.B2(n_206),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

AO22x2_ASAP7_75t_L g261 ( 
.A1(n_209),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_239),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_229),
.A2(n_196),
.B1(n_194),
.B2(n_193),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_183),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_192),
.Y(n_266)
);

AO22x2_ASAP7_75t_L g267 ( 
.A1(n_238),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_229),
.A2(n_191),
.B1(n_190),
.B2(n_186),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_225),
.B(n_185),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

AO22x2_ASAP7_75t_L g272 ( 
.A1(n_238),
.A2(n_246),
.B1(n_234),
.B2(n_249),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_27),
.Y(n_273)
);

AO22x2_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_249),
.B1(n_248),
.B2(n_233),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_233),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_225),
.B(n_230),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_217),
.A2(n_11),
.B1(n_15),
.B2(n_16),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_225),
.B(n_15),
.Y(n_278)
);

AO22x2_ASAP7_75t_L g279 ( 
.A1(n_207),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_230),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_211),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_211),
.Y(n_282)
);

AND2x4_ASAP7_75t_L g283 ( 
.A(n_217),
.B(n_227),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_230),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_207),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

AO22x2_ASAP7_75t_L g287 ( 
.A1(n_210),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_230),
.B(n_30),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_208),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_217),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_210),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g292 ( 
.A1(n_217),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_237),
.B(n_41),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_237),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_237),
.B(n_47),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_211),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_211),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_235),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_297),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_237),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_217),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_263),
.B(n_241),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_289),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_257),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

INVx4_ASAP7_75t_SL g307 ( 
.A(n_283),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

BUFx8_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

INVx4_ASAP7_75t_SL g312 ( 
.A(n_283),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_263),
.B(n_241),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_217),
.Y(n_314)
);

XNOR2x2_ASAP7_75t_L g315 ( 
.A(n_261),
.B(n_267),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_298),
.A2(n_226),
.B(n_215),
.Y(n_316)
);

AND2x2_ASAP7_75t_SL g317 ( 
.A(n_251),
.B(n_241),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_276),
.B(n_235),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_262),
.B(n_236),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_286),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_255),
.B(n_235),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_297),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_297),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_266),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_271),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_268),
.B(n_241),
.Y(n_331)
);

INVxp33_ASAP7_75t_SL g332 ( 
.A(n_264),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_290),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_252),
.B(n_236),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_288),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_268),
.B(n_235),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_271),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_294),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_254),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_287),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_258),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_250),
.B(n_227),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_287),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_L g348 ( 
.A(n_250),
.B(n_228),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_253),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_256),
.B(n_245),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_292),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_261),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_267),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_279),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_279),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_258),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_280),
.B(n_236),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_280),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_284),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_284),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_291),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_258),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_285),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_245),
.Y(n_364)
);

NAND2x1p5_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_214),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_SL g366 ( 
.A(n_329),
.B(n_227),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_299),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_299),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_245),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_334),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_302),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_314),
.Y(n_373)
);

BUFx8_ASAP7_75t_L g374 ( 
.A(n_345),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_317),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_245),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_350),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_305),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_305),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_245),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_346),
.B(n_227),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g386 ( 
.A(n_336),
.B(n_214),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_317),
.B(n_227),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_308),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_326),
.B(n_227),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_304),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_348),
.B(n_227),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g394 ( 
.A(n_336),
.B(n_245),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_306),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_327),
.B(n_343),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_309),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_232),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_310),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_358),
.B(n_232),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_208),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_301),
.B(n_215),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_328),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_301),
.B(n_215),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_311),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

NAND2x1p5_ASAP7_75t_L g407 ( 
.A(n_340),
.B(n_214),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_318),
.B(n_228),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_351),
.B(n_212),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_352),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_324),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_316),
.B(n_228),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_303),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_328),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_303),
.B(n_228),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_322),
.A2(n_226),
.B(n_221),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_309),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_354),
.B(n_277),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_313),
.B(n_239),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_333),
.Y(n_420)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_307),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_313),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_362),
.B(n_212),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_353),
.B(n_221),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_331),
.B(n_228),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_331),
.B(n_228),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_359),
.B(n_221),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_344),
.B(n_347),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_355),
.Y(n_430)
);

BUFx4f_ASAP7_75t_L g431 ( 
.A(n_361),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_300),
.B(n_228),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_359),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_396),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_396),
.B(n_356),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_402),
.B(n_361),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_341),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_427),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_341),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_414),
.Y(n_444)
);

NAND2x1_ASAP7_75t_SL g445 ( 
.A(n_387),
.B(n_315),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_384),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_378),
.B(n_312),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_372),
.B(n_315),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_372),
.B(n_307),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_373),
.B(n_307),
.Y(n_451)
);

NAND2x1_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_307),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_388),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_367),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_431),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_402),
.B(n_404),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_369),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

NOR2x1_ASAP7_75t_L g459 ( 
.A(n_387),
.B(n_338),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_378),
.B(n_312),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_404),
.B(n_398),
.Y(n_462)
);

AND2x2_ASAP7_75t_SL g463 ( 
.A(n_376),
.B(n_291),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_380),
.B(n_285),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

NAND2x1_ASAP7_75t_L g466 ( 
.A(n_421),
.B(n_312),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_398),
.B(n_214),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_423),
.B(n_424),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_401),
.B(n_357),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_376),
.B(n_219),
.Y(n_471)
);

NOR2x1_ASAP7_75t_L g472 ( 
.A(n_419),
.B(n_421),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_401),
.B(n_320),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_369),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_423),
.B(n_49),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_400),
.B(n_431),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g478 ( 
.A(n_373),
.B(n_219),
.Y(n_478)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_374),
.Y(n_479)
);

BUFx4f_ASAP7_75t_L g480 ( 
.A(n_429),
.Y(n_480)
);

NAND2x1p5_ASAP7_75t_L g481 ( 
.A(n_373),
.B(n_219),
.Y(n_481)
);

NOR2x1_ASAP7_75t_SL g482 ( 
.A(n_373),
.B(n_375),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_410),
.B(n_236),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_390),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_381),
.Y(n_485)
);

AND2x2_ASAP7_75t_SL g486 ( 
.A(n_373),
.B(n_222),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_423),
.B(n_50),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_371),
.B(n_239),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_381),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_375),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_437),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_437),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_433),
.B(n_332),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_446),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_444),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_434),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_490),
.B(n_436),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_400),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_435),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_439),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_448),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_448),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_453),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_440),
.B(n_409),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_479),
.Y(n_507)
);

INVx3_ASAP7_75t_SL g508 ( 
.A(n_479),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_460),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_375),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

BUFx2_ASAP7_75t_R g512 ( 
.A(n_470),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_437),
.Y(n_513)
);

NAND2x1p5_ASAP7_75t_L g514 ( 
.A(n_450),
.B(n_375),
.Y(n_514)
);

CKINVDCx11_ASAP7_75t_R g515 ( 
.A(n_464),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_450),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_450),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_440),
.B(n_409),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_474),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_479),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_450),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_456),
.A2(n_407),
.B1(n_383),
.B2(n_375),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_457),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_470),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_448),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_436),
.B(n_429),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_480),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_486),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_480),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_443),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_478),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_473),
.Y(n_533)
);

BUFx4f_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_448),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_456),
.B(n_409),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_478),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_462),
.B(n_424),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_481),
.Y(n_539)
);

INVx6_ASAP7_75t_L g540 ( 
.A(n_530),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_496),
.B(n_433),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_502),
.B(n_469),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_500),
.B(n_462),
.Y(n_543)
);

CKINVDCx11_ASAP7_75t_R g544 ( 
.A(n_507),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_523),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_523),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_534),
.A2(n_463),
.B1(n_438),
.B2(n_476),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_516),
.Y(n_549)
);

BUFx12f_ASAP7_75t_L g550 ( 
.A(n_515),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_528),
.A2(n_438),
.B1(n_455),
.B2(n_458),
.Y(n_551)
);

CKINVDCx6p67_ASAP7_75t_R g552 ( 
.A(n_508),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_500),
.B(n_463),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_SL g554 ( 
.A1(n_534),
.A2(n_363),
.B1(n_275),
.B2(n_332),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_533),
.Y(n_555)
);

INVx8_ASAP7_75t_L g556 ( 
.A(n_521),
.Y(n_556)
);

CKINVDCx6p67_ASAP7_75t_R g557 ( 
.A(n_508),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_534),
.A2(n_484),
.B1(n_275),
.B2(n_471),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_528),
.A2(n_488),
.B1(n_407),
.B2(n_465),
.Y(n_559)
);

CKINVDCx14_ASAP7_75t_R g560 ( 
.A(n_533),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_521),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_494),
.A2(n_468),
.B1(n_488),
.B2(n_487),
.Y(n_562)
);

BUFx12f_ASAP7_75t_L g563 ( 
.A(n_520),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_493),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_493),
.Y(n_565)
);

OAI22xp33_ASAP7_75t_L g566 ( 
.A1(n_528),
.A2(n_363),
.B1(n_464),
.B2(n_465),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_495),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_503),
.A2(n_468),
.B1(n_475),
.B2(n_487),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_495),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_505),
.Y(n_570)
);

NAND2x1p5_ASAP7_75t_L g571 ( 
.A(n_521),
.B(n_449),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_531),
.A2(n_459),
.B(n_483),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_536),
.A2(n_471),
.B1(n_467),
.B2(n_441),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_503),
.A2(n_525),
.B1(n_535),
.B2(n_504),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_505),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_519),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_519),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_520),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_509),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_497),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_L g581 ( 
.A1(n_529),
.A2(n_464),
.B1(n_483),
.B2(n_454),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_509),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_553),
.B(n_498),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_581),
.A2(n_525),
.B1(n_504),
.B2(n_535),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_581),
.A2(n_529),
.B1(n_475),
.B2(n_518),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_542),
.B(n_498),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_558),
.A2(n_529),
.B1(n_506),
.B2(n_538),
.Y(n_587)
);

NAND3xp33_ASAP7_75t_L g588 ( 
.A(n_562),
.B(n_374),
.C(n_364),
.Y(n_588)
);

OAI21xp33_ASAP7_75t_L g589 ( 
.A1(n_558),
.A2(n_445),
.B(n_370),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_548),
.A2(n_529),
.B1(n_512),
.B2(n_407),
.Y(n_590)
);

NAND3xp33_ASAP7_75t_L g591 ( 
.A(n_572),
.B(n_374),
.C(n_377),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_559),
.A2(n_529),
.B1(n_417),
.B2(n_397),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_SL g593 ( 
.A1(n_560),
.A2(n_397),
.B1(n_380),
.B2(n_417),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_545),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_555),
.A2(n_548),
.B1(n_566),
.B2(n_568),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_546),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_547),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_566),
.A2(n_501),
.B1(n_527),
.B2(n_497),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_564),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_565),
.Y(n_600)
);

OAI22xp33_ASAP7_75t_L g601 ( 
.A1(n_541),
.A2(n_527),
.B1(n_530),
.B2(n_501),
.Y(n_601)
);

OAI222xp33_ASAP7_75t_L g602 ( 
.A1(n_554),
.A2(n_386),
.B1(n_467),
.B2(n_522),
.C1(n_418),
.C2(n_489),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_554),
.B(n_543),
.C(n_551),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_574),
.A2(n_530),
.B1(n_392),
.B2(n_391),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_573),
.B(n_510),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_574),
.A2(n_530),
.B1(n_392),
.B2(n_391),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_573),
.A2(n_530),
.B1(n_394),
.B2(n_524),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_567),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_556),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_580),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_569),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_578),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_570),
.A2(n_418),
.B(n_472),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_544),
.A2(n_526),
.B1(n_524),
.B2(n_510),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_575),
.A2(n_385),
.B(n_447),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_576),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_577),
.A2(n_521),
.B1(n_514),
.B2(n_430),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_582),
.A2(n_394),
.B1(n_420),
.B2(n_526),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_540),
.A2(n_394),
.B1(n_526),
.B2(n_399),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_540),
.A2(n_394),
.B1(n_526),
.B2(n_379),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_579),
.B(n_510),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_550),
.A2(n_482),
.B1(n_394),
.B2(n_385),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_549),
.Y(n_623)
);

OAI21xp33_ASAP7_75t_L g624 ( 
.A1(n_571),
.A2(n_424),
.B(n_405),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_552),
.B(n_510),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_540),
.A2(n_394),
.B1(n_379),
.B2(n_405),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_549),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_557),
.A2(n_379),
.B1(n_428),
.B2(n_395),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_563),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_549),
.Y(n_630)
);

OAI21xp33_ASAP7_75t_L g631 ( 
.A1(n_571),
.A2(n_389),
.B(n_426),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_549),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_556),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_SL g634 ( 
.A1(n_556),
.A2(n_539),
.B1(n_537),
.B2(n_532),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_589),
.A2(n_485),
.B1(n_226),
.B2(n_222),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_SL g636 ( 
.A1(n_588),
.A2(n_415),
.B1(n_425),
.B2(n_537),
.Y(n_636)
);

AOI222xp33_ASAP7_75t_L g637 ( 
.A1(n_603),
.A2(n_389),
.B1(n_222),
.B2(n_406),
.C1(n_428),
.C2(n_219),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_591),
.A2(n_395),
.B1(n_379),
.B2(n_537),
.Y(n_638)
);

AOI222xp33_ASAP7_75t_L g639 ( 
.A1(n_590),
.A2(n_602),
.B1(n_587),
.B2(n_583),
.C1(n_585),
.C2(n_586),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_590),
.A2(n_379),
.B1(n_539),
.B2(n_532),
.Y(n_640)
);

OAI221xp5_ASAP7_75t_L g641 ( 
.A1(n_595),
.A2(n_386),
.B1(n_393),
.B2(n_514),
.C(n_481),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_598),
.A2(n_514),
.B1(n_492),
.B2(n_386),
.Y(n_642)
);

OAI222xp33_ASAP7_75t_L g643 ( 
.A1(n_592),
.A2(n_406),
.B1(n_539),
.B2(n_532),
.C1(n_491),
.C2(n_517),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_594),
.Y(n_644)
);

OAI221xp5_ASAP7_75t_L g645 ( 
.A1(n_613),
.A2(n_416),
.B1(n_365),
.B2(n_451),
.C(n_449),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_587),
.A2(n_499),
.B1(n_411),
.B2(n_513),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_615),
.A2(n_447),
.B1(n_461),
.B2(n_499),
.Y(n_647)
);

OA21x2_ASAP7_75t_L g648 ( 
.A1(n_631),
.A2(n_605),
.B(n_624),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_597),
.Y(n_649)
);

AO22x1_ASAP7_75t_L g650 ( 
.A1(n_596),
.A2(n_629),
.B1(n_610),
.B2(n_625),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_584),
.A2(n_605),
.B1(n_601),
.B2(n_614),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_593),
.A2(n_499),
.B1(n_521),
.B2(n_561),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_612),
.A2(n_499),
.B1(n_411),
.B2(n_511),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_604),
.A2(n_411),
.B1(n_511),
.B2(n_513),
.Y(n_654)
);

AOI222xp33_ASAP7_75t_L g655 ( 
.A1(n_607),
.A2(n_382),
.B1(n_220),
.B2(n_223),
.C1(n_461),
.C2(n_451),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_606),
.A2(n_521),
.B1(n_561),
.B2(n_517),
.Y(n_656)
);

AOI222xp33_ASAP7_75t_L g657 ( 
.A1(n_599),
.A2(n_382),
.B1(n_220),
.B2(n_223),
.C1(n_366),
.C2(n_411),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_622),
.A2(n_411),
.B1(n_513),
.B2(n_511),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_633),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_596),
.A2(n_366),
.B1(n_491),
.B2(n_516),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_628),
.A2(n_365),
.B(n_412),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_621),
.B(n_516),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_596),
.A2(n_516),
.B1(n_365),
.B2(n_408),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_617),
.A2(n_516),
.B1(n_220),
.B2(n_223),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_617),
.A2(n_220),
.B1(n_223),
.B2(n_432),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_621),
.B(n_220),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_619),
.A2(n_611),
.B1(n_600),
.B2(n_608),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_634),
.B(n_223),
.C(n_220),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_616),
.A2(n_223),
.B1(n_466),
.B2(n_244),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_633),
.A2(n_244),
.B1(n_243),
.B2(n_231),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_618),
.A2(n_244),
.B1(n_243),
.B2(n_231),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_620),
.A2(n_452),
.B1(n_244),
.B2(n_243),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_626),
.A2(n_244),
.B1(n_243),
.B2(n_231),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_627),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_636),
.B(n_633),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_644),
.B(n_632),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_639),
.B(n_609),
.Y(n_677)
);

OAI21xp33_ASAP7_75t_L g678 ( 
.A1(n_651),
.A2(n_667),
.B(n_638),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_649),
.B(n_674),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_662),
.B(n_623),
.Y(n_680)
);

AOI211xp5_ASAP7_75t_L g681 ( 
.A1(n_650),
.A2(n_630),
.B(n_609),
.C(n_55),
.Y(n_681)
);

AOI221xp5_ASAP7_75t_L g682 ( 
.A1(n_641),
.A2(n_243),
.B1(n_231),
.B2(n_244),
.C(n_57),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_R g683 ( 
.A(n_659),
.B(n_52),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_666),
.B(n_53),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_648),
.B(n_56),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_648),
.B(n_60),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_L g687 ( 
.A(n_637),
.B(n_244),
.C(n_243),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_653),
.B(n_243),
.C(n_231),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_652),
.B(n_231),
.C(n_63),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_647),
.A2(n_231),
.B1(n_64),
.B2(n_66),
.Y(n_690)
);

NAND4xp25_ASAP7_75t_L g691 ( 
.A(n_646),
.B(n_635),
.C(n_640),
.D(n_655),
.Y(n_691)
);

AOI221xp5_ASAP7_75t_L g692 ( 
.A1(n_643),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.C(n_69),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_658),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_648),
.B(n_75),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_635),
.B(n_76),
.C(n_78),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_659),
.B(n_79),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_L g697 ( 
.A1(n_668),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_697)
);

OAI221xp5_ASAP7_75t_L g698 ( 
.A1(n_663),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.C(n_88),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_SL g699 ( 
.A1(n_664),
.A2(n_89),
.B(n_90),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_642),
.B(n_91),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_SL g701 ( 
.A1(n_665),
.A2(n_95),
.B(n_96),
.Y(n_701)
);

NAND3xp33_ASAP7_75t_L g702 ( 
.A(n_678),
.B(n_657),
.C(n_654),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_677),
.A2(n_656),
.B1(n_645),
.B2(n_660),
.Y(n_703)
);

NAND3xp33_ASAP7_75t_L g704 ( 
.A(n_682),
.B(n_669),
.C(n_661),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_L g705 ( 
.A(n_698),
.B(n_670),
.C(n_99),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_679),
.B(n_672),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_676),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_680),
.B(n_672),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_681),
.B(n_671),
.C(n_673),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_700),
.B(n_98),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_685),
.B(n_100),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_686),
.B(n_673),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_694),
.B(n_101),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_675),
.B(n_701),
.C(n_690),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_689),
.Y(n_715)
);

NAND4xp75_ASAP7_75t_L g716 ( 
.A(n_692),
.B(n_103),
.C(n_106),
.D(n_107),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_696),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_684),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_707),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_717),
.B(n_683),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_718),
.B(n_683),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_712),
.B(n_699),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_715),
.B(n_688),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_708),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_702),
.B(n_691),
.Y(n_725)
);

XNOR2xp5_ASAP7_75t_L g726 ( 
.A(n_710),
.B(n_703),
.Y(n_726)
);

XOR2x2_ASAP7_75t_L g727 ( 
.A(n_714),
.B(n_695),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_706),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_728),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_719),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_724),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_723),
.Y(n_732)
);

XOR2x2_ASAP7_75t_L g733 ( 
.A(n_726),
.B(n_702),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_732),
.Y(n_734)
);

OAI22x1_ASAP7_75t_L g735 ( 
.A1(n_731),
.A2(n_725),
.B1(n_721),
.B2(n_720),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_729),
.Y(n_736)
);

XNOR2xp5_ASAP7_75t_L g737 ( 
.A(n_733),
.B(n_727),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_731),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_734),
.Y(n_739)
);

OA22x2_ASAP7_75t_L g740 ( 
.A1(n_737),
.A2(n_738),
.B1(n_735),
.B2(n_734),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_736),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_734),
.Y(n_742)
);

AND4x1_ASAP7_75t_L g743 ( 
.A(n_739),
.B(n_725),
.C(n_723),
.D(n_720),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_740),
.A2(n_727),
.B1(n_722),
.B2(n_730),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_744),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_743),
.A2(n_740),
.B1(n_722),
.B2(n_742),
.Y(n_746)
);

AOI221xp5_ASAP7_75t_L g747 ( 
.A1(n_744),
.A2(n_741),
.B1(n_697),
.B2(n_709),
.C(n_704),
.Y(n_747)
);

AO22x2_ASAP7_75t_L g748 ( 
.A1(n_745),
.A2(n_716),
.B1(n_709),
.B2(n_705),
.Y(n_748)
);

AO22x1_ASAP7_75t_L g749 ( 
.A1(n_746),
.A2(n_713),
.B1(n_711),
.B2(n_693),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_747),
.Y(n_750)
);

NOR2x1_ASAP7_75t_L g751 ( 
.A(n_746),
.B(n_722),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_745),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_745),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_752),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_753),
.B(n_722),
.Y(n_755)
);

NOR2x1_ASAP7_75t_L g756 ( 
.A(n_751),
.B(n_697),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_748),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_SL g758 ( 
.A1(n_750),
.A2(n_687),
.B1(n_109),
.B2(n_111),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_748),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_SL g760 ( 
.A1(n_754),
.A2(n_749),
.B(n_113),
.C(n_114),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_755),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_756),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_759),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_757),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_758),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_764),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_763),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_763),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_762),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_761),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_765),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_760),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_764),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_764),
.Y(n_774)
);

AOI22x1_ASAP7_75t_L g775 ( 
.A1(n_772),
.A2(n_108),
.B1(n_115),
.B2(n_116),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_771),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_SL g777 ( 
.A1(n_772),
.A2(n_121),
.B1(n_122),
.B2(n_126),
.Y(n_777)
);

OAI22x1_ASAP7_75t_L g778 ( 
.A1(n_769),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_774),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_766),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_773),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_770),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_778),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_779),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_781),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_777),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_775),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_SL g788 ( 
.A1(n_783),
.A2(n_768),
.B1(n_767),
.B2(n_776),
.Y(n_788)
);

AOI31xp33_ASAP7_75t_L g789 ( 
.A1(n_786),
.A2(n_782),
.A3(n_780),
.B(n_143),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_788),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_790),
.A2(n_787),
.B1(n_784),
.B2(n_785),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_791),
.Y(n_792)
);

AOI221x1_ASAP7_75t_L g793 ( 
.A1(n_792),
.A2(n_789),
.B1(n_142),
.B2(n_144),
.C(n_146),
.Y(n_793)
);

AOI211xp5_ASAP7_75t_L g794 ( 
.A1(n_793),
.A2(n_140),
.B(n_147),
.C(n_148),
.Y(n_794)
);


endmodule