module fake_jpeg_32169_n_472 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_472);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_472;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_53),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_21),
.A2(n_39),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_7),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_6),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_67),
.Y(n_106)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_64),
.B(n_74),
.Y(n_135)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_16),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_20),
.B(n_6),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_85),
.B(n_43),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_20),
.B(n_6),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_16),
.Y(n_90)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_48),
.A2(n_16),
.B1(n_40),
.B2(n_46),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_97),
.A2(n_108),
.B1(n_124),
.B2(n_19),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_98),
.A2(n_111),
.B1(n_120),
.B2(n_146),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_40),
.B1(n_29),
.B2(n_21),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_53),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_34),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_140),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_55),
.A2(n_40),
.B1(n_37),
.B2(n_38),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_57),
.A2(n_40),
.B1(n_39),
.B2(n_29),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_80),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_35),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_141),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_61),
.A2(n_35),
.B1(n_34),
.B2(n_45),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_129),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_83),
.B1(n_66),
.B2(n_76),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_151),
.A2(n_174),
.B1(n_182),
.B2(n_187),
.Y(n_201)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_153),
.Y(n_220)
);

BUFx4f_ASAP7_75t_SL g154 ( 
.A(n_139),
.Y(n_154)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_113),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_160),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_45),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_162),
.B(n_173),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_97),
.A2(n_60),
.B1(n_39),
.B2(n_43),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_171),
.A2(n_185),
.B(n_33),
.Y(n_214)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_106),
.A2(n_71),
.B1(n_89),
.B2(n_86),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_110),
.A2(n_65),
.B1(n_82),
.B2(n_93),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_177),
.A2(n_179),
.B1(n_180),
.B2(n_183),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_101),
.A2(n_54),
.B1(n_56),
.B2(n_92),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_181),
.Y(n_203)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

BUFx8_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_184),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_119),
.A2(n_32),
.B1(n_46),
.B2(n_19),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_120),
.A2(n_32),
.B1(n_19),
.B2(n_33),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_144),
.A2(n_104),
.B1(n_95),
.B2(n_138),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_193),
.B1(n_38),
.B2(n_37),
.Y(n_225)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_22),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_95),
.A2(n_91),
.B1(n_90),
.B2(n_46),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_139),
.B1(n_105),
.B2(n_134),
.Y(n_204)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_204),
.A2(n_221),
.B1(n_206),
.B2(n_224),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_96),
.B1(n_136),
.B2(n_128),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_205),
.A2(n_211),
.B1(n_221),
.B2(n_224),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_182),
.A2(n_123),
.B1(n_134),
.B2(n_116),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_96),
.B1(n_128),
.B2(n_99),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_214),
.B1(n_161),
.B2(n_149),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_136),
.B1(n_127),
.B2(n_125),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_160),
.A2(n_90),
.B(n_33),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_165),
.B(n_155),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_127),
.B1(n_31),
.B2(n_77),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_171),
.A2(n_31),
.B1(n_77),
.B2(n_11),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_157),
.B1(n_148),
.B2(n_176),
.Y(n_256)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_156),
.B(n_159),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_231),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_156),
.B(n_38),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_150),
.B(n_22),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_38),
.C(n_37),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_235),
.B(n_239),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_185),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_236),
.B(n_240),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_237),
.A2(n_256),
.B(n_217),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_214),
.A2(n_170),
.B1(n_164),
.B2(n_167),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_201),
.A2(n_166),
.B1(n_147),
.B2(n_152),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_193),
.B1(n_189),
.B2(n_188),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_243),
.A2(n_254),
.B1(n_262),
.B2(n_195),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_230),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_250),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_216),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_245),
.Y(n_301)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_169),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_248),
.C(n_257),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_199),
.B(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_153),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_251),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_154),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_200),
.B(n_154),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_168),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_259),
.Y(n_295)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_255),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_203),
.B(n_184),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_201),
.A2(n_205),
.B1(n_226),
.B2(n_204),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_209),
.A2(n_183),
.B1(n_175),
.B2(n_31),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_260),
.A2(n_261),
.B1(n_265),
.B2(n_216),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_211),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_196),
.A2(n_22),
.B1(n_184),
.B2(n_37),
.Y(n_262)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_207),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_268),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_197),
.A2(n_38),
.B1(n_22),
.B2(n_2),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_269),
.B(n_272),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_271),
.A2(n_289),
.B(n_294),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_249),
.B(n_244),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_235),
.A2(n_197),
.B1(n_212),
.B2(n_218),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_273),
.A2(n_279),
.B1(n_285),
.B2(n_254),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_267),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_274),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_236),
.B(n_212),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_275),
.B(n_282),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_253),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_277),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_242),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_233),
.B(n_208),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_241),
.B(n_197),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_283),
.B(n_248),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_234),
.A2(n_218),
.B1(n_227),
.B2(n_202),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_234),
.A2(n_213),
.B(n_227),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_287),
.A2(n_210),
.B(n_194),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_288),
.A2(n_245),
.B1(n_268),
.B2(n_255),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g289 ( 
.A1(n_241),
.A2(n_208),
.B(n_229),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_237),
.A2(n_229),
.B(n_222),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_233),
.B(n_202),
.Y(n_298)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_299),
.A2(n_22),
.B1(n_38),
.B2(n_2),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_247),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_311),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_305),
.B(n_330),
.Y(n_358)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_270),
.Y(n_307)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

OA22x2_ASAP7_75t_L g335 ( 
.A1(n_308),
.A2(n_272),
.B1(n_283),
.B2(n_294),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_279),
.A2(n_259),
.B1(n_238),
.B2(n_240),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_338)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_290),
.B(n_298),
.Y(n_311)
);

AO22x1_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_238),
.B1(n_246),
.B2(n_258),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_289),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_296),
.A2(n_262),
.B(n_264),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_313),
.A2(n_285),
.B(n_289),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_293),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_329),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_295),
.A2(n_261),
.B1(n_260),
.B2(n_252),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_315),
.A2(n_316),
.B1(n_333),
.B2(n_285),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_295),
.A2(n_299),
.B1(n_286),
.B2(n_277),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_271),
.A2(n_245),
.B1(n_216),
.B2(n_195),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_296),
.A2(n_273),
.B1(n_287),
.B2(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_321),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_296),
.A2(n_265),
.B(n_263),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_322),
.A2(n_332),
.B(n_287),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_273),
.A2(n_222),
.B1(n_220),
.B2(n_210),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_325),
.A2(n_278),
.B1(n_286),
.B2(n_301),
.Y(n_342)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_280),
.Y(n_327)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_266),
.C(n_257),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_293),
.B(n_220),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_SL g352 ( 
.A1(n_331),
.A2(n_301),
.B(n_284),
.C(n_281),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_294),
.A2(n_6),
.B(n_12),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_335),
.B(n_336),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_337),
.A2(n_339),
.B(n_350),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_341),
.A2(n_356),
.B1(n_361),
.B2(n_362),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_344),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_323),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_282),
.Y(n_345)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

AOI22x1_ASAP7_75t_L g349 ( 
.A1(n_318),
.A2(n_289),
.B1(n_275),
.B2(n_281),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_352),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_320),
.A2(n_297),
.B(n_284),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_328),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_353),
.B(n_359),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_320),
.A2(n_280),
.B(n_302),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_357),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_316),
.A2(n_274),
.B1(n_291),
.B2(n_302),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_313),
.A2(n_331),
.B(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_307),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_327),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_315),
.A2(n_291),
.B1(n_292),
.B2(n_300),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_304),
.A2(n_292),
.B1(n_300),
.B2(n_2),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_324),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_363),
.B(n_326),
.Y(n_366)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_366),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_314),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_374),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_303),
.C(n_311),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_372),
.C(n_375),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_345),
.B(n_326),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_369),
.B(n_378),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_305),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_383),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_329),
.C(n_330),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_308),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_304),
.C(n_325),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_343),
.B(n_292),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_335),
.B(n_319),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_385),
.C(n_388),
.Y(n_400)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_382),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_312),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_362),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_336),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_335),
.B(n_309),
.C(n_321),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_R g386 ( 
.A(n_352),
.B(n_332),
.Y(n_386)
);

FAx1_ASAP7_75t_SL g407 ( 
.A(n_386),
.B(n_352),
.CI(n_349),
.CON(n_407),
.SN(n_407)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_346),
.B(n_310),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_387),
.A2(n_355),
.B1(n_359),
.B2(n_347),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_312),
.Y(n_388)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_389),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_373),
.A2(n_354),
.B(n_339),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_373),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_365),
.A2(n_338),
.B1(n_341),
.B2(n_335),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_391),
.A2(n_405),
.B1(n_406),
.B2(n_408),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_401),
.Y(n_410)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_377),
.Y(n_399)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_399),
.Y(n_423)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_379),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_360),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_403),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_370),
.A2(n_361),
.B1(n_351),
.B2(n_347),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_349),
.C(n_337),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_375),
.C(n_372),
.Y(n_414)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

FAx1_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_380),
.CI(n_383),
.CON(n_419),
.SN(n_419)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

XNOR2x1_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_411),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_368),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_400),
.C(n_404),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_395),
.B(n_385),
.C(n_374),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_424),
.C(n_400),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_391),
.A2(n_386),
.B1(n_364),
.B2(n_365),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_416),
.B(n_417),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_408),
.A2(n_381),
.B(n_388),
.Y(n_417)
);

BUFx24_ASAP7_75t_SL g418 ( 
.A(n_399),
.Y(n_418)
);

BUFx24_ASAP7_75t_SL g425 ( 
.A(n_418),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_419),
.B(n_420),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_405),
.A2(n_352),
.B1(n_351),
.B2(n_371),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_406),
.A2(n_401),
.B1(n_394),
.B2(n_396),
.Y(n_422)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_422),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_300),
.C(n_1),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_392),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_429),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_397),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_415),
.B(n_398),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_431),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_396),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_433),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_423),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_438),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_402),
.C(n_390),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_412),
.C(n_420),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_410),
.B(n_394),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_407),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_426),
.A2(n_413),
.B1(n_421),
.B2(n_409),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_450),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_445),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_434),
.A2(n_389),
.B(n_419),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_441),
.B(n_440),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_449),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_427),
.A2(n_417),
.B(n_419),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_443),
.A2(n_448),
.B(n_8),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_438),
.A2(n_407),
.B(n_11),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_436),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_425),
.A2(n_8),
.B1(n_9),
.B2(n_3),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_451),
.A2(n_452),
.B(n_450),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_444),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_457),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_0),
.C(n_1),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_0),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_458),
.B(n_3),
.C(n_4),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_SL g459 ( 
.A1(n_451),
.A2(n_439),
.B(n_449),
.C(n_447),
.Y(n_459)
);

AOI21x1_ASAP7_75t_L g466 ( 
.A1(n_459),
.A2(n_460),
.B(n_453),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_461),
.B(n_463),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_3),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_462),
.B(n_455),
.Y(n_465)
);

AO21x1_ASAP7_75t_L g468 ( 
.A1(n_465),
.A2(n_4),
.B(n_5),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_466),
.A2(n_3),
.B(n_4),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_467),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_464),
.C(n_468),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_470),
.B(n_5),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_5),
.Y(n_472)
);


endmodule