module fake_jpeg_373_n_435 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_435);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_435;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_43),
.B(n_56),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2x1_ASAP7_75t_SL g92 ( 
.A(n_55),
.B(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_26),
.B(n_14),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_8),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_77),
.Y(n_103)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_76),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_34),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_80),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_82),
.Y(n_128)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

NAND2x1_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_38),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_33),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_85),
.B(n_87),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_33),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_37),
.B1(n_30),
.B2(n_42),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_90),
.A2(n_123),
.B1(n_44),
.B2(n_53),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_104),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_46),
.A2(n_29),
.B1(n_41),
.B2(n_35),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_28),
.B1(n_39),
.B2(n_15),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_47),
.B(n_15),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_49),
.A2(n_24),
.B1(n_36),
.B2(n_38),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_126),
.B1(n_129),
.B2(n_29),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_122),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_57),
.A2(n_30),
.B1(n_15),
.B2(n_42),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_50),
.A2(n_34),
.B1(n_24),
.B2(n_36),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_62),
.A2(n_24),
.B1(n_36),
.B2(n_38),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_26),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_41),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_35),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_133),
.B(n_140),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_134),
.A2(n_147),
.B1(n_149),
.B2(n_174),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g199 ( 
.A1(n_135),
.A2(n_143),
.B1(n_167),
.B2(n_145),
.Y(n_199)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_136),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_85),
.C(n_87),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_158),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_91),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_86),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_142),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_67),
.B1(n_75),
.B2(n_76),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_143),
.A2(n_109),
.B1(n_100),
.B2(n_121),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_103),
.A2(n_69),
.B1(n_60),
.B2(n_34),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_152),
.B1(n_168),
.B2(n_172),
.Y(n_179)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_42),
.B1(n_44),
.B2(n_53),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_54),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_94),
.A2(n_36),
.B1(n_38),
.B2(n_79),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_48),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_39),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_159),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_92),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_169),
.Y(n_201)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_164),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g165 ( 
.A(n_120),
.B(n_48),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_114),
.C(n_52),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_28),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_176),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_102),
.A2(n_120),
.B1(n_115),
.B2(n_118),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_92),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_88),
.B(n_70),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_82),
.B1(n_81),
.B2(n_78),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_175),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_88),
.A2(n_74),
.B1(n_61),
.B2(n_58),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_93),
.B(n_0),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_86),
.B(n_52),
.C(n_112),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_184),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_180),
.B(n_203),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_151),
.B(n_96),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_132),
.A2(n_127),
.B1(n_118),
.B2(n_111),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_189),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_86),
.B(n_100),
.C(n_93),
.Y(n_190)
);

BUFx24_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_159),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_135),
.A2(n_127),
.B1(n_111),
.B2(n_98),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_213),
.B1(n_215),
.B2(n_218),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_145),
.A2(n_167),
.B1(n_151),
.B2(n_137),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_138),
.A2(n_121),
.B1(n_117),
.B2(n_113),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_139),
.A2(n_96),
.B(n_113),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_210),
.A2(n_156),
.B(n_141),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_144),
.A2(n_107),
.B1(n_45),
.B2(n_31),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_117),
.B1(n_112),
.B2(n_93),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_146),
.B(n_112),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_201),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_165),
.A2(n_31),
.B1(n_16),
.B2(n_21),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_153),
.B1(n_164),
.B2(n_161),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_168),
.A2(n_31),
.B1(n_16),
.B2(n_21),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_154),
.A2(n_16),
.B1(n_31),
.B2(n_21),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_201),
.A2(n_154),
.B1(n_152),
.B2(n_175),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_220),
.A2(n_227),
.B(n_237),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_165),
.C(n_154),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_221),
.B(n_180),
.C(n_214),
.Y(n_267)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_222),
.Y(n_283)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

INVx2_ASAP7_75t_R g227 ( 
.A(n_192),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_180),
.Y(n_268)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_231),
.A2(n_239),
.B1(n_246),
.B2(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_142),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_232),
.B(n_233),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_171),
.C(n_155),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_178),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_238),
.B(n_242),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_162),
.B1(n_173),
.B2(n_163),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_197),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_148),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_243),
.A2(n_249),
.B1(n_251),
.B2(n_188),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_248),
.Y(n_263)
);

OAI22x1_ASAP7_75t_SL g245 ( 
.A1(n_179),
.A2(n_136),
.B1(n_157),
.B2(n_31),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_247),
.B1(n_250),
.B2(n_192),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_204),
.A2(n_31),
.B1(n_21),
.B2(n_3),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_179),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_250)
);

INVx11_ASAP7_75t_L g251 ( 
.A(n_186),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_10),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_253),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_183),
.B(n_10),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_210),
.A2(n_183),
.B(n_214),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_190),
.B(n_198),
.Y(n_280)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_190),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_196),
.A2(n_0),
.B1(n_1),
.B2(n_7),
.Y(n_257)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_259),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_239),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_260),
.B(n_279),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_195),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_261),
.B(n_268),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_272),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_270),
.C(n_271),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_221),
.B(n_216),
.C(n_177),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_205),
.C(n_215),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_205),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_203),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_275),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_224),
.A2(n_185),
.B1(n_213),
.B2(n_218),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_224),
.A2(n_203),
.B1(n_202),
.B2(n_189),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_281),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_225),
.B(n_217),
.C(n_198),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_285),
.C(n_286),
.Y(n_300)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_238),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_280),
.A2(n_236),
.B(n_228),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_203),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_225),
.B(n_203),
.C(n_194),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_191),
.C(n_181),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_212),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_220),
.Y(n_305)
);

AO21x2_ASAP7_75t_L g288 ( 
.A1(n_237),
.A2(n_208),
.B(n_182),
.Y(n_288)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_245),
.A2(n_208),
.B1(n_206),
.B2(n_188),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_289),
.A2(n_231),
.B1(n_235),
.B2(n_256),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_227),
.B(n_206),
.C(n_1),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_247),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_317),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_258),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_301),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_272),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_299),
.B(n_306),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_274),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_303),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_305),
.B(n_270),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_263),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_280),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_308),
.B(n_284),
.Y(n_347)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_227),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_312),
.C(n_316),
.Y(n_345)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_311),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_261),
.B(n_222),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_313),
.A2(n_288),
.B(n_236),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_315),
.A2(n_321),
.B1(n_276),
.B2(n_275),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_268),
.B(n_230),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_282),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_269),
.A2(n_228),
.B(n_236),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_259),
.Y(n_323)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_291),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_320),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_264),
.A2(n_236),
.B1(n_226),
.B2(n_250),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_323),
.A2(n_313),
.B(n_319),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_301),
.A2(n_262),
.B1(n_271),
.B2(n_288),
.Y(n_324)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_267),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_327),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_295),
.A2(n_288),
.B1(n_289),
.B2(n_273),
.Y(n_326)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_241),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_329),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_330),
.A2(n_332),
.B1(n_304),
.B2(n_302),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_321),
.A2(n_269),
.B1(n_285),
.B2(n_281),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_286),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_341),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_303),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_339),
.Y(n_364)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_298),
.B(n_277),
.CI(n_290),
.CON(n_336),
.SN(n_336)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_310),
.Y(n_368)
);

AO22x1_ASAP7_75t_L g338 ( 
.A1(n_293),
.A2(n_318),
.B1(n_308),
.B2(n_315),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_314),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_298),
.B(n_233),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_340),
.A2(n_304),
.B(n_314),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_288),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_302),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_344),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_318),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_346),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_347),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_345),
.B(n_300),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_358),
.Y(n_383)
);

A2O1A1Ixp33_ASAP7_75t_SL g370 ( 
.A1(n_354),
.A2(n_367),
.B(n_323),
.C(n_338),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_300),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_325),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_359),
.B(n_366),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_360),
.A2(n_330),
.B1(n_332),
.B2(n_305),
.Y(n_369)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_362),
.Y(n_385)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_293),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_363),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_316),
.Y(n_366)
);

AOI21xp33_ASAP7_75t_L g375 ( 
.A1(n_368),
.A2(n_336),
.B(n_323),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_369),
.A2(n_372),
.B1(n_374),
.B2(n_376),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_373),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_328),
.C(n_341),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_381),
.C(n_379),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_355),
.A2(n_338),
.B1(n_297),
.B2(n_334),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_265),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_365),
.A2(n_346),
.B1(n_334),
.B2(n_340),
.Y(n_374)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_350),
.A2(n_297),
.B1(n_322),
.B2(n_343),
.Y(n_376)
);

A2O1A1Ixp33_ASAP7_75t_SL g377 ( 
.A1(n_354),
.A2(n_343),
.B(n_309),
.C(n_311),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_377),
.A2(n_357),
.B1(n_322),
.B2(n_363),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_352),
.C(n_349),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_364),
.A2(n_322),
.B1(n_337),
.B2(n_320),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_382),
.A2(n_348),
.B1(n_360),
.B2(n_367),
.Y(n_389)
);

XNOR2x1_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_356),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_387),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_389),
.A2(n_391),
.B1(n_392),
.B2(n_394),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_394),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_384),
.A2(n_351),
.B1(n_368),
.B2(n_294),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_385),
.A2(n_336),
.B1(n_356),
.B2(n_349),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_370),
.A2(n_366),
.B(n_265),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g395 ( 
.A(n_370),
.B(n_292),
.CI(n_291),
.CON(n_395),
.SN(n_395)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_397),
.Y(n_405)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_380),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_398),
.B(n_383),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_383),
.C(n_398),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_399),
.B(n_403),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_401),
.B(n_402),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_393),
.B(n_371),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_379),
.C(n_370),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_223),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_406),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_292),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_408),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_388),
.A2(n_377),
.B1(n_257),
.B2(n_251),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_377),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_410),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_388),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_234),
.Y(n_422)
);

A2O1A1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_405),
.A2(n_377),
.B(n_390),
.C(n_395),
.Y(n_413)
);

AOI321xp33_ASAP7_75t_SL g425 ( 
.A1(n_413),
.A2(n_9),
.A3(n_13),
.B1(n_7),
.B2(n_8),
.C(n_12),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_400),
.A2(n_397),
.B(n_392),
.Y(n_414)
);

AO21x1_ASAP7_75t_L g423 ( 
.A1(n_414),
.A2(n_416),
.B(n_419),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_410),
.A2(n_395),
.B1(n_249),
.B2(n_243),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_403),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_421),
.Y(n_427)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_400),
.C(n_240),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_422),
.B(n_424),
.Y(n_430)
);

AND2x2_ASAP7_75t_SL g424 ( 
.A(n_412),
.B(n_9),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_425),
.A2(n_426),
.B(n_11),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_SL g426 ( 
.A(n_418),
.B(n_9),
.Y(n_426)
);

A2O1A1O1Ixp25_ASAP7_75t_L g428 ( 
.A1(n_423),
.A2(n_413),
.B(n_415),
.C(n_419),
.D(n_426),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_429),
.C(n_11),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_427),
.B(n_11),
.C(n_12),
.Y(n_431)
);

OAI321xp33_ASAP7_75t_L g433 ( 
.A1(n_431),
.A2(n_432),
.A3(n_430),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_13),
.C(n_0),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_1),
.Y(n_435)
);


endmodule