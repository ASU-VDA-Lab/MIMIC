module real_jpeg_19051_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_281, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_281;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_249;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_258;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_0),
.A2(n_3),
.B1(n_18),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_0),
.A2(n_5),
.B1(n_54),
.B2(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_3),
.B1(n_18),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_1),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_1),
.A2(n_5),
.B1(n_30),
.B2(n_65),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_2),
.A2(n_3),
.B1(n_18),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_5),
.B1(n_50),
.B2(n_65),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_50),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_23),
.B(n_27),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_2),
.B(n_28),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_2),
.A2(n_5),
.B(n_10),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_2),
.B(n_37),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_2),
.A2(n_40),
.B(n_41),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_3),
.A2(n_7),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_3),
.A2(n_24),
.B(n_50),
.C(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_4),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_10),
.B1(n_63),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_5),
.A2(n_7),
.B1(n_19),
.B2(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_5),
.B(n_92),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_7),
.A2(n_19),
.B1(n_39),
.B2(n_40),
.Y(n_218)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_9),
.A2(n_18),
.B(n_22),
.C(n_25),
.Y(n_21)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_9),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_274),
.B(n_277),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_67),
.B(n_273),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_31),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_15),
.B(n_31),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_15),
.B(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_15),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_17),
.A2(n_25),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_20),
.A2(n_28),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_21),
.B(n_25),
.Y(n_237)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_38),
.B(n_41),
.C(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_41),
.Y(n_45)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_27),
.A2(n_42),
.B(n_50),
.C(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_28),
.A2(n_48),
.B(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_29),
.B(n_237),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_32),
.B(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_32),
.B(n_271),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_46),
.CI(n_51),
.CON(n_32),
.SN(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_37),
.B1(n_43),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_36),
.B(n_97),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_37),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_38),
.A2(n_44),
.B1(n_97),
.B2(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_38),
.A2(n_250),
.B(n_251),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_40),
.A2(n_50),
.B(n_63),
.C(n_139),
.Y(n_138)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_50),
.B(n_85),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_50),
.B(n_64),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.C(n_58),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_52),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_52),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_52),
.B(n_106),
.C(n_107),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_52),
.A2(n_94),
.B1(n_105),
.B2(n_118),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_52),
.B(n_94),
.C(n_213),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_52),
.A2(n_105),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_55),
.B(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_56),
.A2(n_58),
.B1(n_248),
.B2(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_56),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_57),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_58),
.A2(n_248),
.B1(n_249),
.B2(n_252),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_58),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_66),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_61),
.A2(n_64),
.B1(n_79),
.B2(n_82),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_61),
.A2(n_64),
.B1(n_66),
.B2(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_64),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_65),
.B(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_270),
.B(n_272),
.Y(n_67)
);

OAI321xp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_243),
.A3(n_263),
.B1(n_268),
.B2(n_269),
.C(n_281),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_226),
.B(n_242),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_207),
.B(n_225),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_128),
.B(n_188),
.C(n_206),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_113),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_73),
.B(n_113),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_101),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_93),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_75),
.B(n_93),
.C(n_101),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_83),
.B2(n_84),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_76),
.A2(n_77),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_76),
.A2(n_77),
.B1(n_94),
.B2(n_118),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_76),
.B(n_84),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_77),
.B(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_77),
.B(n_94),
.C(n_161),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B(n_81),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_81),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_84)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_85),
.B(n_91),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_85),
.A2(n_86),
.B1(n_91),
.B2(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_112),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_88),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_91),
.B1(n_92),
.B2(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_98),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_96),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_100),
.A2(n_115),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_100),
.B(n_200),
.C(n_202),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_100),
.A2(n_115),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_100),
.A2(n_115),
.B1(n_257),
.B2(n_261),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_123),
.C(n_125),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_103),
.A2(n_106),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_103),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_103),
.B(n_232),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_145),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_121),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_153),
.C(n_156),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_120),
.C(n_122),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_114),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_115),
.B(n_248),
.C(n_252),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_115),
.B(n_261),
.C(n_262),
.Y(n_271)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_120),
.B(n_122),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_135),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_187),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_182),
.B(n_186),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_170),
.B(n_181),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_158),
.B(n_169),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_148),
.B(n_157),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_140),
.B(n_147),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_136),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_144),
.B(n_146),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_150),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_156),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_156),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_173),
.C(n_180),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_156),
.B(n_196),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_160),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_164),
.B1(n_165),
.B2(n_167),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_164),
.B(n_167),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_171),
.B(n_172),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_178),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_179),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_184),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_190),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_204),
.B2(n_205),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_198),
.B2(n_199),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_199),
.C(n_205),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_204),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_209),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_224),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_216),
.C(n_224),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_221),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_221),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_236),
.B(n_239),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_228),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_240),
.B2(n_241),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_234),
.C(n_241),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_245),
.C(n_253),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_245),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_236),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_240),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_255),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_249),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_253),
.A2(n_254),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_266),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);


endmodule