module fake_jpeg_3691_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx12f_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_0),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_40),
.B1(n_46),
.B2(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_62),
.B1(n_59),
.B2(n_53),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_71),
.B1(n_50),
.B2(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_48),
.B1(n_41),
.B2(n_45),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_49),
.B1(n_44),
.B2(n_47),
.Y(n_91)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_41),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_81),
.Y(n_102)
);

INVx5_ASAP7_75t_SL g80 ( 
.A(n_65),
.Y(n_80)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_45),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_48),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

BUFx2_ASAP7_75t_SL g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_67),
.B1(n_66),
.B2(n_46),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_91),
.B1(n_75),
.B2(n_82),
.Y(n_110)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_47),
.B(n_2),
.C(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_74),
.Y(n_108)
);

AOI22x1_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_57),
.B1(n_19),
.B2(n_20),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_16),
.B1(n_38),
.B2(n_37),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_82),
.B1(n_77),
.B2(n_74),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_108),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_114),
.B1(n_120),
.B2(n_9),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_1),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_117),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_96),
.B(n_102),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_5),
.B(n_6),
.Y(n_128)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_39),
.B1(n_36),
.B2(n_34),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_101),
.B1(n_92),
.B2(n_96),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_1),
.B(n_4),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_118),
.Y(n_129)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_123),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

AOI22x1_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_107),
.B1(n_121),
.B2(n_126),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_31),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_128),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_30),
.C(n_26),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_130),
.C(n_18),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_7),
.B(n_8),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_120),
.B1(n_114),
.B2(n_13),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_23),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_139),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_144),
.Y(n_146)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_142),
.B(n_136),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_124),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_149),
.B(n_124),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_152),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_141),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_149),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_153),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_143),
.Y(n_157)
);

AOI321xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_148),
.A3(n_138),
.B1(n_24),
.B2(n_25),
.C(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_10),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_12),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_13),
.B(n_14),
.C(n_135),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_14),
.Y(n_162)
);


endmodule