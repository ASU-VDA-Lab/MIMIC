module fake_jpeg_4141_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_32),
.Y(n_52)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_46),
.Y(n_61)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_57),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_24),
.B1(n_22),
.B2(n_15),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_55),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_24),
.B1(n_15),
.B2(n_22),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_25),
.B1(n_16),
.B2(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_24),
.B1(n_27),
.B2(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_59),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_67),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_69),
.B1(n_19),
.B2(n_18),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_28),
.B1(n_29),
.B2(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_42),
.Y(n_84)
);

NOR2xp67_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_20),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_47),
.B1(n_49),
.B2(n_19),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_49),
.B1(n_60),
.B2(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_67),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_73),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_85),
.B1(n_89),
.B2(n_69),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_46),
.B1(n_55),
.B2(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_91),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_46),
.B1(n_55),
.B2(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_18),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_18),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_102),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_95),
.B1(n_85),
.B2(n_82),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_75),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_94),
.Y(n_123)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx9p33_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_107),
.Y(n_125)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_111),
.Y(n_116)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_9),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_77),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_61),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_113),
.A2(n_63),
.B(n_2),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_81),
.B(n_63),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_112),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_117),
.B1(n_118),
.B2(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_95),
.B1(n_78),
.B2(n_79),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_82),
.B1(n_80),
.B2(n_61),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_120),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_127),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_113),
.A2(n_68),
.B1(n_70),
.B2(n_77),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_129),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_14),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_1),
.C(n_2),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_137),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_127),
.B(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_144),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_108),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_110),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_104),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_158),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_145),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_151),
.C(n_157),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_123),
.C(n_115),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_142),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_98),
.B1(n_109),
.B2(n_114),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_138),
.B1(n_139),
.B2(n_99),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_98),
.B1(n_128),
.B2(n_99),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_131),
.C(n_112),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_102),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_105),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_143),
.C(n_147),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_181)
);

OA21x2_ASAP7_75t_SL g164 ( 
.A1(n_160),
.A2(n_143),
.B(n_144),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_172),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_170),
.C(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_3),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_105),
.C(n_104),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_171),
.A2(n_167),
.B(n_162),
.Y(n_180)
);

OA21x2_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_97),
.B(n_106),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_178),
.C(n_165),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_162),
.A2(n_161),
.B1(n_153),
.B2(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_181),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_150),
.C(n_156),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_170),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_189),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_163),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_176),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_188),
.A2(n_178),
.B(n_166),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_192),
.C(n_195),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_171),
.B1(n_182),
.B2(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_185),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_5),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_8),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_7),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_196),
.A2(n_197),
.B(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_183),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_195),
.B(n_183),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_8),
.B1(n_9),
.B2(n_201),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_9),
.Y(n_203)
);


endmodule