module fake_jpeg_30900_n_534 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_534);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_10),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_53),
.B(n_54),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_22),
.B(n_9),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_57),
.B(n_67),
.Y(n_157)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_59),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_60),
.Y(n_153)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_11),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_11),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_69),
.B(n_77),
.Y(n_139)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_70),
.Y(n_138)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_26),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_81),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_40),
.B(n_11),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_87),
.B(n_92),
.Y(n_148)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_45),
.B(n_11),
.Y(n_92)
);

BUFx4f_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_45),
.B(n_8),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_100),
.Y(n_107)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_20),
.B(n_8),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_106),
.A2(n_108),
.B1(n_109),
.B2(n_121),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_47),
.B1(n_33),
.B2(n_20),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_47),
.B1(n_31),
.B2(n_29),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_31),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_113),
.B(n_124),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_48),
.C(n_44),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_118),
.B(n_13),
.C(n_2),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_50),
.A2(n_48),
.B1(n_41),
.B2(n_44),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_63),
.B(n_29),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_71),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_126),
.A2(n_136),
.B1(n_27),
.B2(n_18),
.Y(n_208)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_95),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_91),
.B(n_41),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_55),
.Y(n_154)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_91),
.B(n_42),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_155),
.B(n_163),
.Y(n_212)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_56),
.Y(n_158)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_70),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_63),
.B(n_52),
.Y(n_164)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx11_ASAP7_75t_L g246 ( 
.A(n_165),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_107),
.B(n_42),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_168),
.B(n_222),
.Y(n_228)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_170),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_104),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_171),
.B(n_195),
.Y(n_233)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_173),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_178),
.Y(n_258)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_117),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_129),
.A2(n_66),
.B1(n_65),
.B2(n_62),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_183),
.A2(n_205),
.B1(n_160),
.B2(n_137),
.Y(n_240)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_102),
.Y(n_184)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_43),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_185),
.B(n_208),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_186),
.Y(n_270)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_187),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_18),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_188),
.B(n_196),
.Y(n_260)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_133),
.Y(n_189)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_189),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_59),
.B1(n_60),
.B2(n_82),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_190),
.A2(n_206),
.B1(n_221),
.B2(n_162),
.Y(n_241)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_191),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_192),
.B(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_193),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_131),
.A2(n_99),
.B1(n_79),
.B2(n_74),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_194),
.A2(n_199),
.B1(n_115),
.B2(n_156),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_145),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_18),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_139),
.B(n_35),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_198),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_126),
.A2(n_90),
.B1(n_72),
.B2(n_58),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_131),
.A2(n_51),
.B1(n_46),
.B2(n_37),
.Y(n_199)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_143),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_161),
.B(n_27),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_202),
.B(n_203),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_125),
.B(n_27),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_73),
.B1(n_78),
.B2(n_93),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_L g206 ( 
.A1(n_144),
.A2(n_80),
.B1(n_30),
.B2(n_27),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_210),
.Y(n_254)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_213),
.B(n_215),
.Y(n_275)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_214),
.A2(n_220),
.B1(n_224),
.B2(n_225),
.Y(n_264)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_153),
.B(n_27),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_103),
.Y(n_231)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g263 ( 
.A(n_217),
.Y(n_263)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_111),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_218),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_106),
.A2(n_27),
.B(n_18),
.C(n_37),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_223),
.Y(n_227)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_120),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g221 ( 
.A1(n_119),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_115),
.B(n_12),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_119),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_140),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_166),
.A2(n_159),
.B1(n_146),
.B2(n_122),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_230),
.A2(n_241),
.B1(n_4),
.B2(n_6),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_231),
.B(n_253),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_234),
.A2(n_199),
.B1(n_194),
.B2(n_187),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_128),
.B1(n_160),
.B2(n_137),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_236),
.A2(n_240),
.B1(n_206),
.B2(n_214),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_177),
.B(n_156),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_242),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_200),
.B(n_132),
.Y(n_242)
);

CKINVDCx12_ASAP7_75t_R g245 ( 
.A(n_182),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_145),
.B(n_3),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_247),
.B(n_250),
.Y(n_302)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_138),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_138),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_197),
.B(n_152),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_265),
.Y(n_281)
);

OA22x2_ASAP7_75t_L g259 ( 
.A1(n_198),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_SL g303 ( 
.A1(n_259),
.A2(n_4),
.B(n_14),
.C(n_15),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_190),
.B(n_132),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_172),
.B(n_162),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_225),
.C(n_217),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_176),
.B(n_0),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_180),
.B(n_0),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_277),
.B(n_285),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_279),
.B(n_318),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_236),
.A2(n_165),
.B1(n_204),
.B2(n_173),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_280),
.A2(n_229),
.B1(n_232),
.B2(n_248),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_183),
.B1(n_167),
.B2(n_169),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_282),
.A2(n_299),
.B1(n_312),
.B2(n_240),
.Y(n_324)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_260),
.B(n_181),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_284),
.B(n_291),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_233),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_289),
.Y(n_330)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

OAI32xp33_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_205),
.A3(n_201),
.B1(n_211),
.B2(n_179),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_290),
.B(n_296),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_186),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_237),
.A2(n_174),
.B(n_3),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_294),
.A2(n_246),
.B(n_263),
.Y(n_341)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_237),
.A2(n_14),
.B(n_3),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_297),
.A2(n_306),
.B(n_264),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_0),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_298),
.B(n_305),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_259),
.A2(n_4),
.B1(n_6),
.B2(n_14),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_300),
.A2(n_273),
.B1(n_270),
.B2(n_243),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_304),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_303),
.A2(n_241),
.B(n_235),
.C(n_246),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_274),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_231),
.B(n_0),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_15),
.B(n_16),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_228),
.B(n_261),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_307),
.B(n_309),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_253),
.B(n_0),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_308),
.B(n_314),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_257),
.B(n_15),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_256),
.Y(n_310)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_310),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_248),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_311),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_252),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_255),
.B(n_16),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_227),
.B(n_17),
.C(n_244),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_259),
.C(n_268),
.Y(n_326)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_227),
.B(n_17),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_243),
.Y(n_319)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_319),
.Y(n_360)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_258),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_L g338 ( 
.A1(n_320),
.A2(n_235),
.B(n_263),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_321),
.A2(n_322),
.B1(n_324),
.B2(n_341),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_285),
.A2(n_259),
.B1(n_263),
.B2(n_232),
.Y(n_322)
);

XNOR2x1_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_298),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_250),
.C(n_258),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_357),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_329),
.Y(n_379)
);

OA22x2_ASAP7_75t_L g374 ( 
.A1(n_333),
.A2(n_345),
.B1(n_310),
.B2(n_316),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_297),
.A2(n_249),
.B(n_226),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_337),
.A2(n_340),
.B(n_351),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_338),
.A2(n_355),
.B(n_356),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_304),
.A2(n_273),
.B1(n_229),
.B2(n_249),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_339),
.A2(n_347),
.B1(n_350),
.B2(n_358),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_302),
.A2(n_226),
.B(n_251),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_342),
.A2(n_311),
.B1(n_319),
.B2(n_320),
.Y(n_361)
);

AO22x1_ASAP7_75t_L g345 ( 
.A1(n_303),
.A2(n_251),
.B1(n_270),
.B2(n_281),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_284),
.A2(n_281),
.B1(n_302),
.B2(n_305),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_290),
.A2(n_303),
.B1(n_306),
.B2(n_276),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_278),
.A2(n_314),
.B(n_279),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_276),
.A2(n_308),
.B(n_291),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_303),
.A2(n_294),
.B(n_315),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_287),
.C(n_286),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_303),
.A2(n_277),
.B1(n_289),
.B2(n_282),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_361),
.A2(n_394),
.B1(n_360),
.B2(n_353),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_330),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_363),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_287),
.Y(n_364)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_364),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_365),
.B(n_368),
.C(n_346),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_334),
.A2(n_303),
.B1(n_307),
.B2(n_292),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_367),
.A2(n_392),
.B1(n_393),
.B2(n_341),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_312),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_350),
.A2(n_309),
.B1(n_295),
.B2(n_313),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_369),
.A2(n_333),
.B1(n_324),
.B2(n_331),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_339),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_386),
.Y(n_402)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_371),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_283),
.Y(n_372)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_372),
.Y(n_411)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

A2O1A1Ixp33_ASAP7_75t_SL g415 ( 
.A1(n_374),
.A2(n_333),
.B(n_337),
.C(n_329),
.Y(n_415)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_375),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_288),
.Y(n_376)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_376),
.Y(n_424)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_349),
.Y(n_378)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_378),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_348),
.B(n_319),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_380),
.B(n_389),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_330),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_381),
.B(n_384),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_332),
.B(n_293),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_323),
.Y(n_385)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_385),
.Y(n_407)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_354),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_387),
.B(n_352),
.Y(n_419)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_389),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_354),
.Y(n_389)
);

INVx6_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_352),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_334),
.A2(n_335),
.B1(n_345),
.B2(n_358),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_334),
.A2(n_317),
.B1(n_335),
.B2(n_345),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_401),
.A2(n_416),
.B1(n_420),
.B2(n_421),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_408),
.C(n_418),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_405),
.A2(n_413),
.B1(n_374),
.B2(n_362),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_383),
.A2(n_340),
.B(n_356),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_406),
.A2(n_394),
.B(n_390),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_351),
.Y(n_408)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_412),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_392),
.A2(n_326),
.B1(n_347),
.B2(n_333),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_333),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_371),
.Y(n_441)
);

OAI21xp33_ASAP7_75t_SL g431 ( 
.A1(n_415),
.A2(n_422),
.B(n_367),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_377),
.A2(n_366),
.B1(n_369),
.B2(n_370),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_363),
.B(n_331),
.Y(n_417)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_417),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_327),
.C(n_357),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_419),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_366),
.A2(n_332),
.B1(n_325),
.B2(n_355),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_383),
.A2(n_379),
.B1(n_374),
.B2(n_393),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_372),
.Y(n_422)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_423),
.Y(n_436)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_425),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_426),
.A2(n_435),
.B1(n_444),
.B2(n_416),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_376),
.Y(n_429)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_429),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_431),
.A2(n_414),
.B1(n_415),
.B2(n_411),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_364),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_433),
.B(n_439),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_406),
.A2(n_380),
.B(n_362),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_434),
.A2(n_438),
.B(n_441),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_405),
.A2(n_368),
.B1(n_361),
.B2(n_385),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_365),
.C(n_325),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_445),
.C(n_447),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_421),
.A2(n_378),
.B(n_375),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_409),
.Y(n_439)
);

BUFx5_ASAP7_75t_L g440 ( 
.A(n_398),
.Y(n_440)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_440),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_410),
.B(n_373),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_443),
.A2(n_395),
.B1(n_411),
.B2(n_424),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_413),
.A2(n_388),
.B1(n_391),
.B2(n_386),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_353),
.C(n_359),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_359),
.C(n_360),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_448),
.B(n_401),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_398),
.Y(n_449)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_409),
.Y(n_450)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_450),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_395),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_451),
.Y(n_465)
);

XOR2x1_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_434),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_458),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_426),
.A2(n_425),
.B1(n_402),
.B2(n_424),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_456),
.A2(n_460),
.B1(n_464),
.B2(n_471),
.Y(n_478)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_432),
.B(n_402),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_430),
.A2(n_444),
.B1(n_435),
.B2(n_436),
.Y(n_459)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_459),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_436),
.A2(n_397),
.B1(n_399),
.B2(n_400),
.Y(n_461)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_461),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_428),
.A2(n_414),
.B1(n_415),
.B2(n_422),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_412),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_466),
.B(n_470),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_415),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_442),
.A2(n_414),
.B1(n_415),
.B2(n_403),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_407),
.C(n_437),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_472),
.B(n_468),
.C(n_458),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_480),
.C(n_481),
.Y(n_496)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_462),
.Y(n_475)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_475),
.Y(n_492)
);

MAJx2_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_428),
.C(n_446),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_479),
.B(n_453),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_448),
.C(n_450),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_438),
.C(n_427),
.Y(n_481)
);

CKINVDCx14_ASAP7_75t_R g482 ( 
.A(n_469),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_485),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_460),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_484),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_440),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_465),
.B(n_429),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_486),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_427),
.C(n_446),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_488),
.B(n_454),
.C(n_452),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_483),
.A2(n_456),
.B(n_452),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_491),
.B(n_497),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_503),
.Y(n_512)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_480),
.Y(n_498)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_498),
.Y(n_504)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_478),
.Y(n_499)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_499),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_474),
.B(n_455),
.C(n_471),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_502),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_477),
.A2(n_467),
.B(n_441),
.Y(n_501)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_501),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_478),
.A2(n_454),
.B(n_464),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_463),
.Y(n_507)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_507),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_488),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_510),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_473),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_497),
.A2(n_476),
.B1(n_467),
.B2(n_487),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_511),
.B(n_514),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_489),
.Y(n_514)
);

AOI321xp33_ASAP7_75t_L g515 ( 
.A1(n_509),
.A2(n_496),
.A3(n_494),
.B1(n_479),
.B2(n_491),
.C(n_473),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_518),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_496),
.C(n_500),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_489),
.C(n_481),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_519),
.B(n_520),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_514),
.B(n_512),
.C(n_510),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_521),
.B(n_512),
.Y(n_522)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_522),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_516),
.A2(n_513),
.B(n_505),
.Y(n_524)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_524),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_523),
.B(n_525),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_526),
.C(n_517),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_495),
.C(n_463),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_492),
.B(n_502),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_511),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_441),
.B(n_501),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_503),
.Y(n_534)
);


endmodule