module real_jpeg_27079_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_321, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;
input n_321;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_0),
.A2(n_7),
.B1(n_20),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_0),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_106),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_0),
.A2(n_42),
.B1(n_46),
.B2(n_106),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_0),
.A2(n_48),
.B1(n_50),
.B2(n_106),
.Y(n_195)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_2),
.B(n_50),
.Y(n_92)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_2),
.Y(n_97)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_2),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_5),
.A2(n_20),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_20),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_5),
.A2(n_42),
.B1(n_46),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_5),
.B(n_33),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_54),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_42),
.B(n_60),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_5),
.A2(n_45),
.B(n_48),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_5),
.B(n_58),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_6),
.A2(n_7),
.B1(n_20),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_48),
.B1(n_50),
.B2(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_6),
.A2(n_42),
.B1(n_46),
.B2(n_72),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_72),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_7),
.A2(n_11),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_11),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_21),
.B1(n_48),
.B2(n_50),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_11),
.A2(n_21),
.B1(n_42),
.B2(n_46),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_16),
.C(n_282),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_81),
.B(n_317),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_34),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_16),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_29),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_17),
.A2(n_25),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_18),
.B(n_104),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_20),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_23),
.Y(n_24)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_22),
.B(n_31),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_22),
.A2(n_25),
.B(n_31),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_24),
.Y(n_127)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_25),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_26),
.B(n_28),
.Y(n_125)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_27),
.A2(n_58),
.B(n_61),
.C(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_27),
.B(n_59),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_27),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_27),
.A2(n_54),
.B(n_154),
.C(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_29),
.B(n_117),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_35),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_73),
.C(n_75),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_36),
.A2(n_37),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_55),
.C(n_69),
.Y(n_37)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_38),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_38),
.B(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_38),
.B(n_55),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_51),
.B(n_52),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_39),
.A2(n_99),
.B(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_40),
.B(n_53),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_40),
.B(n_100),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_40),
.B(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_46),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_42),
.A2(n_44),
.B(n_54),
.C(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_47),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_47),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_47),
.B(n_53),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_48),
.Y(n_50)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_50),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_51),
.B(n_54),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_51),
.A2(n_166),
.B(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_54),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_64),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_62),
.B(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_57),
.A2(n_65),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_58),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_68),
.Y(n_141)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_63),
.B(n_66),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_66),
.B(n_112),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_66),
.A2(n_259),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_69),
.A2(n_70),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_73),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_73),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_73),
.A2(n_75),
.B1(n_243),
.B2(n_314),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_75),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_76),
.B(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_79),
.B(n_292),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_310),
.B(n_316),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_287),
.A3(n_305),
.B1(n_308),
.B2(n_309),
.C(n_321),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_267),
.B(n_286),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_247),
.B(n_266),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_147),
.B(n_229),
.C(n_246),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_133),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_87),
.B(n_133),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_113),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_102),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_89),
.B(n_102),
.C(n_113),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_90),
.B(n_98),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_93),
.B(n_94),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_92),
.A2(n_96),
.B(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_92),
.B(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_94),
.B(n_194),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_96),
.B(n_146),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_96),
.B(n_195),
.Y(n_200)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_99),
.B(n_176),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_101),
.B(n_164),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.C(n_109),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_105),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_107),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_108),
.B(n_291),
.C(n_295),
.Y(n_304)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_123),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_115),
.B(n_120),
.C(n_123),
.Y(n_244)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_128),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_130),
.B(n_193),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.C(n_139),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_134),
.A2(n_135),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_139),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_141),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_145),
.B(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_228),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_221),
.B(n_227),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_178),
.B(n_220),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_167),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_151),
.B(n_167),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.C(n_162),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_152),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_153),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_157),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_156),
.A2(n_157),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_156),
.B(n_263),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_156),
.A2(n_157),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_157),
.A2(n_278),
.B(n_283),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_161),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_166),
.B(n_175),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_174),
.C(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_215),
.B(n_219),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_196),
.B(n_214),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_181),
.B(n_186),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_191),
.C(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_203),
.B(n_213),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_207),
.B(n_212),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_216),
.B(n_217),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_223),
.Y(n_227)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_231),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_244),
.B2(n_245),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_238),
.C(n_245),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_236),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_248),
.B(n_249),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_265),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_261),
.B2(n_262),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_262),
.C(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_255),
.C(n_258),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_263),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_268),
.B(n_269),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_284),
.B2(n_285),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_277),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_277),
.C(n_285),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B(n_276),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_275),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_289),
.C(n_297),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_276),
.B(n_289),
.CI(n_297),
.CON(n_307),
.SN(n_307)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_298),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_298),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_293),
.B2(n_294),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_290),
.A2(n_291),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_300),
.C(n_304),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_306),
.B(n_307),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_307),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_312),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_313),
.Y(n_315)
);


endmodule