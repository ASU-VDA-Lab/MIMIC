module fake_jpeg_11019_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_45),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_56),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_66),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_19),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_24),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_51),
.A2(n_28),
.B1(n_23),
.B2(n_25),
.Y(n_112)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_14),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_14),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_35),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_32),
.B(n_14),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_24),
.Y(n_69)
);

CKINVDCx10_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_114),
.Y(n_120)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_33),
.B1(n_35),
.B2(n_32),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_73),
.A2(n_100),
.B1(n_110),
.B2(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_79),
.B(n_81),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_34),
.B1(n_37),
.B2(n_26),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_80),
.A2(n_92),
.B1(n_72),
.B2(n_116),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_43),
.B(n_12),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_82),
.B(n_88),
.Y(n_142)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_83),
.B(n_89),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_17),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_26),
.B1(n_36),
.B2(n_28),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_12),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_95),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_44),
.A2(n_26),
.B1(n_40),
.B2(n_36),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_109),
.B1(n_42),
.B2(n_38),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_67),
.A2(n_26),
.B1(n_30),
.B2(n_38),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_26),
.C(n_30),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_39),
.C(n_42),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_29),
.Y(n_130)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_54),
.A2(n_26),
.B1(n_40),
.B2(n_36),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_59),
.A2(n_28),
.B1(n_40),
.B2(n_23),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_69),
.B(n_13),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_13),
.B(n_18),
.Y(n_147)
);

CKINVDCx12_ASAP7_75t_R g113 ( 
.A(n_60),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_113),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_17),
.Y(n_114)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_17),
.B1(n_25),
.B2(n_23),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_118),
.A2(n_134),
.B1(n_137),
.B2(n_139),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_136),
.C(n_138),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_130),
.Y(n_185)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_87),
.A2(n_104),
.B(n_74),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_42),
.B1(n_38),
.B2(n_31),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_31),
.C(n_30),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_31),
.B1(n_27),
.B2(n_21),
.Y(n_139)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_27),
.C(n_21),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_3),
.C(n_4),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_27),
.B1(n_21),
.B2(n_18),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_102),
.B1(n_94),
.B2(n_91),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_18),
.B(n_29),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_86),
.B(n_84),
.C(n_99),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_85),
.A2(n_18),
.B1(n_13),
.B2(n_11),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_145),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_189)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_0),
.B(n_1),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_0),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_0),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_154),
.B(n_1),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_156),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_130),
.B(n_128),
.C(n_154),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_158),
.B(n_170),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_166),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_103),
.B1(n_75),
.B2(n_105),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_164),
.B(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_91),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_168),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_120),
.A2(n_76),
.A3(n_77),
.B1(n_115),
.B2(n_96),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_103),
.B1(n_70),
.B2(n_93),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_94),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_SL g172 ( 
.A(n_120),
.B(n_99),
.C(n_29),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_179),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_124),
.B1(n_138),
.B2(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_175),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_134),
.A2(n_93),
.B1(n_70),
.B2(n_102),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_77),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_76),
.Y(n_179)
);

BUFx4f_ASAP7_75t_SL g180 ( 
.A(n_155),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_129),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_115),
.B1(n_2),
.B2(n_3),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_135),
.B1(n_126),
.B2(n_119),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_189),
.B1(n_125),
.B2(n_152),
.Y(n_204)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_6),
.Y(n_219)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_123),
.C(n_130),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_223),
.C(n_219),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_211),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_167),
.A2(n_144),
.B1(n_141),
.B2(n_139),
.Y(n_202)
);

AOI22x1_ASAP7_75t_L g233 ( 
.A1(n_202),
.A2(n_168),
.B1(n_185),
.B2(n_172),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_208),
.A2(n_215),
.B(n_182),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_167),
.A2(n_140),
.B1(n_119),
.B2(n_132),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_216),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_125),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_127),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_218),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_128),
.B(n_122),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_160),
.A2(n_153),
.B1(n_122),
.B2(n_133),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_157),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_223),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_179),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_174),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_146),
.C(n_7),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_160),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_7),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_193),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_195),
.Y(n_250)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_196),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_231),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_164),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_241),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_246),
.B1(n_204),
.B2(n_201),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_213),
.A2(n_166),
.B1(n_189),
.B2(n_175),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_236),
.A2(n_240),
.B1(n_247),
.B2(n_248),
.Y(n_276)
);

NAND2x1_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_187),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_252),
.B(n_200),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_213),
.A2(n_192),
.B1(n_178),
.B2(n_163),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_191),
.A3(n_184),
.B1(n_176),
.B2(n_173),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_220),
.A2(n_178),
.B1(n_163),
.B2(n_173),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_194),
.A2(n_10),
.B1(n_182),
.B2(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_215),
.A2(n_208),
.B(n_200),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_194),
.A2(n_210),
.B1(n_202),
.B2(n_207),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_197),
.C(n_207),
.Y(n_259)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_257),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_262),
.C(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_221),
.C(n_209),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_228),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_263),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_237),
.B1(n_236),
.B2(n_240),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_212),
.C(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_231),
.A2(n_201),
.B1(n_203),
.B2(n_227),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_271),
.B1(n_232),
.B2(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_275),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_234),
.A2(n_201),
.B1(n_203),
.B2(n_224),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_195),
.C(n_205),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_245),
.C(n_252),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_274),
.A2(n_258),
.B1(n_276),
.B2(n_264),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_282),
.B1(n_288),
.B2(n_266),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_253),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_292),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_281),
.A2(n_276),
.B1(n_258),
.B2(n_268),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_274),
.A2(n_230),
.B1(n_229),
.B2(n_234),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_290),
.C(n_257),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_233),
.C(n_244),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_264),
.A2(n_246),
.B1(n_233),
.B2(n_237),
.Y(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_239),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_305),
.B1(n_307),
.B2(n_237),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_272),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_297),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_262),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_300),
.A2(n_281),
.B1(n_290),
.B2(n_289),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_287),
.B(n_273),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_302),
.Y(n_316)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

XNOR2x2_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_239),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_293),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_268),
.C(n_256),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_286),
.C(n_282),
.Y(n_311)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_312),
.B1(n_309),
.B2(n_306),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_297),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_278),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_315),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

FAx1_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_248),
.CI(n_247),
.CON(n_315),
.SN(n_315)
);

A2O1A1Ixp33_ASAP7_75t_SL g317 ( 
.A1(n_304),
.A2(n_298),
.B(n_302),
.C(n_285),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_307),
.B1(n_284),
.B2(n_279),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_285),
.C(n_284),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_296),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_321),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_327),
.Y(n_332)
);

AO221x1_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_287),
.B1(n_279),
.B2(n_261),
.C(n_267),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_325),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_303),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_300),
.C(n_317),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_314),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_318),
.B1(n_311),
.B2(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_329),
.B(n_330),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_315),
.B1(n_260),
.B2(n_270),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_319),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_319),
.C(n_317),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_337),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_330),
.Y(n_338)
);

AOI322xp5_ASAP7_75t_L g337 ( 
.A1(n_332),
.A2(n_317),
.A3(n_242),
.B1(n_235),
.B2(n_225),
.C1(n_205),
.C2(n_226),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_338),
.A2(n_335),
.B(n_332),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_338),
.B(n_339),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_R g342 ( 
.A(n_341),
.B(n_333),
.C(n_235),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_235),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_203),
.C(n_225),
.Y(n_344)
);


endmodule