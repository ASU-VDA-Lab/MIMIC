module real_jpeg_28535_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_292;
wire n_215;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_293;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_216;
wire n_213;
wire n_179;
wire n_244;
wire n_128;
wire n_133;
wire n_202;
wire n_295;
wire n_138;
wire n_257;
wire n_25;
wire n_217;
wire n_210;
wire n_127;
wire n_206;
wire n_53;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_0),
.A2(n_74),
.B1(n_75),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_0),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_123),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_123),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_0),
.A2(n_45),
.B1(n_48),
.B2(n_123),
.Y(n_244)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_1),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_2),
.A2(n_42),
.B1(n_74),
.B2(n_75),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_3),
.A2(n_55),
.B1(n_74),
.B2(n_75),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_3),
.A2(n_45),
.B1(n_48),
.B2(n_55),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_5),
.A2(n_38),
.B1(n_45),
.B2(n_48),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_7),
.A2(n_74),
.B1(n_75),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_7),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_170),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_170),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_7),
.A2(n_45),
.B1(n_48),
.B2(n_170),
.Y(n_257)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_9),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_70),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_27),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_9),
.A2(n_27),
.B(n_209),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_168),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_9),
.A2(n_45),
.B(n_49),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_9),
.B(n_117),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_9),
.A2(n_86),
.B1(n_89),
.B2(n_257),
.Y(n_260)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_12),
.A2(n_74),
.B1(n_75),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_12),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_149),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_149),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_12),
.A2(n_45),
.B1(n_48),
.B2(n_149),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_13),
.A2(n_36),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_13),
.A2(n_36),
.B1(n_45),
.B2(n_48),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_14),
.Y(n_208)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_15),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_100),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_19),
.B(n_100),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_83),
.B2(n_84),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_56),
.B2(n_57),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_23),
.A2(n_24),
.B(n_39),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_25),
.B(n_67),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_25),
.A2(n_31),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_25),
.A2(n_31),
.B1(n_164),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_25),
.A2(n_31),
.B1(n_193),
.B2(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_28),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_27),
.B(n_71),
.Y(n_182)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_28),
.A2(n_78),
.B1(n_167),
.B2(n_182),
.Y(n_181)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_28),
.A2(n_32),
.A3(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_31),
.B(n_145),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_33),
.B1(n_47),
.B2(n_49),
.Y(n_53)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_33),
.B(n_207),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_33),
.A2(n_47),
.B(n_168),
.C(n_236),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_35),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_50),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_40),
.A2(n_52),
.B(n_217),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_43),
.B(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_52),
.B(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_44),
.A2(n_52),
.B1(n_95),
.B2(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_44),
.A2(n_50),
.B(n_115),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_44),
.A2(n_52),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_44),
.A2(n_52),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_44),
.A2(n_52),
.B1(n_216),
.B2(n_234),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_44),
.B(n_168),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_48),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_52),
.A2(n_61),
.B(n_96),
.Y(n_161)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_68),
.B1(n_81),
.B2(n_82),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_64),
.A2(n_66),
.B(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_64),
.A2(n_178),
.B(n_179),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B(n_76),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_80),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_69),
.A2(n_121),
.B1(n_122),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_69),
.A2(n_121),
.B1(n_148),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_71),
.B(n_75),
.C(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_70),
.B(n_98),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_70),
.A2(n_77),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_75),
.Y(n_78)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_75),
.B(n_168),
.CON(n_167),
.SN(n_167)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_93),
.B(n_97),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_97),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_85),
.A2(n_94),
.B1(n_104),
.B2(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B(n_91),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_86),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_86),
.A2(n_89),
.B1(n_139),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_86),
.A2(n_113),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_86),
.A2(n_249),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_87),
.A2(n_92),
.B(n_141),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_87),
.A2(n_88),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_92),
.Y(n_113)
);

INVx11_ASAP7_75t_L g258 ( 
.A(n_88),
.Y(n_258)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_112),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_90),
.A2(n_110),
.B(n_184),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_94),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_97),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.C(n_106),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_105),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_106),
.A2(n_107),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_116),
.C(n_119),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_109),
.B(n_114),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_119),
.B1(n_120),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B(n_124),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_153),
.B(n_303),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_150),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_129),
.B(n_150),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.C(n_136),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_130),
.A2(n_131),
.B1(n_134),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_134),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_136),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.C(n_146),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_137),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_142),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_143),
.Y(n_293)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_297),
.B(n_302),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_197),
.B(n_283),
.C(n_296),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_185),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_156),
.B(n_185),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_171),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_158),
.B(n_159),
.C(n_171),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_166),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_168),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_180),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_173),
.B(n_177),
.C(n_180),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_183),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_186),
.A2(n_187),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_191),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_196),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_196),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_282),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_275),
.B(n_281),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_227),
.B(n_274),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_218),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_201),
.B(n_218),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_211),
.C(n_214),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_202),
.A2(n_203),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_205),
.Y(n_225)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_225),
.C(n_226),
.Y(n_276)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_268),
.B(n_273),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_245),
.B(n_267),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_230),
.B(n_237),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_232),
.B1(n_235),
.B2(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_244),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_253),
.B(n_266),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_251),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_259),
.B(n_265),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_255),
.B(n_256),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_294),
.B2(n_295),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_291),
.C(n_295),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);


endmodule