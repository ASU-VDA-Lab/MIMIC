module fake_jpeg_25521_n_144 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_45),
.Y(n_47)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_2),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_12),
.Y(n_45)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_24),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_26),
.B1(n_28),
.B2(n_22),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_37),
.B1(n_23),
.B2(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_59),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_15),
.B1(n_28),
.B2(n_17),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_15),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_72),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_86),
.B1(n_63),
.B2(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_73),
.Y(n_99)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_19),
.B(n_25),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g100 ( 
.A(n_81),
.B(n_61),
.C(n_4),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_50),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_57),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_94),
.B(n_81),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_83),
.B(n_74),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_104),
.B1(n_78),
.B2(n_67),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_57),
.Y(n_94)
);

OAI21x1_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_3),
.B(n_5),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_82),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_46),
.B(n_53),
.C(n_50),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_102),
.A2(n_84),
.B1(n_77),
.B2(n_72),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_55),
.B1(n_65),
.B2(n_57),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_113),
.B1(n_89),
.B2(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_73),
.C(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_65),
.B1(n_78),
.B2(n_76),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_47),
.C(n_92),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_101),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_115),
.A2(n_116),
.B(n_102),
.Y(n_119)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_99),
.B(n_96),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_118),
.B(n_121),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_99),
.B(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_122),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_100),
.B(n_94),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_97),
.B(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_10),
.C(n_11),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_126),
.B(n_131),
.Y(n_133)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_132),
.B(n_105),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_108),
.C(n_67),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_128),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_133),
.B1(n_10),
.B2(n_6),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_129),
.B(n_6),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_138),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_139),
.Y(n_144)
);


endmodule