module fake_jpeg_2964_n_99 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_41),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_35),
.B1(n_29),
.B2(n_30),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_32),
.B1(n_28),
.B2(n_40),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_32),
.B1(n_28),
.B2(n_34),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_15),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_56),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_3),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_57),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_42),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_42),
.C(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_5),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_42),
.B1(n_49),
.B2(n_46),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_65),
.B1(n_16),
.B2(n_18),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_42),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_4),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_73),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_5),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_76),
.C(n_11),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_6),
.B(n_7),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_83),
.B1(n_70),
.B2(n_22),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_65),
.C(n_14),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_84),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_13),
.C(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_69),
.C(n_24),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_89),
.C(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_91),
.B(n_20),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_93),
.A2(n_26),
.B(n_92),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_81),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_85),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_85),
.Y(n_99)
);


endmodule