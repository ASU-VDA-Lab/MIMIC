module fake_netlist_5_833_n_467 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_467);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_467;

wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_451;
wire n_408;
wire n_376;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_155;
wire n_423;
wire n_284;
wire n_245;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_275;
wire n_252;
wire n_295;
wire n_330;
wire n_147;
wire n_373;
wire n_307;
wire n_439;
wire n_150;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_186;
wire n_191;
wire n_171;
wire n_153;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_325;
wire n_449;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_457;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_264;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_243;
wire n_183;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_422;
wire n_415;
wire n_355;
wire n_336;
wire n_337;
wire n_430;
wire n_313;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_311;
wire n_208;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_165;
wire n_213;
wire n_342;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_461;
wire n_333;
wire n_309;
wire n_462;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_463;
wire n_239;
wire n_466;
wire n_420;
wire n_310;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_174;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_441;
wire n_450;
wire n_312;
wire n_429;
wire n_345;
wire n_210;
wire n_365;
wire n_176;
wire n_182;
wire n_354;
wire n_237;
wire n_425;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_246;
wire n_179;
wire n_410;
wire n_269;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_202;
wire n_266;
wire n_272;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_426;
wire n_409;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_391;
wire n_434;
wire n_175;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_278;

INVx2_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_30),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_22),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_27),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_9),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_0),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_19),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_18),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_59),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_40),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_107),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_15),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_38),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_53),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_47),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_82),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_21),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_0),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_90),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_123),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_50),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_L g180 ( 
.A(n_73),
.B(n_113),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_28),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_11),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_83),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_24),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_35),
.Y(n_187)
);

INVxp33_ASAP7_75t_SL g188 ( 
.A(n_62),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_100),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_14),
.B(n_91),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_58),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_2),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_78),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_93),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_45),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_71),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_110),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_66),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_3),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_64),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_118),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_1),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_96),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_43),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_97),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_26),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_76),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_16),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_79),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_57),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_141),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_56),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_142),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_1),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_3),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_176),
.B(n_195),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_4),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_4),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_148),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_158),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_149),
.B(n_5),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_150),
.A2(n_152),
.B(n_151),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_157),
.Y(n_236)
);

BUFx8_ASAP7_75t_L g237 ( 
.A(n_163),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_153),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_160),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_155),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_154),
.A2(n_5),
.B(n_6),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_178),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_166),
.B(n_187),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_182),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_177),
.B(n_6),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_161),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_164),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_167),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_168),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_232),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_179),
.B1(n_189),
.B2(n_188),
.Y(n_258)
);

BUFx8_ASAP7_75t_SL g259 ( 
.A(n_249),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_186),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_249),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

OR2x2_ASAP7_75t_SL g266 ( 
.A(n_224),
.B(n_225),
.Y(n_266)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

CKINVDCx8_ASAP7_75t_R g269 ( 
.A(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_227),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_223),
.B(n_169),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_223),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_237),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_248),
.B(n_172),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_172),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_170),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_228),
.A2(n_147),
.B1(n_203),
.B2(n_218),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_219),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_242),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_191),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_235),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_224),
.Y(n_293)
);

NAND3xp33_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_251),
.C(n_225),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_253),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_264),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_269),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_243),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_254),
.Y(n_300)
);

BUFx4f_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_256),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_200),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_245),
.B1(n_237),
.B2(n_247),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_287),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_212),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_267),
.B(n_288),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_226),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_284),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_259),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_217),
.Y(n_321)
);

NAND2xp33_ASAP7_75t_L g322 ( 
.A(n_273),
.B(n_171),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_236),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_268),
.B(n_236),
.Y(n_324)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_263),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_257),
.A2(n_190),
.B1(n_181),
.B2(n_156),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_263),
.A2(n_180),
.B1(n_206),
.B2(n_173),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_265),
.B(n_174),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_265),
.B(n_175),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_330),
.Y(n_332)
);

HAxp5_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_7),
.CON(n_333),
.SN(n_333)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_293),
.A2(n_245),
.B1(n_205),
.B2(n_202),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

OAI21x1_ASAP7_75t_L g336 ( 
.A1(n_292),
.A2(n_215),
.B(n_214),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_300),
.A2(n_298),
.B1(n_321),
.B2(n_331),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_304),
.A2(n_199),
.B1(n_220),
.B2(n_213),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_299),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_L g340 ( 
.A1(n_322),
.A2(n_196),
.B(n_211),
.C(n_210),
.Y(n_340)
);

NOR3xp33_ASAP7_75t_L g341 ( 
.A(n_294),
.B(n_276),
.C(n_208),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_305),
.A2(n_207),
.B(n_201),
.C(n_198),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_297),
.B(n_194),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_308),
.A2(n_185),
.B(n_184),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

AOI222xp33_ASAP7_75t_L g349 ( 
.A1(n_296),
.A2(n_183),
.B1(n_7),
.B2(n_10),
.C1(n_12),
.C2(n_13),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_291),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_328),
.A2(n_8),
.B1(n_20),
.B2(n_23),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_315),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_325),
.B(n_25),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_327),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_323),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_313),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_291),
.Y(n_359)
);

BUFx4f_ASAP7_75t_L g360 ( 
.A(n_324),
.Y(n_360)
);

INVx6_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_326),
.Y(n_362)
);

AND3x1_ASAP7_75t_SL g363 ( 
.A(n_320),
.B(n_33),
.C(n_34),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_325),
.B(n_36),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_L g367 ( 
.A1(n_301),
.A2(n_37),
.B(n_39),
.C(n_42),
.Y(n_367)
);

OAI221xp5_ASAP7_75t_L g368 ( 
.A1(n_337),
.A2(n_338),
.B1(n_349),
.B2(n_342),
.C(n_346),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_301),
.Y(n_369)
);

AO32x2_ASAP7_75t_L g370 ( 
.A1(n_363),
.A2(n_329),
.A3(n_326),
.B1(n_318),
.B2(n_307),
.Y(n_370)
);

OAI21x1_ASAP7_75t_L g371 ( 
.A1(n_336),
.A2(n_318),
.B(n_307),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_350),
.A2(n_316),
.B(n_46),
.Y(n_373)
);

OAI21x1_ASAP7_75t_L g374 ( 
.A1(n_335),
.A2(n_345),
.B(n_352),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_353),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_334),
.A2(n_319),
.B1(n_316),
.B2(n_49),
.Y(n_376)
);

AOI221xp5_ASAP7_75t_L g377 ( 
.A1(n_341),
.A2(n_316),
.B1(n_48),
.B2(n_51),
.C(n_52),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_44),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_343),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_54),
.Y(n_380)
);

OAI221xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_55),
.B1(n_60),
.B2(n_63),
.C(n_65),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_335),
.A2(n_67),
.B(n_68),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_361),
.Y(n_384)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_362),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_332),
.B(n_69),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_351),
.A2(n_70),
.B1(n_72),
.B2(n_75),
.Y(n_388)
);

AO21x2_ASAP7_75t_L g389 ( 
.A1(n_358),
.A2(n_77),
.B(n_84),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_358),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_360),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_356),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_333),
.B(n_104),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_383),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_388),
.A2(n_364),
.B1(n_355),
.B2(n_360),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_375),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_394),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_372),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_371),
.A2(n_365),
.B(n_344),
.Y(n_400)
);

OA21x2_ASAP7_75t_L g401 ( 
.A1(n_374),
.A2(n_367),
.B(n_359),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_368),
.A2(n_340),
.B(n_362),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_105),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_145),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_388),
.A2(n_109),
.B1(n_112),
.B2(n_114),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_376),
.A2(n_115),
.B1(n_117),
.B2(n_119),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_387),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_376),
.A2(n_120),
.B1(n_121),
.B2(n_125),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_382),
.A2(n_126),
.B(n_127),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

OAI321xp33_ASAP7_75t_L g411 ( 
.A1(n_392),
.A2(n_128),
.A3(n_129),
.B1(n_131),
.B2(n_132),
.C(n_134),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_380),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_393),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_397),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_369),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_407),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_378),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_404),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_403),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_378),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_398),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_384),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_402),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_400),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_405),
.A2(n_377),
.B1(n_391),
.B2(n_392),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_401),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_426),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_386),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_408),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_396),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_406),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_415),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_420),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_416),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_405),
.Y(n_437)
);

OAI31xp33_ASAP7_75t_L g438 ( 
.A1(n_425),
.A2(n_412),
.A3(n_381),
.B(n_396),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_417),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_411),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_434),
.B(n_421),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_SL g442 ( 
.A(n_438),
.B(n_412),
.C(n_390),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_389),
.Y(n_443)
);

NAND4xp25_ASAP7_75t_L g444 ( 
.A(n_440),
.B(n_373),
.C(n_411),
.D(n_370),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_439),
.B(n_389),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_370),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_433),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_435),
.Y(n_449)
);

OAI211xp5_ASAP7_75t_SL g450 ( 
.A1(n_449),
.A2(n_438),
.B(n_430),
.C(n_436),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_448),
.B(n_437),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_429),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_451),
.B(n_445),
.Y(n_453)
);

AOI221xp5_ASAP7_75t_L g454 ( 
.A1(n_453),
.A2(n_452),
.B1(n_442),
.B2(n_450),
.C(n_444),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_454),
.A2(n_446),
.B1(n_443),
.B2(n_431),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_455),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_456),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_457),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_458),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_458),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_460),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_461),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_461),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_463),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_462),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_464),
.A2(n_465),
.B(n_459),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_466),
.A2(n_447),
.B1(n_409),
.B2(n_401),
.Y(n_467)
);


endmodule