module fake_jpeg_3324_n_208 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_208);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_11),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_11),
.B(n_47),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_52),
.Y(n_77)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_81),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_62),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_84),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_51),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_71),
.B1(n_72),
.B2(n_58),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_90),
.B1(n_77),
.B2(n_68),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_58),
.B1(n_68),
.B2(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_82),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_67),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_86),
.B1(n_91),
.B2(n_80),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_112),
.B1(n_1),
.B2(n_3),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_101),
.B(n_113),
.Y(n_141)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_75),
.B(n_64),
.C(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_77),
.B1(n_76),
.B2(n_78),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_55),
.B1(n_70),
.B2(n_2),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_57),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_64),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_22),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_60),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_0),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_82),
.C(n_70),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_50),
.C(n_37),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_74),
.B1(n_61),
.B2(n_55),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_135),
.B1(n_117),
.B2(n_6),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_130),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_26),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_10),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_139),
.B1(n_7),
.B2(n_8),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_138),
.B(n_4),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_19),
.B1(n_49),
.B2(n_44),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_103),
.C(n_101),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_149),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_147),
.B1(n_148),
.B2(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_146),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_25),
.B1(n_43),
.B2(n_41),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_161),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_152)
);

NOR4xp25_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_158),
.C(n_159),
.D(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_36),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_150),
.C(n_148),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_12),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_160),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_13),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_18),
.B1(n_14),
.B2(n_16),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_164),
.A2(n_124),
.B1(n_137),
.B2(n_17),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_161),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_168),
.B(n_180),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_16),
.C(n_17),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_147),
.C(n_156),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_185),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_18),
.B1(n_162),
.B2(n_171),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_169),
.B1(n_175),
.B2(n_162),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_170),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_172),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_SL g192 ( 
.A(n_187),
.B(n_174),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_197),
.B(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_196),
.Y(n_201)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_174),
.C(n_166),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_190),
.B(n_191),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_193),
.B1(n_183),
.B2(n_167),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_202),
.A2(n_201),
.B(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_203),
.Y(n_205)
);

AOI31xp67_ASAP7_75t_SL g206 ( 
.A1(n_205),
.A2(n_192),
.A3(n_182),
.B(n_178),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_173),
.B(n_184),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_176),
.Y(n_208)
);


endmodule