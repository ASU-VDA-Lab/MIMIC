module fake_netlist_1_8014_n_30 (n_1, n_2, n_4, n_3, n_5, n_0, n_30);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_6;
wire n_29;
wire n_7;
wire n_27;
CKINVDCx6p67_ASAP7_75t_R g6 ( .A(n_4), .Y(n_6) );
CKINVDCx20_ASAP7_75t_R g7 ( .A(n_3), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_1), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_0), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
INVx2_ASAP7_75t_SL g12 ( .A(n_11), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
CKINVDCx8_ASAP7_75t_R g14 ( .A(n_8), .Y(n_14) );
INVxp67_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_14), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_13), .Y(n_17) );
NAND2xp33_ASAP7_75t_SL g18 ( .A(n_12), .B(n_7), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_17), .B(n_15), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
INVxp67_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_19), .B(n_15), .Y(n_23) );
AOI211xp5_ASAP7_75t_SL g24 ( .A1(n_22), .A2(n_21), .B(n_20), .C(n_6), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVxp33_ASAP7_75t_SL g26 ( .A(n_25), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_25), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_24), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
AOI22xp5_ASAP7_75t_SL g30 ( .A1(n_29), .A2(n_26), .B1(n_28), .B2(n_16), .Y(n_30) );
endmodule