module fake_jpeg_13185_n_625 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_625);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_625;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_15),
.B(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_61),
.B(n_64),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_66),
.B(n_71),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_67),
.Y(n_209)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_72),
.B(n_74),
.Y(n_151)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_73),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_77),
.B(n_79),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_78),
.Y(n_196)
);

INVx2_ASAP7_75t_R g79 ( 
.A(n_19),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_22),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_80),
.B(n_86),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_82),
.Y(n_173)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_83),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_84),
.Y(n_187)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_25),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_24),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_87),
.B(n_93),
.Y(n_176)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_90),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_26),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_97),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_41),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_98),
.B(n_99),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_41),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_101),
.Y(n_213)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_24),
.B(n_2),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_104),
.B(n_109),
.Y(n_199)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_37),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_31),
.B(n_3),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_119),
.B(n_122),
.Y(n_212)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_120),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_42),
.Y(n_124)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

BUFx16f_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

BUFx16f_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_30),
.Y(n_128)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_80),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_132),
.B(n_84),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_76),
.A2(n_32),
.B1(n_82),
.B2(n_60),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_137),
.A2(n_143),
.B(n_117),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_73),
.A2(n_29),
.B1(n_40),
.B2(n_50),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_138),
.A2(n_146),
.B1(n_91),
.B2(n_78),
.Y(n_253)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_142),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_70),
.A2(n_32),
.B1(n_30),
.B2(n_45),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_100),
.A2(n_59),
.B1(n_50),
.B2(n_40),
.Y(n_146)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_156),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_29),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_158),
.B(n_189),
.Y(n_233)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_85),
.A2(n_32),
.B1(n_55),
.B2(n_54),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_164),
.A2(n_183),
.B1(n_143),
.B2(n_176),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_169),
.Y(n_276)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_179),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_79),
.B(n_52),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_188),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_62),
.A2(n_52),
.B1(n_55),
.B2(n_54),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_80),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_126),
.B(n_53),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

INVx6_ASAP7_75t_SL g192 ( 
.A(n_127),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_192),
.Y(n_255)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_193),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_113),
.B(n_58),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_200),
.B(n_6),
.Y(n_269)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_127),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_116),
.B(n_53),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_208),
.B(n_211),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_118),
.B(n_49),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_131),
.A2(n_128),
.B1(n_48),
.B2(n_49),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_215),
.A2(n_242),
.B1(n_268),
.B2(n_284),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_198),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_216),
.B(n_258),
.Y(n_305)
);

CKINVDCx12_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_217),
.Y(n_319)
);

CKINVDCx12_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_218),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_219),
.B(n_245),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_220),
.A2(n_224),
.B1(n_196),
.B2(n_144),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_221),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_48),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_222),
.B(n_265),
.Y(n_308)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_223),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_132),
.A2(n_121),
.B1(n_123),
.B2(n_69),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_95),
.C(n_106),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_225),
.B(n_282),
.C(n_137),
.Y(n_300)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_130),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g329 ( 
.A(n_227),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_229),
.Y(n_307)
);

HAxp5_ASAP7_75t_SL g231 ( 
.A(n_172),
.B(n_120),
.CON(n_231),
.SN(n_231)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_231),
.B(n_234),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_232),
.A2(n_280),
.B(n_140),
.Y(n_314)
);

NAND3xp33_ASAP7_75t_SL g234 ( 
.A(n_145),
.B(n_96),
.C(n_108),
.Y(n_234)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_149),
.Y(n_238)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_239),
.Y(n_327)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_134),
.Y(n_240)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_240),
.Y(n_299)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_141),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_241),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_131),
.A2(n_58),
.B1(n_42),
.B2(n_81),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_153),
.Y(n_243)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_243),
.Y(n_295)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_150),
.Y(n_244)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_244),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_145),
.B(n_58),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_246),
.Y(n_342)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_153),
.Y(n_248)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_249),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_250),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_212),
.A2(n_58),
.B(n_42),
.C(n_6),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_252),
.B(n_254),
.Y(n_333)
);

OA22x2_ASAP7_75t_L g298 ( 
.A1(n_253),
.A2(n_164),
.B1(n_271),
.B2(n_196),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_159),
.B(n_4),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_185),
.Y(n_257)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_159),
.B(n_5),
.Y(n_258)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_170),
.Y(n_259)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_198),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_270),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_176),
.A2(n_94),
.B1(n_63),
.B2(n_7),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_262),
.A2(n_271),
.B1(n_191),
.B2(n_136),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_147),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_173),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_269),
.A2(n_276),
.B1(n_279),
.B2(n_247),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_151),
.B(n_8),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_182),
.A2(n_168),
.B1(n_155),
.B2(n_165),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_139),
.Y(n_272)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_180),
.Y(n_273)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_151),
.B(n_9),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_275),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_199),
.B(n_9),
.Y(n_275)
);

NAND4xp25_ASAP7_75t_L g277 ( 
.A(n_199),
.B(n_9),
.C(n_10),
.D(n_11),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_285),
.Y(n_328)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_135),
.Y(n_278)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_147),
.B(n_9),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_281),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_200),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_166),
.B(n_13),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_169),
.B(n_133),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_167),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_148),
.B(n_14),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_173),
.A2(n_14),
.B1(n_18),
.B2(n_201),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_286),
.A2(n_163),
.B1(n_175),
.B2(n_202),
.Y(n_316)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_152),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_288),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_183),
.B(n_14),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_157),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_289),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_298),
.A2(n_318),
.B1(n_323),
.B2(n_331),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_300),
.B(n_314),
.Y(n_354)
);

AO22x1_ASAP7_75t_L g312 ( 
.A1(n_231),
.A2(n_129),
.B1(n_163),
.B2(n_140),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_312),
.A2(n_335),
.B(n_251),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_317),
.A2(n_321),
.B1(n_343),
.B2(n_344),
.Y(n_381)
);

AO22x1_ASAP7_75t_SL g320 ( 
.A1(n_224),
.A2(n_203),
.B1(n_197),
.B2(n_178),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_320),
.B(n_322),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_283),
.A2(n_184),
.B1(n_195),
.B2(n_206),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_281),
.B(n_195),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_225),
.A2(n_154),
.B1(n_162),
.B2(n_205),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_282),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_339),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_253),
.A2(n_142),
.B1(n_232),
.B2(n_233),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_259),
.A2(n_238),
.B1(n_276),
.B2(n_223),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_332),
.A2(n_346),
.B1(n_250),
.B2(n_264),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_222),
.A2(n_228),
.B(n_282),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_255),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_340),
.B(n_251),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_269),
.A2(n_252),
.B1(n_244),
.B2(n_240),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_269),
.A2(n_237),
.B1(n_230),
.B2(n_260),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_265),
.B(n_280),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_264),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_278),
.A2(n_272),
.B1(n_287),
.B2(n_239),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_330),
.Y(n_349)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_349),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_319),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_366),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_331),
.A2(n_300),
.B1(n_326),
.B2(n_333),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_351),
.A2(n_362),
.B(n_363),
.Y(n_406)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_352),
.Y(n_404)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_302),
.Y(n_353)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_298),
.A2(n_248),
.B1(n_227),
.B2(n_249),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_357),
.A2(n_338),
.B1(n_294),
.B2(n_297),
.Y(n_393)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_317),
.A2(n_284),
.B1(n_221),
.B2(n_243),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_359),
.A2(n_388),
.B1(n_391),
.B2(n_318),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_305),
.B(n_235),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_361),
.B(n_370),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_363),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_295),
.Y(n_364)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

INVx11_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_263),
.Y(n_366)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_347),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_367),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_307),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_373),
.Y(n_412)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_327),
.Y(n_371)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_371),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_323),
.A2(n_235),
.B1(n_236),
.B2(n_256),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_372),
.A2(n_329),
.B1(n_337),
.B2(n_325),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_301),
.Y(n_373)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_297),
.Y(n_374)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_374),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_315),
.B(n_236),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_375),
.B(n_382),
.Y(n_421)
);

INVx4_ASAP7_75t_SL g376 ( 
.A(n_312),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_376),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_377),
.A2(n_387),
.B1(n_392),
.B2(n_341),
.Y(n_395)
);

CKINVDCx12_ASAP7_75t_R g378 ( 
.A(n_312),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_378),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_290),
.B(n_263),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_380),
.Y(n_413)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_293),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_343),
.B(n_256),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_384),
.Y(n_424)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_291),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_322),
.B(n_226),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_301),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_314),
.B(n_226),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_296),
.Y(n_423)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_329),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_313),
.A2(n_250),
.B1(n_321),
.B2(n_333),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_310),
.B(n_315),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_389),
.B(n_390),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_340),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_313),
.A2(n_306),
.B1(n_308),
.B2(n_290),
.Y(n_391)
);

INVx13_ASAP7_75t_L g392 ( 
.A(n_341),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_393),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_394),
.B(n_416),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_395),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_360),
.A2(n_387),
.B1(n_359),
.B2(n_371),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_397),
.A2(n_406),
.B(n_386),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_354),
.B(n_335),
.C(n_308),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_423),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_369),
.A2(n_345),
.B1(n_298),
.B2(n_336),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_410),
.B1(n_417),
.B2(n_427),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_415),
.A2(n_430),
.B1(n_372),
.B2(n_348),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_324),
.Y(n_416)
);

OAI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_369),
.A2(n_298),
.B1(n_320),
.B2(n_342),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_320),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_382),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_386),
.A2(n_292),
.B(n_311),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_422),
.A2(n_358),
.B(n_353),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_354),
.B(n_293),
.C(n_309),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_429),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_348),
.A2(n_329),
.B1(n_294),
.B2(n_342),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_354),
.B(n_375),
.C(n_351),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_381),
.A2(n_309),
.B1(n_303),
.B2(n_296),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_398),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_431),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_398),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_444),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_350),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_435),
.B(n_437),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_436),
.B(n_443),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_403),
.B(n_380),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_407),
.Y(n_438)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_438),
.Y(n_465)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_414),
.Y(n_440)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_440),
.Y(n_469)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_396),
.Y(n_442)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_442),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_415),
.A2(n_390),
.B1(n_362),
.B2(n_370),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_412),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_396),
.Y(n_445)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_445),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_401),
.B(n_349),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_446),
.B(n_461),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_412),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_462),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_418),
.A2(n_360),
.B1(n_355),
.B2(n_381),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_448),
.B(n_449),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_418),
.A2(n_430),
.B1(n_419),
.B2(n_420),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_451),
.A2(n_405),
.B(n_423),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_376),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_457),
.Y(n_472)
);

INVx13_ASAP7_75t_L g453 ( 
.A(n_411),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_453),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_408),
.A2(n_391),
.B1(n_388),
.B2(n_382),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_454),
.A2(n_399),
.B1(n_428),
.B2(n_402),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_416),
.B(n_303),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_455),
.Y(n_487)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_456),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_420),
.A2(n_376),
.B1(n_352),
.B2(n_374),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_458),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_459),
.A2(n_422),
.B(n_437),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_401),
.B(n_377),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_404),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_400),
.B(n_413),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_463),
.B(n_464),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_400),
.B(n_413),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_451),
.A2(n_406),
.B(n_428),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_470),
.B(n_494),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_473),
.B(n_481),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_474),
.A2(n_454),
.B1(n_441),
.B2(n_434),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_439),
.B(n_421),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_489),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_435),
.B(n_411),
.Y(n_477)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_394),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_444),
.B(n_424),
.Y(n_482)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_482),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_427),
.Y(n_484)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_484),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_486),
.A2(n_443),
.B1(n_448),
.B2(n_436),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_439),
.B(n_421),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_489),
.B(n_493),
.C(n_495),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_447),
.B(n_424),
.Y(n_490)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_490),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_426),
.C(n_399),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_456),
.A2(n_407),
.B(n_409),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_409),
.C(n_425),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_446),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_496),
.B(n_464),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_498),
.A2(n_467),
.B1(n_482),
.B2(n_466),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_499),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_506),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_481),
.A2(n_450),
.B1(n_441),
.B2(n_457),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_502),
.A2(n_468),
.B1(n_484),
.B2(n_474),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_471),
.Y(n_504)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_504),
.Y(n_527)
);

NOR2xp67_ASAP7_75t_SL g507 ( 
.A(n_495),
.B(n_461),
.Y(n_507)
);

AOI21xp33_ASAP7_75t_L g545 ( 
.A1(n_507),
.A2(n_513),
.B(n_497),
.Y(n_545)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_475),
.Y(n_510)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_510),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_463),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_511),
.B(n_512),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_452),
.Y(n_512)
);

OA21x2_ASAP7_75t_L g514 ( 
.A1(n_472),
.A2(n_452),
.B(n_432),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_514),
.B(n_492),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_481),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_515),
.B(n_518),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_493),
.B(n_459),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_516),
.B(n_521),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_476),
.B(n_462),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_517),
.B(n_522),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_487),
.B(n_483),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_425),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_520),
.Y(n_526)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_475),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_486),
.B(n_458),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_470),
.B(n_445),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_491),
.B(n_442),
.C(n_438),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_524),
.C(n_465),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_311),
.C(n_325),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_471),
.A2(n_433),
.B1(n_431),
.B2(n_440),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_525),
.A2(n_481),
.B1(n_478),
.B2(n_494),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_528),
.B(n_544),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_483),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_529),
.Y(n_555)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_530),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_531),
.A2(n_536),
.B1(n_539),
.B2(n_410),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_480),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_532),
.B(n_547),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_509),
.B(n_472),
.C(n_480),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_533),
.B(n_535),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_509),
.B(n_468),
.C(n_490),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_498),
.A2(n_502),
.B1(n_505),
.B2(n_508),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_500),
.A2(n_478),
.B1(n_465),
.B2(n_485),
.Y(n_542)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_542),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_467),
.C(n_473),
.Y(n_544)
);

OA21x2_ASAP7_75t_SL g565 ( 
.A1(n_545),
.A2(n_365),
.B(n_479),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_501),
.A2(n_466),
.B(n_477),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_546),
.A2(n_523),
.B(n_524),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_511),
.B(n_328),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_549),
.B(n_488),
.Y(n_558)
);

A2O1A1O1Ixp25_ASAP7_75t_L g550 ( 
.A1(n_533),
.A2(n_512),
.B(n_501),
.C(n_514),
.D(n_522),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_550),
.B(n_543),
.Y(n_577)
);

INVx13_ASAP7_75t_L g551 ( 
.A(n_549),
.Y(n_551)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_551),
.Y(n_571)
);

NOR3xp33_ASAP7_75t_SL g552 ( 
.A(n_537),
.B(n_514),
.C(n_485),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_552),
.B(n_553),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_526),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_554),
.A2(n_534),
.B(n_546),
.Y(n_569)
);

OAI322xp33_ASAP7_75t_L g557 ( 
.A1(n_538),
.A2(n_506),
.A3(n_517),
.B1(n_492),
.B2(n_488),
.C1(n_525),
.C2(n_469),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_557),
.A2(n_565),
.B(n_540),
.Y(n_574)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_558),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_543),
.B(n_469),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_560),
.B(n_548),
.Y(n_580)
);

BUFx12_ASAP7_75t_L g561 ( 
.A(n_528),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_561),
.B(n_541),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_527),
.B(n_479),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_563),
.B(n_542),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_530),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_564),
.A2(n_539),
.B1(n_531),
.B2(n_527),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_567),
.A2(n_479),
.B1(n_364),
.B2(n_453),
.Y(n_583)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_569),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_570),
.B(n_572),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_568),
.B(n_535),
.C(n_534),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_568),
.B(n_541),
.C(n_544),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_573),
.B(n_559),
.C(n_555),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_574),
.B(n_578),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_576),
.B(n_579),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_577),
.A2(n_581),
.B1(n_583),
.B2(n_562),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_560),
.B(n_548),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_553),
.B(n_540),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_580),
.B(n_567),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_554),
.B(n_414),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_582),
.B(n_563),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_585),
.B(n_590),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_575),
.A2(n_558),
.B1(n_562),
.B2(n_564),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_587),
.A2(n_584),
.B1(n_571),
.B2(n_591),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_592),
.B(n_582),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_573),
.B(n_556),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_593),
.B(n_594),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_572),
.B(n_556),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_580),
.B(n_569),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_595),
.B(n_590),
.C(n_589),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_596),
.B(n_597),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_577),
.B(n_561),
.Y(n_597)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_599),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_600),
.B(n_603),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_588),
.B(n_566),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_601),
.B(n_605),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_596),
.B(n_570),
.Y(n_605)
);

AOI31xp67_ASAP7_75t_L g606 ( 
.A1(n_586),
.A2(n_552),
.A3(n_551),
.B(n_550),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_606),
.B(n_607),
.C(n_595),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_586),
.A2(n_566),
.B(n_578),
.Y(n_607)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_608),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_605),
.B(n_561),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_610),
.A2(n_611),
.B(n_613),
.Y(n_616)
);

NAND5xp2_ASAP7_75t_L g611 ( 
.A(n_604),
.B(n_585),
.C(n_453),
.D(n_392),
.E(n_367),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_598),
.B(n_364),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_614),
.A2(n_612),
.B(n_609),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_617),
.B(n_618),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_614),
.A2(n_602),
.B(n_600),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_615),
.B(n_334),
.C(n_338),
.Y(n_620)
);

AO221x1_ASAP7_75t_L g621 ( 
.A1(n_620),
.A2(n_616),
.B1(n_295),
.B2(n_338),
.C(n_334),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_621),
.B(n_619),
.Y(n_622)
);

AO21x1_ASAP7_75t_L g623 ( 
.A1(n_622),
.A2(n_384),
.B(n_291),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_623),
.A2(n_292),
.B(n_304),
.Y(n_624)
);

OAI31xp33_ASAP7_75t_L g625 ( 
.A1(n_624),
.A2(n_299),
.A3(n_304),
.B(n_350),
.Y(n_625)
);


endmodule