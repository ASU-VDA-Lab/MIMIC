module fake_jpeg_24491_n_249 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

AND2x4_ASAP7_75t_SL g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_39),
.B(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_22),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_16),
.B1(n_25),
.B2(n_20),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.Y(n_61)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_24),
.B(n_18),
.C(n_26),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_22),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_25),
.B1(n_17),
.B2(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_62),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_14),
.Y(n_96)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_40),
.A2(n_24),
.B(n_18),
.C(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_20),
.B1(n_17),
.B2(n_27),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_45),
.C(n_50),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_63),
.C(n_60),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_57),
.B1(n_28),
.B2(n_17),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_63),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_58),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_67),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_109),
.Y(n_121)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_104),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_78),
.C(n_77),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_61),
.B1(n_59),
.B2(n_76),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_107),
.B1(n_28),
.B2(n_86),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_80),
.B(n_78),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_113),
.B1(n_95),
.B2(n_92),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_115),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_79),
.A2(n_60),
.B1(n_36),
.B2(n_38),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_108),
.Y(n_122)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_77),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_68),
.B(n_46),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx2_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_120),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_92),
.C(n_74),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_115),
.B1(n_105),
.B2(n_107),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_113),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_88),
.Y(n_128)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_132),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_74),
.C(n_86),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_65),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_153),
.B1(n_130),
.B2(n_133),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_131),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_142),
.B(n_144),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_125),
.C(n_126),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_129),
.B(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_147),
.Y(n_174)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_108),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_111),
.B1(n_95),
.B2(n_41),
.Y(n_152)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_120),
.A2(n_111),
.B(n_47),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_137),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_23),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_139),
.B1(n_153),
.B2(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_151),
.C(n_119),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_172),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_127),
.B1(n_135),
.B2(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_137),
.B(n_122),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_15),
.B(n_23),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_134),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_70),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_22),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_14),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_194),
.B1(n_173),
.B2(n_175),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_143),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_SL g202 ( 
.A(n_183),
.B(n_188),
.C(n_190),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_169),
.A2(n_156),
.B1(n_147),
.B2(n_117),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_167),
.B1(n_172),
.B2(n_165),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_187),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_23),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_20),
.B(n_21),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_46),
.B1(n_53),
.B2(n_41),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_164),
.C(n_163),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_53),
.C(n_62),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_178),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_205),
.B(n_207),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_75),
.B1(n_66),
.B2(n_28),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_206),
.B1(n_14),
.B2(n_1),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_165),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_177),
.B1(n_171),
.B2(n_42),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_208),
.A2(n_171),
.B(n_181),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_182),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_217),
.C(n_203),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_187),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_14),
.Y(n_229)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_SL g213 ( 
.A(n_202),
.B(n_188),
.C(n_186),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_219),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_15),
.C(n_82),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_15),
.B(n_64),
.C(n_82),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_226),
.C(n_3),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_195),
.B1(n_204),
.B2(n_203),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_1),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_229),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_209),
.A3(n_218),
.B1(n_213),
.B2(n_217),
.C1(n_215),
.C2(n_216),
.Y(n_231)
);

OAI21x1_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_5),
.B(n_6),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_13),
.Y(n_232)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_5),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_3),
.B(n_4),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_4),
.Y(n_238)
);

OAI31xp33_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_228),
.A3(n_221),
.B(n_6),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_237),
.A2(n_5),
.B(n_9),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_241),
.Y(n_242)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_230),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_12),
.C(n_14),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_240),
.B(n_238),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_245),
.A2(n_246),
.B(n_242),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_12),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_12),
.Y(n_249)
);


endmodule