module real_aes_14325_n_14 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_14);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_14;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_34;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_35;
wire n_15;
wire n_27;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_0), .Y(n_26) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_1), .B(n_7), .C(n_21), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_2), .Y(n_23) );
NOR2xp33_ASAP7_75t_R g25 ( .A(n_3), .B(n_12), .Y(n_25) );
NOR2xp33_ASAP7_75t_R g28 ( .A(n_3), .B(n_29), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_3), .Y(n_35) );
NAND2xp33_ASAP7_75t_R g37 ( .A(n_3), .B(n_12), .Y(n_37) );
NAND5xp2_ASAP7_75t_SL g17 ( .A(n_4), .B(n_5), .C(n_18), .D(n_23), .E(n_24), .Y(n_17) );
AOI22xp33_ASAP7_75t_R g31 ( .A1(n_6), .A2(n_11), .B1(n_32), .B2(n_36), .Y(n_31) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_8), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_9), .Y(n_24) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_10), .Y(n_30) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_12), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g34 ( .A(n_12), .B(n_35), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_13), .Y(n_21) );
OAI221xp5_ASAP7_75t_R g14 ( .A1(n_15), .A2(n_26), .B1(n_27), .B2(n_30), .C(n_31), .Y(n_14) );
NAND2xp33_ASAP7_75t_R g15 ( .A(n_16), .B(n_25), .Y(n_15) );
NAND2xp33_ASAP7_75t_R g27 ( .A(n_16), .B(n_28), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_17), .Y(n_16) );
NOR2xp33_ASAP7_75t_R g32 ( .A(n_17), .B(n_33), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g36 ( .A(n_17), .B(n_37), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
NAND2xp33_ASAP7_75t_R g19 ( .A(n_20), .B(n_22), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_34), .Y(n_33) );
endmodule