module fake_jpeg_9726_n_19 (n_3, n_2, n_1, n_0, n_4, n_19);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_19;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_18;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g5 ( 
.A(n_1),
.B(n_3),
.Y(n_5)
);

INVx4_ASAP7_75t_SL g6 ( 
.A(n_0),
.Y(n_6)
);

MAJIxp5_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_0),
.C(n_2),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_2),
.B(n_1),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_4),
.Y(n_9)
);

AO21x1_ASAP7_75t_SL g10 ( 
.A1(n_6),
.A2(n_4),
.B(n_1),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_10),
.A2(n_8),
.B(n_5),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g11 ( 
.A1(n_9),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_11)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_12),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_3),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_14),
.A2(n_10),
.B1(n_6),
.B2(n_3),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_12),
.C(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_16),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_17),
.A2(n_15),
.B(n_0),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_17),
.B(n_2),
.Y(n_19)
);


endmodule