module fake_jpeg_30341_n_63 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_4),
.B(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_8),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_3),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_25),
.B1(n_4),
.B2(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_0),
.CI(n_2),
.CON(n_32),
.SN(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_23),
.B1(n_26),
.B2(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_40),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_23),
.B1(n_13),
.B2(n_22),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_3),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_6),
.B(n_7),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_10),
.C(n_14),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_21),
.C(n_6),
.Y(n_50)
);

NOR3xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_37),
.C(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_49),
.B(n_7),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_55),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_51),
.A2(n_54),
.B(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_54),
.Y(n_59)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_54),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

OAI221xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_56),
.B1(n_61),
.B2(n_55),
.C(n_59),
.Y(n_63)
);


endmodule