module fake_jpeg_15409_n_293 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_40),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_61),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_31),
.B1(n_32),
.B2(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_19),
.B1(n_30),
.B2(n_29),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_37),
.B1(n_19),
.B2(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_38),
.B1(n_33),
.B2(n_30),
.Y(n_84)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_34),
.B(n_28),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_28),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_78),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_37),
.CI(n_33),
.CON(n_77),
.SN(n_77)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_55),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_17),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_49),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_39),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_33),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_39),
.C(n_20),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_96),
.C(n_109),
.Y(n_138)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_71),
.Y(n_117)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_104),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

FAx1_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_50),
.CI(n_39),
.CON(n_103),
.SN(n_103)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_76),
.B(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_109),
.Y(n_114)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_112),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_27),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_68),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_50),
.B1(n_58),
.B2(n_82),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_122),
.B(n_130),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_87),
.B1(n_71),
.B2(n_79),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_106),
.B1(n_107),
.B2(n_100),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_133),
.B1(n_135),
.B2(n_137),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_69),
.Y(n_160)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_93),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_76),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_131),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_20),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_138),
.C(n_139),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_73),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_104),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_88),
.A2(n_63),
.B1(n_75),
.B2(n_46),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_0),
.B(n_85),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_16),
.B(n_21),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_63),
.B1(n_46),
.B2(n_85),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_90),
.A2(n_23),
.B1(n_22),
.B2(n_29),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_69),
.C(n_20),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_136),
.A2(n_113),
.B1(n_94),
.B2(n_105),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_153),
.C(n_160),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_101),
.B1(n_97),
.B2(n_108),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_146),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_147),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_148),
.B(n_154),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_165),
.Y(n_178)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_23),
.B1(n_22),
.B2(n_29),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_124),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_99),
.B1(n_98),
.B2(n_23),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_22),
.B1(n_21),
.B2(n_26),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_138),
.B1(n_135),
.B2(n_131),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_18),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_25),
.C(n_26),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_25),
.C(n_27),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_137),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_168),
.B(n_16),
.Y(n_182)
);

XOR2x1_ASAP7_75t_SL g168 ( 
.A(n_120),
.B(n_127),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_119),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_192),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_116),
.B1(n_118),
.B2(n_139),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_182),
.B1(n_185),
.B2(n_194),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_8),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_155),
.B(n_168),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_133),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_25),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_170),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_16),
.B(n_0),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_195),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_158),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_199),
.C(n_201),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_159),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_163),
.B1(n_159),
.B2(n_169),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_200),
.A2(n_205),
.B1(n_215),
.B2(n_218),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_161),
.C(n_183),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_166),
.C(n_167),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_214),
.C(n_217),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_157),
.B1(n_165),
.B2(n_25),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_195),
.B1(n_189),
.B2(n_171),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_177),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_180),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_170),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_181),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_191),
.C(n_174),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_217),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_228),
.C(n_230),
.Y(n_248)
);

INVxp33_ASAP7_75t_SL g220 ( 
.A(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_173),
.B(n_182),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_227),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_191),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_234),
.B1(n_208),
.B2(n_200),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_190),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_233),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_172),
.B1(n_176),
.B2(n_194),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_172),
.C(n_5),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_215),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_204),
.B(n_4),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_240),
.B(n_244),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_242),
.B(n_243),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_213),
.B1(n_203),
.B2(n_196),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_232),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_224),
.C(n_232),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_205),
.B1(n_6),
.B2(n_7),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_7),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_4),
.C(n_6),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_228),
.C(n_221),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_4),
.B(n_7),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_224),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_258),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_249),
.C(n_239),
.Y(n_269)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_235),
.C(n_8),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_256),
.B(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_242),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_242),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_10),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_252),
.C(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_237),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_262),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_274),
.B(n_271),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_238),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_279),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_269),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_263),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_285),
.C(n_278),
.Y(n_287)
);

O2A1O1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_287),
.A2(n_288),
.B(n_11),
.C(n_12),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_276),
.C(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

AO221x1_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_286),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_12),
.C(n_13),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_14),
.Y(n_293)
);


endmodule