module fake_jpeg_20042_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_45),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_43),
.Y(n_58)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_0),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_18),
.Y(n_89)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_22),
.B1(n_19),
.B2(n_32),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_23),
.B1(n_30),
.B2(n_32),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_29),
.B1(n_19),
.B2(n_32),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_39),
.B1(n_35),
.B2(n_29),
.Y(n_93)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_16),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_33),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_35),
.Y(n_94)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g105 ( 
.A(n_68),
.Y(n_105)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_73),
.Y(n_114)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_36),
.B1(n_37),
.B2(n_45),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_99),
.B1(n_39),
.B2(n_58),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_89),
.Y(n_122)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_36),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_98),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_25),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_18),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_121)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_50),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_27),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_54),
.A2(n_37),
.B1(n_39),
.B2(n_35),
.Y(n_99)
);

AO22x1_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_41),
.B1(n_38),
.B2(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_107),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_102),
.A2(n_124),
.B1(n_91),
.B2(n_66),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_42),
.C(n_38),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_20),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_43),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_59),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_29),
.B1(n_23),
.B2(n_34),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_95),
.B1(n_79),
.B2(n_65),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_72),
.B(n_40),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_59),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_41),
.B1(n_48),
.B2(n_52),
.Y(n_124)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_137),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_27),
.B1(n_34),
.B2(n_30),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_132),
.B(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_34),
.B(n_30),
.C(n_23),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_134),
.A2(n_43),
.B(n_24),
.C(n_17),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_40),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_80),
.Y(n_163)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_138),
.B(n_141),
.Y(n_187)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_145),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_65),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_154),
.B1(n_125),
.B2(n_119),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_31),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_146),
.B(n_148),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_121),
.B(n_113),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_31),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_20),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_20),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_79),
.B1(n_66),
.B2(n_41),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_102),
.B1(n_124),
.B2(n_112),
.Y(n_162)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_41),
.B1(n_78),
.B2(n_71),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_166),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_162),
.A2(n_176),
.B1(n_24),
.B2(n_1),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_163),
.B(n_171),
.Y(n_223)
);

XOR2x2_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_107),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_100),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_193),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_134),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_100),
.B1(n_122),
.B2(n_112),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_128),
.B1(n_123),
.B2(n_106),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_180),
.A2(n_183),
.B1(n_137),
.B2(n_145),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_135),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_185),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_126),
.B1(n_115),
.B2(n_127),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_28),
.Y(n_214)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_147),
.A2(n_103),
.B(n_0),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_131),
.A2(n_43),
.B(n_31),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_43),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_156),
.B(n_139),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_194),
.A2(n_202),
.B(n_191),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_159),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_198),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_155),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_199),
.B(n_203),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_206),
.B1(n_209),
.B2(n_188),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_130),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_165),
.B(n_103),
.Y(n_203)
);

AND2x6_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_144),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_160),
.A2(n_69),
.B1(n_90),
.B2(n_41),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_171),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_210),
.B(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_28),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_28),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_172),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_177),
.A2(n_64),
.B1(n_42),
.B2(n_26),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

AOI32xp33_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_26),
.A3(n_42),
.B1(n_24),
.B2(n_64),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_217),
.Y(n_238)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_9),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_179),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_192),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_235),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_187),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_194),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_198),
.C(n_204),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_230),
.C(n_239),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_183),
.C(n_178),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_202),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_26),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_201),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_175),
.C(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_223),
.C(n_200),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_248),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_244),
.A2(n_213),
.B1(n_222),
.B2(n_181),
.Y(n_252)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_209),
.B1(n_222),
.B2(n_195),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_243),
.B1(n_239),
.B2(n_240),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_250),
.B(n_42),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_257),
.B1(n_264),
.B2(n_266),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_256),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_236),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_219),
.B1(n_217),
.B2(n_189),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_219),
.CI(n_185),
.CON(n_258),
.SN(n_258)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_265),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_173),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_227),
.A2(n_174),
.B1(n_184),
.B2(n_164),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_246),
.B(n_174),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_233),
.A2(n_172),
.B1(n_24),
.B2(n_0),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_248),
.B1(n_238),
.B2(n_226),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_280),
.B1(n_1),
.B2(n_4),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_279),
.B1(n_253),
.B2(n_266),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_263),
.A2(n_226),
.B(n_237),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_281),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_255),
.B1(n_242),
.B2(n_234),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_237),
.B1(n_245),
.B2(n_230),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_64),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_42),
.C(n_2),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_286),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_269),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_42),
.C(n_2),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_291),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_264),
.C(n_250),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_290),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_283),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_258),
.C(n_257),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_295),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_258),
.C(n_3),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_273),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_1),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_299),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_280),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_270),
.B1(n_285),
.B2(n_7),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_270),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_306),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_276),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_288),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_286),
.C(n_6),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_5),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_296),
.B(n_290),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_303),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_292),
.Y(n_314)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_318),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_302),
.A2(n_301),
.B(n_7),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_310),
.B(n_305),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_5),
.C(n_7),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_320),
.B(n_312),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_8),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_322),
.B(n_316),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_320),
.C(n_10),
.Y(n_327)
);

OAI211xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_327),
.B(n_325),
.C(n_324),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_323),
.C(n_10),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_9),
.B(n_11),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_13),
.C(n_14),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_13),
.C(n_14),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_14),
.B1(n_15),
.B2(n_325),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_15),
.Y(n_334)
);


endmodule