module fake_jpeg_11428_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_62),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_0),
.B(n_1),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_61),
.Y(n_74)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_58),
.B1(n_57),
.B2(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_SL g67 ( 
.A(n_53),
.Y(n_67)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_58),
.B(n_57),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_50),
.C(n_3),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_51),
.B1(n_45),
.B2(n_52),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_45),
.B1(n_52),
.B2(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_80),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_55),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_82),
.B1(n_81),
.B2(n_79),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_93),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_88),
.B1(n_94),
.B2(n_24),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_50),
.B1(n_49),
.B2(n_48),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_47),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_19),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_17),
.B1(n_35),
.B2(n_34),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g109 ( 
.A(n_98),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_15),
.B(n_16),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_20),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_113),
.C(n_37),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_4),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_111),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_5),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_112),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_7),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_7),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_8),
.C(n_9),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_9),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_25),
.B1(n_33),
.B2(n_31),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_126),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_21),
.B1(n_22),
.B2(n_26),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_27),
.B(n_28),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_127),
.A2(n_110),
.B(n_107),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_130),
.A2(n_127),
.B1(n_123),
.B2(n_117),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_106),
.C(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_136),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_125),
.B(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_135),
.Y(n_139)
);

OAI31xp33_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_137),
.A3(n_122),
.B(n_121),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_131),
.Y(n_141)
);

OAI321xp33_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_132),
.A3(n_103),
.B1(n_120),
.B2(n_119),
.C(n_115),
.Y(n_142)
);

OAI31xp33_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_118),
.A3(n_116),
.B(n_128),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_106),
.Y(n_144)
);


endmodule