module fake_netlist_1_8798_n_14 (n_1, n_2, n_0, n_14);
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
NAND2xp5_ASAP7_75t_L g4 ( .A(n_2), .B(n_1), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
AOI22xp5_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_6) );
AO31x2_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_1), .A3(n_2), .B(n_0), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
AND2x4_ASAP7_75t_L g9 ( .A(n_6), .B(n_3), .Y(n_9) );
AO22x1_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_5), .B1(n_7), .B2(n_2), .Y(n_10) );
AOI21xp33_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_5), .B(n_2), .Y(n_11) );
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_9), .B1(n_8), .B2(n_0), .Y(n_12) );
AOI221xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_0), .B1(n_9), .B2(n_11), .C(n_10), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
endmodule