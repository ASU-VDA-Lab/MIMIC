module real_aes_670_n_367 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_367);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_367;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_963;
wire n_865;
wire n_537;
wire n_884;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_892;
wire n_994;
wire n_372;
wire n_528;
wire n_495;
wire n_578;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_755;
wire n_409;
wire n_860;
wire n_781;
wire n_909;
wire n_996;
wire n_523;
wire n_748;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_973;
wire n_960;
wire n_504;
wire n_671;
wire n_725;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_970;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_769;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_733;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_869;
wire n_613;
wire n_387;
wire n_957;
wire n_995;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_1003;
wire n_533;
wire n_1000;
wire n_727;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_691;
wire n_765;
wire n_481;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_0), .A2(n_350), .B1(n_482), .B2(n_483), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_1), .A2(n_80), .B1(n_448), .B2(n_452), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_2), .A2(n_258), .B1(n_660), .B2(n_661), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g985 ( .A1(n_3), .A2(n_103), .B1(n_413), .B2(n_417), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_4), .A2(n_168), .B1(n_660), .B2(n_777), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_5), .A2(n_261), .B1(n_555), .B2(n_558), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_6), .A2(n_328), .B1(n_438), .B2(n_494), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_7), .A2(n_35), .B1(n_430), .B2(n_828), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_8), .A2(n_26), .B1(n_408), .B2(n_536), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_9), .A2(n_329), .B1(n_434), .B2(n_437), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_10), .A2(n_83), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_11), .A2(n_65), .B1(n_488), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_12), .A2(n_363), .B1(n_475), .B2(n_609), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_13), .A2(n_202), .B1(n_400), .B2(n_407), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_14), .A2(n_143), .B1(n_428), .B2(n_526), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_15), .A2(n_43), .B1(n_444), .B2(n_774), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_16), .A2(n_178), .B1(n_437), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_17), .A2(n_121), .B1(n_483), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_18), .A2(n_226), .B1(n_479), .B2(n_480), .Y(n_568) );
AO222x2_ASAP7_75t_L g564 ( .A1(n_19), .A2(n_193), .B1(n_239), .B2(n_472), .C1(n_475), .C2(n_476), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_20), .A2(n_147), .B1(n_424), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_21), .A2(n_22), .B1(n_549), .B2(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_23), .A2(n_349), .B1(n_491), .B2(n_733), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_24), .A2(n_180), .B1(n_494), .B2(n_495), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_25), .A2(n_216), .B1(n_658), .B2(n_690), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_27), .A2(n_232), .B1(n_555), .B2(n_556), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_28), .A2(n_172), .B1(n_519), .B2(n_947), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_29), .A2(n_122), .B1(n_512), .B2(n_877), .Y(n_951) );
AO22x1_ASAP7_75t_L g764 ( .A1(n_30), .A2(n_221), .B1(n_700), .B2(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_31), .A2(n_123), .B1(n_511), .B2(n_512), .Y(n_510) );
INVx1_ASAP7_75t_SL g388 ( .A(n_32), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g966 ( .A(n_32), .B(n_40), .Y(n_966) );
INVx1_ASAP7_75t_L g925 ( .A(n_33), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_34), .A2(n_215), .B1(n_656), .B2(n_658), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g902 ( .A1(n_36), .A2(n_313), .B1(n_833), .B2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_37), .A2(n_186), .B1(n_482), .B2(n_483), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_38), .A2(n_77), .B1(n_479), .B2(n_480), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_39), .B(n_472), .Y(n_546) );
AO22x2_ASAP7_75t_L g390 ( .A1(n_40), .A2(n_338), .B1(n_387), .B2(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_41), .B(n_472), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_42), .A2(n_292), .B1(n_690), .B2(n_691), .Y(n_689) );
XOR2xp5_ASAP7_75t_L g701 ( .A(n_44), .B(n_702), .Y(n_701) );
XOR2xp5_ASAP7_75t_L g736 ( .A(n_44), .B(n_737), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_45), .A2(n_82), .B1(n_690), .B2(n_845), .Y(n_948) );
INVx1_ASAP7_75t_L g389 ( .A(n_46), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_47), .A2(n_81), .B1(n_428), .B2(n_526), .Y(n_712) );
XNOR2xp5_ASAP7_75t_L g856 ( .A(n_48), .B(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_49), .A2(n_96), .B1(n_498), .B2(n_560), .Y(n_758) );
AOI22xp33_ASAP7_75t_SL g792 ( .A1(n_50), .A2(n_315), .B1(n_624), .B2(n_769), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_51), .A2(n_294), .B1(n_656), .B2(n_658), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_52), .A2(n_347), .B1(n_909), .B2(n_912), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_53), .A2(n_278), .B1(n_437), .B2(n_682), .Y(n_937) );
AO22x1_ASAP7_75t_L g766 ( .A1(n_54), .A2(n_359), .B1(n_698), .B2(n_706), .Y(n_766) );
AOI222xp33_ASAP7_75t_L g979 ( .A1(n_55), .A2(n_980), .B1(n_994), .B2(n_996), .C1(n_998), .C2(n_1001), .Y(n_979) );
XNOR2x1_ASAP7_75t_L g981 ( .A(n_55), .B(n_982), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_56), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_57), .A2(n_224), .B1(n_488), .B2(n_553), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_58), .A2(n_166), .B1(n_479), .B2(n_607), .Y(n_606) );
AO22x2_ASAP7_75t_L g397 ( .A1(n_59), .A2(n_175), .B1(n_387), .B2(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_60), .A2(n_353), .B1(n_418), .B2(n_892), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_61), .A2(n_334), .B1(n_444), .B2(n_639), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_62), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_63), .A2(n_129), .B1(n_487), .B2(n_488), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_64), .A2(n_146), .B1(n_917), .B2(n_918), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_66), .A2(n_209), .B1(n_434), .B2(n_661), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_67), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_68), .A2(n_138), .B1(n_685), .B2(n_686), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_69), .A2(n_317), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_70), .A2(n_207), .B1(n_414), .B2(n_532), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_71), .A2(n_376), .B1(n_377), .B2(n_464), .Y(n_375) );
INVx1_ASAP7_75t_L g464 ( .A(n_71), .Y(n_464) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_72), .A2(n_88), .B1(n_183), .B2(n_472), .C1(n_482), .C2(n_567), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_73), .A2(n_271), .B1(n_497), .B2(n_498), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_74), .A2(n_241), .B1(n_518), .B2(n_880), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_75), .A2(n_185), .B1(n_497), .B2(n_558), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_76), .A2(n_101), .B1(n_448), .B2(n_452), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_78), .A2(n_364), .B1(n_482), .B2(n_567), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_79), .A2(n_346), .B1(n_482), .B2(n_567), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_84), .B(n_381), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_85), .A2(n_164), .B1(n_424), .B2(n_930), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_86), .A2(n_131), .B1(n_487), .B2(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_87), .A2(n_191), .B1(n_682), .B2(n_777), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_89), .A2(n_114), .B1(n_488), .B2(n_553), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_90), .A2(n_251), .B1(n_706), .B2(n_708), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_91), .A2(n_196), .B1(n_498), .B2(n_560), .Y(n_559) );
OA22x2_ASAP7_75t_L g600 ( .A1(n_92), .A2(n_601), .B1(n_602), .B2(n_603), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_92), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_93), .A2(n_100), .B1(n_558), .B2(n_560), .Y(n_614) );
XNOR2xp5_ASAP7_75t_L g996 ( .A(n_94), .B(n_997), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_95), .A2(n_285), .B1(n_497), .B2(n_558), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_97), .A2(n_284), .B1(n_413), .B2(n_417), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_98), .A2(n_127), .B1(n_490), .B2(n_491), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_99), .A2(n_341), .B1(n_488), .B2(n_553), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_102), .A2(n_214), .B1(n_497), .B2(n_498), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_104), .A2(n_358), .B1(n_497), .B2(n_498), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_105), .A2(n_244), .B1(n_627), .B2(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_106), .A2(n_323), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_107), .A2(n_243), .B1(n_779), .B2(n_798), .Y(n_797) );
XNOR2xp5_ASAP7_75t_L g561 ( .A(n_108), .B(n_562), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_109), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_110), .A2(n_342), .B1(n_463), .B2(n_497), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_111), .A2(n_201), .B1(n_475), .B2(n_476), .Y(n_747) );
AO22x2_ASAP7_75t_L g394 ( .A1(n_112), .A2(n_275), .B1(n_387), .B2(n_395), .Y(n_394) );
AOI222xp33_ASAP7_75t_SL g989 ( .A1(n_113), .A2(n_262), .B1(n_333), .B2(n_527), .C1(n_590), .C2(n_990), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_115), .A2(n_135), .B1(n_697), .B2(n_698), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_116), .Y(n_861) );
XOR2x2_ASAP7_75t_L g883 ( .A(n_117), .B(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_118), .A2(n_276), .B1(n_686), .B2(n_733), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_119), .A2(n_356), .B1(n_685), .B2(n_686), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_120), .A2(n_316), .B1(n_514), .B2(n_915), .Y(n_914) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_124), .A2(n_157), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_125), .A2(n_194), .B1(n_448), .B2(n_452), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_126), .A2(n_197), .B1(n_625), .B2(n_665), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_128), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_130), .A2(n_161), .B1(n_480), .B2(n_536), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_132), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_133), .A2(n_167), .B1(n_479), .B2(n_480), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_134), .A2(n_293), .B1(n_556), .B2(n_576), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_136), .A2(n_223), .B1(n_833), .B2(n_903), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_137), .A2(n_326), .B1(n_488), .B2(n_553), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_139), .A2(n_250), .B1(n_424), .B2(n_428), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_140), .A2(n_159), .B1(n_774), .B2(n_775), .Y(n_773) );
AOI222xp33_ASAP7_75t_L g952 ( .A1(n_141), .A2(n_163), .B1(n_210), .B2(n_381), .C1(n_697), .C2(n_698), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g575 ( .A1(n_142), .A2(n_289), .B1(n_556), .B2(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_144), .A2(n_298), .B1(n_625), .B2(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_145), .B(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_148), .A2(n_327), .B1(n_488), .B2(n_553), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_149), .A2(n_257), .B1(n_475), .B2(n_609), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_150), .B(n_621), .Y(n_620) );
AO21x2_ASAP7_75t_L g824 ( .A1(n_151), .A2(n_825), .B(n_846), .Y(n_824) );
INVx1_ASAP7_75t_L g848 ( .A(n_151), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_152), .A2(n_234), .B1(n_518), .B2(n_519), .Y(n_517) );
AO22x2_ASAP7_75t_L g810 ( .A1(n_153), .A2(n_811), .B1(n_822), .B2(n_823), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_153), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_154), .A2(n_309), .B1(n_448), .B2(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_155), .B(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_156), .A2(n_227), .B1(n_463), .B2(n_639), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_158), .A2(n_176), .B1(n_448), .B2(n_452), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_160), .A2(n_354), .B1(n_682), .B2(n_683), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_162), .A2(n_331), .B1(n_534), .B2(n_538), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_165), .A2(n_291), .B1(n_475), .B2(n_476), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_169), .A2(n_264), .B1(n_549), .B2(n_567), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_170), .A2(n_310), .B1(n_414), .B2(n_418), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_171), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_173), .A2(n_188), .B1(n_401), .B2(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_174), .A2(n_268), .B1(n_434), .B2(n_718), .Y(n_992) );
INVx1_ASAP7_75t_L g965 ( .A(n_175), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_177), .A2(n_272), .B1(n_407), .B2(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_179), .A2(n_319), .B1(n_514), .B2(n_516), .Y(n_513) );
AO222x2_ASAP7_75t_SL g827 ( .A1(n_181), .A2(n_269), .B1(n_325), .B2(n_590), .C1(n_828), .C2(n_829), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_182), .A2(n_286), .B1(n_555), .B2(n_556), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_184), .A2(n_365), .B1(n_497), .B2(n_498), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_187), .A2(n_240), .B1(n_490), .B2(n_498), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_189), .A2(n_235), .B1(n_479), .B2(n_480), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_190), .A2(n_307), .B1(n_635), .B2(n_636), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g876 ( .A1(n_192), .A2(n_282), .B1(n_877), .B2(n_878), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_195), .A2(n_273), .B1(n_529), .B2(n_531), .Y(n_905) );
XNOR2x2_ASAP7_75t_L g761 ( .A(n_198), .B(n_762), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_199), .A2(n_274), .B1(n_495), .B2(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_200), .B(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_203), .B(n_698), .Y(n_862) );
NAND2xp5_ASAP7_75t_SL g906 ( .A(n_204), .B(n_522), .Y(n_906) );
XNOR2x1_ASAP7_75t_L g647 ( .A(n_205), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g975 ( .A(n_206), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_208), .A2(n_295), .B1(n_627), .B2(n_628), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_211), .A2(n_366), .B1(n_494), .B2(n_718), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_212), .A2(n_941), .B1(n_953), .B2(n_954), .Y(n_940) );
INVx1_ASAP7_75t_L g954 ( .A(n_212), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_213), .B(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g932 ( .A1(n_217), .A2(n_344), .B1(n_408), .B2(n_700), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_218), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_219), .A2(n_230), .B1(n_529), .B2(n_531), .Y(n_528) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_220), .A2(n_321), .B1(n_488), .B2(n_572), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_222), .A2(n_324), .B1(n_636), .B2(n_909), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_225), .B(n_771), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_228), .A2(n_280), .B1(n_624), .B2(n_625), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_229), .A2(n_302), .B1(n_531), .B2(n_672), .Y(n_671) );
XNOR2x1_ASAP7_75t_L g543 ( .A(n_231), .B(n_544), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_233), .A2(n_300), .B1(n_538), .B2(n_627), .Y(n_943) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_236), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_237), .A2(n_303), .B1(n_558), .B2(n_560), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_238), .A2(n_357), .B1(n_658), .B2(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_242), .A2(n_301), .B1(n_401), .B2(n_670), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_245), .Y(n_837) );
XOR2x2_ASAP7_75t_L g899 ( .A(n_246), .B(n_900), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_247), .A2(n_360), .B1(n_414), .B2(n_532), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_248), .A2(n_351), .B1(n_635), .B2(n_654), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_249), .Y(n_860) );
INVx1_ASAP7_75t_L g978 ( .A(n_252), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_253), .A2(n_320), .B1(n_441), .B2(n_444), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g873 ( .A1(n_254), .A2(n_340), .B1(n_512), .B2(n_660), .Y(n_873) );
XNOR2x1_ASAP7_75t_L g617 ( .A(n_255), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g499 ( .A(n_256), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_259), .A2(n_263), .B1(n_497), .B2(n_498), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_260), .A2(n_283), .B1(n_457), .B2(n_461), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_265), .A2(n_306), .B1(n_556), .B2(n_576), .Y(n_755) );
OA22x2_ASAP7_75t_L g578 ( .A1(n_266), .A2(n_579), .B1(n_580), .B2(n_594), .Y(n_578) );
INVx1_ASAP7_75t_L g594 ( .A(n_266), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_267), .B(n_667), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_270), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_275), .B(n_964), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_277), .A2(n_332), .B1(n_670), .B2(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_279), .A2(n_336), .B1(n_462), .B2(n_633), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_281), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_287), .A2(n_305), .B1(n_529), .B2(n_531), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_288), .A2(n_312), .B1(n_441), .B2(n_556), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_290), .A2(n_322), .B1(n_530), .B2(n_698), .Y(n_790) );
INVx3_ASAP7_75t_L g387 ( .A(n_296), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_297), .A2(n_311), .B1(n_518), .B2(n_654), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_299), .Y(n_840) );
OA22x2_ASAP7_75t_L g504 ( .A1(n_304), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_304), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_308), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_314), .B(n_590), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_318), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_330), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_335), .A2(n_343), .B1(n_479), .B2(n_607), .Y(n_750) );
INVx1_ASAP7_75t_L g759 ( .A(n_337), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_339), .B(n_771), .Y(n_896) );
INVx1_ASAP7_75t_L g960 ( .A(n_345), .Y(n_960) );
AND2x4_ASAP7_75t_L g977 ( .A(n_345), .B(n_961), .Y(n_977) );
AO21x1_ASAP7_75t_L g1002 ( .A1(n_345), .A2(n_973), .B(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g961 ( .A(n_348), .Y(n_961) );
AND2x2_ASAP7_75t_R g1000 ( .A(n_348), .B(n_960), .Y(n_1000) );
INVxp67_ASAP7_75t_L g974 ( .A(n_352), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_355), .B(n_771), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_361), .Y(n_864) );
XNOR2xp5_ASAP7_75t_L g678 ( .A(n_362), .B(n_679), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_967), .B(n_970), .Y(n_367) );
AOI21xp33_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_642), .B(n_957), .Y(n_368) );
INVx1_ASAP7_75t_L g968 ( .A(n_369), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_615), .B1(n_640), .B2(n_641), .Y(n_369) );
XOR2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_501), .Y(n_370) );
XNOR2xp5_ASAP7_75t_L g640 ( .A(n_371), .B(n_501), .Y(n_640) );
BUFx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI22x1_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_465), .B2(n_500), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx2_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_432), .Y(n_377) );
NAND4xp25_ASAP7_75t_SL g378 ( .A(n_379), .B(n_399), .C(n_412), .D(n_423), .Y(n_378) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx3_ASAP7_75t_SL g524 ( .A(n_382), .Y(n_524) );
INVx3_ASAP7_75t_L g590 ( .A(n_382), .Y(n_590) );
INVx4_ASAP7_75t_SL g621 ( .A(n_382), .Y(n_621) );
BUFx2_ASAP7_75t_L g668 ( .A(n_382), .Y(n_668) );
INVx4_ASAP7_75t_SL g771 ( .A(n_382), .Y(n_771) );
INVx6_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_392), .Y(n_383) );
AND2x4_ASAP7_75t_L g409 ( .A(n_384), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g430 ( .A(n_384), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g472 ( .A(n_384), .B(n_392), .Y(n_472) );
AND2x2_ASAP7_75t_L g480 ( .A(n_384), .B(n_410), .Y(n_480) );
AND2x2_ASAP7_75t_L g483 ( .A(n_384), .B(n_431), .Y(n_483) );
AND2x2_ASAP7_75t_L g567 ( .A(n_384), .B(n_431), .Y(n_567) );
AND2x2_ASAP7_75t_L g607 ( .A(n_384), .B(n_410), .Y(n_607) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_390), .Y(n_384) );
AND2x2_ASAP7_75t_L g405 ( .A(n_385), .B(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_385), .Y(n_422) );
INVx2_ASAP7_75t_L g427 ( .A(n_385), .Y(n_427) );
OAI22x1_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_388), .B2(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g391 ( .A(n_387), .Y(n_391) );
INVx2_ASAP7_75t_L g395 ( .A(n_387), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_387), .Y(n_398) );
INVx2_ASAP7_75t_L g406 ( .A(n_390), .Y(n_406) );
AND2x2_ASAP7_75t_L g426 ( .A(n_390), .B(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g455 ( .A(n_390), .Y(n_455) );
AND2x4_ASAP7_75t_L g436 ( .A(n_392), .B(n_405), .Y(n_436) );
AND2x4_ASAP7_75t_L g443 ( .A(n_392), .B(n_439), .Y(n_443) );
AND2x2_ASAP7_75t_L g460 ( .A(n_392), .B(n_426), .Y(n_460) );
AND2x6_ASAP7_75t_L g497 ( .A(n_392), .B(n_426), .Y(n_497) );
AND2x2_ASAP7_75t_L g555 ( .A(n_392), .B(n_405), .Y(n_555) );
AND2x2_ASAP7_75t_L g560 ( .A(n_392), .B(n_439), .Y(n_560) );
AND2x2_ASAP7_75t_L g576 ( .A(n_392), .B(n_405), .Y(n_576) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_396), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g404 ( .A(n_394), .Y(n_404) );
AND2x4_ASAP7_75t_L g416 ( .A(n_394), .B(n_396), .Y(n_416) );
AND2x2_ASAP7_75t_L g421 ( .A(n_394), .B(n_397), .Y(n_421) );
INVxp67_ASAP7_75t_L g431 ( .A(n_396), .Y(n_431) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g403 ( .A(n_397), .B(n_404), .Y(n_403) );
BUFx6f_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g537 ( .A(n_402), .Y(n_537) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_402), .Y(n_627) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
AND2x4_ASAP7_75t_L g446 ( .A(n_403), .B(n_439), .Y(n_446) );
AND2x2_ASAP7_75t_L g451 ( .A(n_403), .B(n_426), .Y(n_451) );
AND2x4_ASAP7_75t_L g479 ( .A(n_403), .B(n_405), .Y(n_479) );
AND2x6_ASAP7_75t_L g498 ( .A(n_403), .B(n_439), .Y(n_498) );
AND2x2_ASAP7_75t_L g553 ( .A(n_403), .B(n_426), .Y(n_553) );
AND2x2_ASAP7_75t_SL g572 ( .A(n_403), .B(n_426), .Y(n_572) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_404), .Y(n_411) );
AND2x2_ASAP7_75t_L g415 ( .A(n_405), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g475 ( .A(n_405), .B(n_416), .Y(n_475) );
AND2x4_ASAP7_75t_L g439 ( .A(n_406), .B(n_427), .Y(n_439) );
BUFx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g540 ( .A(n_409), .Y(n_540) );
INVx1_ASAP7_75t_L g629 ( .A(n_409), .Y(n_629) );
BUFx4f_ASAP7_75t_L g670 ( .A(n_409), .Y(n_670) );
BUFx3_ASAP7_75t_L g794 ( .A(n_409), .Y(n_794) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g530 ( .A(n_415), .Y(n_530) );
BUFx5_ASAP7_75t_L g697 ( .A(n_415), .Y(n_697) );
INVx2_ASAP7_75t_L g707 ( .A(n_415), .Y(n_707) );
AND2x4_ASAP7_75t_L g425 ( .A(n_416), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g463 ( .A(n_416), .B(n_439), .Y(n_463) );
AND2x2_ASAP7_75t_L g482 ( .A(n_416), .B(n_426), .Y(n_482) );
AND2x2_ASAP7_75t_L g549 ( .A(n_416), .B(n_426), .Y(n_549) );
AND2x2_ASAP7_75t_L g558 ( .A(n_416), .B(n_439), .Y(n_558) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g532 ( .A(n_419), .Y(n_532) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx12f_ASAP7_75t_L g698 ( .A(n_420), .Y(n_698) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AND2x4_ASAP7_75t_L g438 ( .A(n_421), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g454 ( .A(n_421), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_SL g476 ( .A(n_421), .B(n_422), .Y(n_476) );
AND2x4_ASAP7_75t_L g488 ( .A(n_421), .B(n_455), .Y(n_488) );
AND2x4_ASAP7_75t_L g556 ( .A(n_421), .B(n_439), .Y(n_556) );
AND2x2_ASAP7_75t_SL g609 ( .A(n_421), .B(n_422), .Y(n_609) );
BUFx4f_ASAP7_75t_SL g526 ( .A(n_424), .Y(n_526) );
BUFx2_ASAP7_75t_L g828 ( .A(n_424), .Y(n_828) );
BUFx2_ASAP7_75t_L g990 ( .A(n_424), .Y(n_990) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx2_ASAP7_75t_L g624 ( .A(n_425), .Y(n_624) );
BUFx3_ASAP7_75t_L g665 ( .A(n_425), .Y(n_665) );
BUFx2_ASAP7_75t_L g695 ( .A(n_425), .Y(n_695) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g527 ( .A(n_429), .Y(n_527) );
INVx2_ASAP7_75t_SL g625 ( .A(n_429), .Y(n_625) );
INVx2_ASAP7_75t_L g769 ( .A(n_429), .Y(n_769) );
INVx2_ASAP7_75t_L g829 ( .A(n_429), .Y(n_829) );
OAI22xp33_ASAP7_75t_L g867 ( .A1(n_429), .A2(n_868), .B1(n_869), .B2(n_870), .Y(n_867) );
INVx1_ASAP7_75t_L g930 ( .A(n_429), .Y(n_930) );
INVx6_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND4xp25_ASAP7_75t_L g432 ( .A(n_433), .B(n_440), .C(n_447), .D(n_456), .Y(n_432) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g511 ( .A(n_435), .Y(n_511) );
INVx2_ASAP7_75t_L g660 ( .A(n_435), .Y(n_660) );
INVx3_ASAP7_75t_L g688 ( .A(n_435), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_435), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_714) );
INVx1_ASAP7_75t_SL g917 ( .A(n_435), .Y(n_917) );
INVx6_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx3_ASAP7_75t_L g494 ( .A(n_436), .Y(n_494) );
BUFx3_ASAP7_75t_L g633 ( .A(n_436), .Y(n_633) );
BUFx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx3_ASAP7_75t_L g495 ( .A(n_438), .Y(n_495) );
BUFx2_ASAP7_75t_SL g512 ( .A(n_438), .Y(n_512) );
INVx2_ASAP7_75t_L g662 ( .A(n_438), .Y(n_662) );
BUFx2_ASAP7_75t_SL g918 ( .A(n_438), .Y(n_918) );
INVx2_ASAP7_75t_L g515 ( .A(n_441), .Y(n_515) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_441), .Y(n_651) );
INVx4_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_SL g490 ( .A(n_442), .Y(n_490) );
INVx3_ASAP7_75t_L g639 ( .A(n_442), .Y(n_639) );
INVx2_ASAP7_75t_SL g682 ( .A(n_442), .Y(n_682) );
INVx2_ASAP7_75t_L g733 ( .A(n_442), .Y(n_733) );
INVx2_ASAP7_75t_SL g877 ( .A(n_442), .Y(n_877) );
INVx8_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g519 ( .A(n_445), .Y(n_519) );
INVx2_ASAP7_75t_SL g654 ( .A(n_445), .Y(n_654) );
INVx2_ASAP7_75t_L g686 ( .A(n_445), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_445), .A2(n_720), .B1(n_721), .B2(n_723), .Y(n_719) );
INVx2_ASAP7_75t_L g775 ( .A(n_445), .Y(n_775) );
INVx1_ASAP7_75t_SL g878 ( .A(n_445), .Y(n_878) );
INVx2_ASAP7_75t_L g912 ( .A(n_445), .Y(n_912) );
INVx8_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g657 ( .A(n_450), .Y(n_657) );
INVx1_ASAP7_75t_L g779 ( .A(n_450), .Y(n_779) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx3_ASAP7_75t_L g487 ( .A(n_451), .Y(n_487) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_451), .Y(n_690) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g658 ( .A(n_453), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_453), .A2(n_726), .B1(n_727), .B2(n_729), .Y(n_725) );
INVx2_ASAP7_75t_L g798 ( .A(n_453), .Y(n_798) );
INVx2_ASAP7_75t_L g845 ( .A(n_453), .Y(n_845) );
INVx5_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g586 ( .A(n_454), .Y(n_586) );
BUFx3_ASAP7_75t_L g691 ( .A(n_454), .Y(n_691) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_SL g518 ( .A(n_459), .Y(n_518) );
INVx3_ASAP7_75t_L g635 ( .A(n_459), .Y(n_635) );
INVx2_ASAP7_75t_L g774 ( .A(n_459), .Y(n_774) );
INVx2_ASAP7_75t_SL g947 ( .A(n_459), .Y(n_947) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g685 ( .A(n_460), .Y(n_685) );
BUFx2_ASAP7_75t_L g911 ( .A(n_460), .Y(n_911) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g881 ( .A(n_462), .Y(n_881) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_463), .Y(n_491) );
INVx2_ASAP7_75t_L g637 ( .A(n_463), .Y(n_637) );
BUFx3_ASAP7_75t_L g777 ( .A(n_463), .Y(n_777) );
INVx1_ASAP7_75t_SL g500 ( .A(n_465), .Y(n_500) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
XOR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_499), .Y(n_467) );
NAND2x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_484), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_477), .Y(n_469) );
OAI21xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_473), .B(n_474), .Y(n_470) );
INVx2_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_481), .Y(n_477) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_492), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_489), .Y(n_485) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_491), .Y(n_516) );
INVx2_ASAP7_75t_L g735 ( .A(n_491), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .Y(n_492) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_495), .Y(n_718) );
XOR2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_598), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_541), .B2(n_597), .Y(n_502) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_520), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .C(n_513), .D(n_517), .Y(n_508) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND4xp25_ASAP7_75t_SL g520 ( .A(n_521), .B(n_525), .C(n_528), .D(n_533), .Y(n_520) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OAI21xp33_ASAP7_75t_SL g788 ( .A1(n_523), .A2(n_789), .B(n_790), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g859 ( .A1(n_523), .A2(n_673), .B1(n_860), .B2(n_861), .C(n_862), .Y(n_859) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g869 ( .A(n_526), .Y(n_869) );
BUFx6f_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g673 ( .A(n_530), .Y(n_673) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
INVx4_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g700 ( .A(n_537), .Y(n_700) );
INVx1_ASAP7_75t_L g834 ( .A(n_537), .Y(n_834) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_539), .A2(n_864), .B1(n_865), .B2(n_866), .Y(n_863) );
BUFx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g765 ( .A(n_540), .Y(n_765) );
INVx1_ASAP7_75t_L g597 ( .A(n_541), .Y(n_597) );
OA22x2_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_578), .B1(n_595), .B2(n_596), .Y(n_541) );
INVx1_ASAP7_75t_L g596 ( .A(n_542), .Y(n_596) );
XOR2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_561), .Y(n_542) );
OR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_551), .Y(n_544) );
NAND4xp25_ASAP7_75t_SL g545 ( .A(n_546), .B(n_547), .C(n_548), .D(n_550), .Y(n_545) );
NAND4xp25_ASAP7_75t_SL g551 ( .A(n_552), .B(n_554), .C(n_557), .D(n_559), .Y(n_551) );
NAND2x1_ASAP7_75t_L g562 ( .A(n_563), .B(n_569), .Y(n_562) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_574), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
INVx1_ASAP7_75t_L g595 ( .A(n_578), .Y(n_595) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NOR2xp67_ASAP7_75t_L g580 ( .A(n_581), .B(n_588), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .C(n_587), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NAND4xp25_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .C(n_592), .D(n_593), .Y(n_588) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NOR2x1_ASAP7_75t_L g603 ( .A(n_604), .B(n_610), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .C(n_608), .Y(n_604) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .C(n_613), .D(n_614), .Y(n_610) );
INVx2_ASAP7_75t_L g641 ( .A(n_615), .Y(n_641) );
BUFx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g674 ( .A(n_616), .Y(n_674) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_630), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .C(n_623), .D(n_626), .Y(n_619) );
INVx2_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
NAND4xp25_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .C(n_634), .D(n_638), .Y(n_630) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g652 ( .A(n_637), .Y(n_652) );
INVx2_ASAP7_75t_L g683 ( .A(n_637), .Y(n_683) );
INVxp67_ASAP7_75t_L g969 ( .A(n_642), .Y(n_969) );
XNOR2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_851), .Y(n_642) );
XOR2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_739), .Y(n_643) );
XOR2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_675), .Y(n_644) );
XOR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_674), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NOR2x1_ASAP7_75t_L g648 ( .A(n_649), .B(n_663), .Y(n_648) );
NAND4xp25_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .C(n_655), .D(n_659), .Y(n_649) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g728 ( .A(n_657), .Y(n_728) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .C(n_669), .D(n_671), .Y(n_663) );
INVx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_701), .B1(n_736), .B2(n_738), .Y(n_676) );
INVx1_ASAP7_75t_L g738 ( .A(n_677), .Y(n_738) );
BUFx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2xp67_ASAP7_75t_L g679 ( .A(n_680), .B(n_692), .Y(n_679) );
NAND4xp25_ASAP7_75t_L g680 ( .A(n_681), .B(n_684), .C(n_687), .D(n_689), .Y(n_680) );
BUFx3_ASAP7_75t_L g722 ( .A(n_685), .Y(n_722) );
NAND4xp25_ASAP7_75t_SL g692 ( .A(n_693), .B(n_694), .C(n_696), .D(n_699), .Y(n_692) );
BUFx3_ASAP7_75t_L g708 ( .A(n_698), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_713), .C(n_724), .Y(n_702) );
AND3x1_ASAP7_75t_L g737 ( .A(n_703), .B(n_713), .C(n_724), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_710), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_705), .B(n_709), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g892 ( .A(n_707), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_719), .Y(n_713) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_730), .Y(n_724) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_734), .B2(n_735), .Y(n_730) );
OAI221xp5_ASAP7_75t_SL g836 ( .A1(n_732), .A2(n_837), .B1(n_838), .B2(n_840), .C(n_841), .Y(n_836) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g915 ( .A(n_735), .Y(n_915) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_807), .B1(n_849), .B2(n_850), .Y(n_739) );
INVx1_ASAP7_75t_SL g849 ( .A(n_740), .Y(n_849) );
AOI22x1_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_782), .B1(n_804), .B2(n_805), .Y(n_740) );
BUFx2_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g804 ( .A(n_742), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_760), .B1(n_761), .B2(n_781), .Y(n_742) );
INVx3_ASAP7_75t_SL g781 ( .A(n_743), .Y(n_781) );
OA22x2_ASAP7_75t_L g922 ( .A1(n_743), .A2(n_781), .B1(n_923), .B2(n_924), .Y(n_922) );
XOR2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_759), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_752), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_747), .B(n_748), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_756), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_772), .Y(n_762) );
NOR3xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .C(n_767), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g767 ( .A(n_768), .B(n_770), .Y(n_767) );
AND4x1_ASAP7_75t_L g772 ( .A(n_773), .B(n_776), .C(n_778), .D(n_780), .Y(n_772) );
BUFx2_ASAP7_75t_L g839 ( .A(n_777), .Y(n_839) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g806 ( .A(n_785), .Y(n_806) );
XNOR2x1_ASAP7_75t_L g785 ( .A(n_786), .B(n_803), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_795), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_791), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
BUFx6f_ASAP7_75t_SL g903 ( .A(n_794), .Y(n_903) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_800), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_799), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
INVxp67_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVxp33_ASAP7_75t_L g850 ( .A(n_808), .Y(n_850) );
XNOR2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_824), .Y(n_808) );
INVx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g823 ( .A(n_811), .Y(n_823) );
NOR2xp67_ASAP7_75t_L g811 ( .A(n_812), .B(n_817), .Y(n_811) );
NAND4xp25_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .C(n_815), .D(n_816), .Y(n_812) );
NAND4xp25_ASAP7_75t_SL g817 ( .A(n_818), .B(n_819), .C(n_820), .D(n_821), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_835), .C(n_842), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_830), .Y(n_826) );
NOR4xp25_ASAP7_75t_L g846 ( .A(n_827), .B(n_830), .C(n_836), .D(n_847), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_832), .Y(n_830) );
INVx1_ASAP7_75t_L g865 ( .A(n_833), .Y(n_865) );
BUFx3_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVxp67_ASAP7_75t_SL g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_SL g847 ( .A(n_842), .B(n_848), .Y(n_847) );
AND2x2_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
OAI22xp5_ASAP7_75t_SL g851 ( .A1(n_852), .A2(n_919), .B1(n_920), .B2(n_956), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_853), .Y(n_956) );
OA22x2_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B1(n_898), .B2(n_899), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_882), .B1(n_883), .B2(n_897), .Y(n_855) );
INVx1_ASAP7_75t_L g897 ( .A(n_856), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_871), .Y(n_857) );
NOR3xp33_ASAP7_75t_L g858 ( .A(n_859), .B(n_863), .C(n_867), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_875), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_876), .B(n_879), .Y(n_875) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
NOR3xp33_ASAP7_75t_L g884 ( .A(n_885), .B(n_890), .C(n_894), .Y(n_884) );
NAND4xp25_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .C(n_888), .D(n_889), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_893), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_895), .B(n_896), .Y(n_894) );
INVx4_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
NOR2x1_ASAP7_75t_L g900 ( .A(n_901), .B(n_907), .Y(n_900) );
NAND4xp25_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .C(n_905), .D(n_906), .Y(n_901) );
NAND4xp25_ASAP7_75t_L g907 ( .A(n_908), .B(n_913), .C(n_914), .D(n_916), .Y(n_907) );
INVx2_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
OAI22xp33_ASAP7_75t_R g920 ( .A1(n_921), .A2(n_922), .B1(n_938), .B2(n_955), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
XNOR2x2_ASAP7_75t_SL g924 ( .A(n_925), .B(n_926), .Y(n_924) );
OR2x2_ASAP7_75t_L g926 ( .A(n_927), .B(n_933), .Y(n_926) );
NAND4xp25_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .C(n_931), .D(n_932), .Y(n_927) );
NAND4xp25_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .C(n_936), .D(n_937), .Y(n_933) );
INVx1_ASAP7_75t_SL g955 ( .A(n_938), .Y(n_955) );
BUFx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_SL g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g953 ( .A(n_941), .Y(n_953) );
NAND4xp75_ASAP7_75t_L g941 ( .A(n_942), .B(n_945), .C(n_949), .D(n_952), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_943), .B(n_944), .Y(n_942) );
AND2x2_ASAP7_75t_L g945 ( .A(n_946), .B(n_948), .Y(n_945) );
AND2x2_ASAP7_75t_L g949 ( .A(n_950), .B(n_951), .Y(n_949) );
INVx4_ASAP7_75t_R g957 ( .A(n_958), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_962), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_959), .B(n_963), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_960), .B(n_961), .Y(n_959) );
INVx1_ASAP7_75t_L g1003 ( .A(n_961), .Y(n_1003) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_966), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_968), .B(n_969), .Y(n_967) );
OAI21xp5_ASAP7_75t_L g970 ( .A1(n_971), .A2(n_978), .B(n_979), .Y(n_970) );
OR2x2_ASAP7_75t_L g971 ( .A(n_972), .B(n_976), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
NOR2xp33_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .Y(n_973) );
INVxp67_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVxp67_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
INVx2_ASAP7_75t_L g997 ( .A(n_982), .Y(n_997) );
NAND4xp75_ASAP7_75t_L g982 ( .A(n_983), .B(n_986), .C(n_989), .D(n_991), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_984), .B(n_985), .Y(n_983) );
AND2x2_ASAP7_75t_L g986 ( .A(n_987), .B(n_988), .Y(n_986) );
AND2x2_ASAP7_75t_SL g991 ( .A(n_992), .B(n_993), .Y(n_991) );
CKINVDCx6p67_ASAP7_75t_R g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_SL g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_1002), .Y(n_1001) );
endmodule