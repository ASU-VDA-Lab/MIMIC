module real_jpeg_2282_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_2),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_2),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_42),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_3),
.A2(n_32),
.B1(n_40),
.B2(n_43),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_3),
.A2(n_32),
.B1(n_55),
.B2(n_56),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_3),
.B(n_40),
.C(n_52),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_3),
.B(n_51),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_3),
.B(n_27),
.C(n_37),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_3),
.B(n_70),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_3),
.B(n_21),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_22),
.C(n_24),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_3),
.B(n_35),
.Y(n_146)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_106),
.B1(n_164),
.B2(n_165),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_13),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_105),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_83),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_15),
.B(n_83),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_64),
.C(n_74),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_16),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_49),
.B2(n_63),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_33),
.B1(n_34),
.B2(n_48),
.Y(n_18)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_34),
.C(n_63),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B(n_31),
.Y(n_19)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_20),
.A2(n_30),
.B1(n_31),
.B2(n_98),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_20),
.A2(n_30),
.B1(n_31),
.B2(n_98),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

AO22x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_23),
.B(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_24),
.B(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

AOI22x1_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_29),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_27),
.B(n_139),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_33),
.A2(n_34),
.B1(n_96),
.B2(n_97),
.Y(n_155)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_34),
.B(n_96),
.C(n_154),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B(n_44),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_35),
.A2(n_39),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_40),
.Y(n_43)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_43),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_40),
.B(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_59),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_52),
.B(n_55),
.C(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_60),
.B1(n_61),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_55),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_74),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_73),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_67),
.A2(n_68),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_68),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_68),
.B(n_134),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_68),
.B(n_116),
.C(n_146),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.C(n_79),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_91),
.B1(n_112),
.B2(n_115),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_79),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_131),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_82),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_82),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_80),
.B(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_103),
.B2(n_104),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_97),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_125),
.B(n_163),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_110),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.C(n_117),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_137),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_116),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_117),
.B1(n_147),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_157),
.B(n_162),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_151),
.B(n_156),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_142),
.B(n_150),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_136),
.B(n_141),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_133),
.B(n_135),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_138),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_149),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_149),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_153),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_161),
.Y(n_162)
);


endmodule