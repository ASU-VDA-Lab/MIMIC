module fake_jpeg_10769_n_175 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_83),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_0),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_54),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_56),
.B(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_101),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_60),
.B1(n_58),
.B2(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_70),
.B1(n_66),
.B2(n_64),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_82),
.B(n_68),
.Y(n_101)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_75),
.B1(n_63),
.B2(n_62),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_109),
.B1(n_118),
.B2(n_5),
.Y(n_133)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_75),
.B1(n_63),
.B2(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_75),
.B(n_56),
.C(n_57),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_53),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_52),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_116),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_73),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_60),
.B1(n_58),
.B2(n_49),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_67),
.B1(n_59),
.B2(n_65),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_120),
.B1(n_57),
.B2(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_134),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_138),
.B(n_8),
.Y(n_151)
);

AO22x2_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_15),
.B1(n_43),
.B2(n_37),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_13),
.C(n_36),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_130),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_12),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_6),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_6),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_136),
.B(n_141),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_44),
.B1(n_25),
.B2(n_26),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_7),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_128),
.B(n_127),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_148),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_140),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_151),
.B(n_153),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_156),
.B1(n_33),
.B2(n_35),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_23),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_31),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_138),
.B1(n_131),
.B2(n_135),
.C(n_129),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_161),
.A2(n_144),
.B(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_165),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_160),
.A2(n_145),
.B1(n_143),
.B2(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_164),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_166),
.B1(n_168),
.B2(n_161),
.C(n_145),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_157),
.B(n_159),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_173),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_150),
.Y(n_175)
);


endmodule