module real_aes_14748_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_892;
wire n_372;
wire n_528;
wire n_202;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_931;
wire n_683;
wire n_904;
wire n_174;
wire n_780;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_917;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g286 ( .A(n_0), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_1), .Y(n_139) );
OA21x2_ASAP7_75t_L g124 ( .A1(n_2), .A2(n_47), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g185 ( .A(n_2), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_3), .B(n_175), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_4), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_5), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_6), .B(n_322), .Y(n_637) );
AND2x2_ASAP7_75t_L g190 ( .A(n_7), .B(n_154), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_8), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_9), .B(n_263), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_10), .B(n_263), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_11), .B(n_576), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_12), .B(n_166), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_13), .B(n_147), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_14), .B(n_285), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_15), .Y(n_611) );
BUFx3_ASAP7_75t_L g131 ( .A(n_16), .Y(n_131) );
INVx1_ASAP7_75t_L g145 ( .A(n_16), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_17), .B(n_153), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_18), .B(n_162), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_19), .Y(n_634) );
BUFx10_ASAP7_75t_L g108 ( .A(n_20), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_21), .B(n_203), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_22), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_23), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_24), .B(n_563), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g302 ( .A(n_25), .B(n_129), .C(n_300), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_26), .B(n_203), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_27), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_28), .B(n_162), .Y(n_655) );
NAND2xp33_ASAP7_75t_L g566 ( .A(n_29), .B(n_134), .Y(n_566) );
INVx1_ASAP7_75t_L g151 ( .A(n_30), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_31), .A2(n_146), .B(n_164), .C(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_32), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_33), .B(n_141), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_34), .B(n_175), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_35), .B(n_231), .Y(n_626) );
INVx1_ASAP7_75t_L g549 ( .A(n_36), .Y(n_549) );
AND3x2_ASAP7_75t_L g916 ( .A(n_36), .B(n_103), .C(n_105), .Y(n_916) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_37), .B(n_265), .Y(n_264) );
AO221x1_ASAP7_75t_L g573 ( .A1(n_38), .A2(n_80), .B1(n_203), .B2(n_230), .C(n_277), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_39), .B(n_623), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_40), .B(n_143), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_41), .Y(n_913) );
AND2x4_ASAP7_75t_L g150 ( .A(n_42), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_43), .B(n_153), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_44), .B(n_254), .Y(n_282) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_45), .B(n_143), .C(n_146), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_46), .B(n_153), .Y(n_316) );
INVx1_ASAP7_75t_L g184 ( .A(n_47), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_48), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_49), .A2(n_174), .B(n_284), .C(n_287), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g109 ( .A1(n_50), .A2(n_110), .B1(n_111), .B2(n_892), .Y(n_109) );
INVx1_ASAP7_75t_L g892 ( .A(n_50), .Y(n_892) );
INVx1_ASAP7_75t_L g125 ( .A(n_51), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_52), .Y(n_608) );
A2O1A1Ixp33_ASAP7_75t_L g668 ( .A1(n_53), .A2(n_669), .B(n_670), .C(n_672), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_54), .B(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g671 ( .A(n_55), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_56), .B(n_254), .Y(n_639) );
AND2x4_ASAP7_75t_L g924 ( .A(n_57), .B(n_925), .Y(n_924) );
INVx3_ASAP7_75t_L g217 ( .A(n_58), .Y(n_217) );
NOR2xp67_ASAP7_75t_L g104 ( .A(n_59), .B(n_72), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_60), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g925 ( .A(n_61), .Y(n_925) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_62), .B(n_213), .Y(n_327) );
INVx1_ASAP7_75t_L g229 ( .A(n_63), .Y(n_229) );
AND2x2_ASAP7_75t_L g628 ( .A(n_64), .B(n_254), .Y(n_628) );
INVx1_ASAP7_75t_L g579 ( .A(n_65), .Y(n_579) );
AOI31xp33_ASAP7_75t_L g895 ( .A1(n_66), .A2(n_896), .A3(n_902), .B(n_904), .Y(n_895) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_66), .B(n_897), .Y(n_910) );
INVx1_ASAP7_75t_L g939 ( .A(n_66), .Y(n_939) );
INVx2_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_68), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_69), .B(n_133), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_70), .B(n_129), .Y(n_128) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_71), .A2(n_74), .B1(n_563), .B2(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_73), .B(n_146), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_75), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g278 ( .A(n_76), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_77), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_78), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_79), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g678 ( .A(n_81), .B(n_154), .Y(n_678) );
INVx1_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
BUFx3_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
INVx1_ASAP7_75t_L g180 ( .A(n_82), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_83), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g215 ( .A(n_84), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_85), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_86), .B(n_182), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_87), .B(n_165), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_88), .B(n_154), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g905 ( .A(n_89), .Y(n_905) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_90), .B(n_623), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_91), .B(n_254), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_92), .B(n_325), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_93), .Y(n_207) );
INVx1_ASAP7_75t_L g202 ( .A(n_94), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g660 ( .A(n_95), .Y(n_660) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_96), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_97), .B(n_213), .Y(n_319) );
AOI21xp33_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_917), .B(n_926), .Y(n_98) );
OAI21xp5_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_109), .B(n_893), .Y(n_99) );
BUFx4f_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OR2x6_ASAP7_75t_L g101 ( .A(n_102), .B(n_107), .Y(n_101) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_104), .B(n_549), .Y(n_901) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g900 ( .A(n_106), .Y(n_900) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_107), .B(n_937), .Y(n_936) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g911 ( .A(n_108), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_108), .B(n_916), .Y(n_915) );
OR2x6_ASAP7_75t_SL g930 ( .A(n_108), .B(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OAI22x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_544), .B1(n_545), .B2(n_550), .Y(n_112) );
INVx1_ASAP7_75t_L g903 ( .A(n_113), .Y(n_903) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_442), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_364), .C(n_415), .Y(n_114) );
OAI221xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_256), .B1(n_304), .B2(n_309), .C(n_333), .Y(n_115) );
AOI211xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_191), .B(n_238), .C(n_246), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g539 ( .A(n_118), .B(n_242), .Y(n_539) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_156), .Y(n_118) );
INVx1_ASAP7_75t_L g240 ( .A(n_119), .Y(n_240) );
AND2x2_ASAP7_75t_L g394 ( .A(n_119), .B(n_340), .Y(n_394) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_119), .Y(n_439) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g249 ( .A(n_120), .Y(n_249) );
INVx3_ASAP7_75t_L g342 ( .A(n_120), .Y(n_342) );
AND2x2_ASAP7_75t_L g370 ( .A(n_120), .B(n_251), .Y(n_370) );
AND2x2_ASAP7_75t_L g377 ( .A(n_120), .B(n_378), .Y(n_377) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_126), .B(n_152), .Y(n_121) );
OAI21x1_ASAP7_75t_L g222 ( .A1(n_122), .A2(n_223), .B(n_237), .Y(n_222) );
OAI21x1_ASAP7_75t_L g631 ( .A1(n_122), .A2(n_632), .B(n_639), .Y(n_631) );
BUFx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVxp67_ASAP7_75t_L g661 ( .A(n_123), .Y(n_661) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g155 ( .A(n_124), .Y(n_155) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_124), .Y(n_254) );
INVx1_ASAP7_75t_L g186 ( .A(n_125), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_138), .B(n_148), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_132), .B(n_135), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g231 ( .A(n_130), .Y(n_231) );
INVx2_ASAP7_75t_L g563 ( .A(n_130), .Y(n_563) );
INVx2_ASAP7_75t_L g623 ( .A(n_130), .Y(n_623) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_131), .Y(n_134) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_131), .Y(n_209) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g141 ( .A(n_134), .Y(n_141) );
INVx3_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
INVx2_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
INVx2_ASAP7_75t_L g263 ( .A(n_134), .Y(n_263) );
INVx3_ASAP7_75t_L g277 ( .A(n_134), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_135), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_135), .A2(n_268), .B(n_269), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_135), .A2(n_626), .B(n_627), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_135), .A2(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g677 ( .A(n_135), .Y(n_677) );
BUFx10_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g300 ( .A(n_136), .Y(n_300) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx3_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
O2A1O1Ixp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_142), .C(n_146), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_140), .A2(n_657), .B(n_658), .Y(n_656) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
INVx2_ASAP7_75t_L g322 ( .A(n_144), .Y(n_322) );
INVx1_ASAP7_75t_L g326 ( .A(n_144), .Y(n_326) );
INVx1_ASAP7_75t_L g609 ( .A(n_144), .Y(n_609) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g167 ( .A(n_145), .Y(n_167) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_147), .B(n_205), .Y(n_204) );
NOR3xp33_ASAP7_75t_L g214 ( .A(n_147), .B(n_205), .C(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g230 ( .A(n_147), .Y(n_230) );
INVx1_ASAP7_75t_L g592 ( .A(n_147), .Y(n_592) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_148), .A2(n_294), .B(n_298), .Y(n_293) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_SL g331 ( .A(n_149), .Y(n_331) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g189 ( .A(n_150), .Y(n_189) );
INVx3_ASAP7_75t_L g205 ( .A(n_150), .Y(n_205) );
BUFx6f_ASAP7_75t_SL g236 ( .A(n_150), .Y(n_236) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_153), .Y(n_292) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OR2x2_ASAP7_75t_L g351 ( .A(n_157), .B(n_308), .Y(n_351) );
AO31x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_181), .A3(n_187), .B(n_190), .Y(n_157) );
AO31x2_ASAP7_75t_L g362 ( .A1(n_158), .A2(n_181), .A3(n_187), .B(n_190), .Y(n_362) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_159), .A2(n_252), .B(n_255), .Y(n_251) );
AOI22x1_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_169), .B1(n_170), .B2(n_177), .Y(n_159) );
OAI22x1_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B1(n_164), .B2(n_168), .Y(n_160) );
INVxp67_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g265 ( .A(n_166), .Y(n_265) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_166), .Y(n_280) );
INVx2_ASAP7_75t_L g297 ( .A(n_166), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_166), .B(n_611), .Y(n_610) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_167), .Y(n_203) );
INVx1_ASAP7_75t_L g287 ( .A(n_169), .Y(n_287) );
AOI21x1_ASAP7_75t_L g294 ( .A1(n_169), .A2(n_295), .B(n_296), .Y(n_294) );
AOI21xp5_ASAP7_75t_SL g619 ( .A1(n_169), .A2(n_620), .B(n_621), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .B1(n_174), .B2(n_176), .Y(n_170) );
INVxp67_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVxp67_ASAP7_75t_L g225 ( .A(n_172), .Y(n_225) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21x1_ASAP7_75t_SL g275 ( .A1(n_177), .A2(n_276), .B(n_279), .Y(n_275) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_178), .A2(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_178), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g211 ( .A(n_179), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_179), .A2(n_561), .B(n_562), .Y(n_560) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx3_ASAP7_75t_L g266 ( .A(n_180), .Y(n_266) );
INVxp67_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OAI21xp33_ASAP7_75t_L g288 ( .A1(n_182), .A2(n_189), .B(n_282), .Y(n_288) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_183), .B(n_331), .Y(n_600) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .Y(n_183) );
AOI21x1_ASAP7_75t_L g198 ( .A1(n_184), .A2(n_185), .B(n_186), .Y(n_198) );
BUFx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g255 ( .A(n_190), .Y(n_255) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI322xp5_ASAP7_75t_L g365 ( .A1(n_192), .A2(n_366), .A3(n_370), .B1(n_371), .B2(n_374), .C1(n_381), .C2(n_389), .Y(n_365) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g389 ( .A(n_194), .B(n_341), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_194), .B(n_341), .Y(n_404) );
AND2x2_ASAP7_75t_L g457 ( .A(n_194), .B(n_370), .Y(n_457) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_221), .Y(n_194) );
INVx3_ASAP7_75t_L g244 ( .A(n_195), .Y(n_244) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_199), .B(n_219), .Y(n_195) );
AO21x1_ASAP7_75t_L g379 ( .A1(n_196), .A2(n_199), .B(n_219), .Y(n_379) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_SL g219 ( .A(n_197), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_197), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_R g577 ( .A(n_198), .B(n_205), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_212), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_204), .B1(n_206), .B2(n_210), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
INVx1_ASAP7_75t_L g218 ( .A(n_203), .Y(n_218) );
INVx2_ASAP7_75t_L g270 ( .A(n_203), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_205), .B(n_211), .Y(n_210) );
NOR3xp33_ASAP7_75t_L g216 ( .A(n_205), .B(n_211), .C(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g567 ( .A(n_205), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_205), .B(n_254), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
INVx2_ASAP7_75t_L g213 ( .A(n_208), .Y(n_213) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g235 ( .A(n_209), .Y(n_235) );
INVx2_ASAP7_75t_L g285 ( .A(n_209), .Y(n_285) );
INVx2_ASAP7_75t_L g576 ( .A(n_209), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B1(n_216), .B2(n_218), .Y(n_212) );
INVx1_ASAP7_75t_L g245 ( .A(n_221), .Y(n_245) );
AND2x2_ASAP7_75t_L g250 ( .A(n_221), .B(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g308 ( .A(n_221), .Y(n_308) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_221), .Y(n_399) );
INVx2_ASAP7_75t_L g412 ( .A(n_221), .Y(n_412) );
AND2x2_ASAP7_75t_L g422 ( .A(n_221), .B(n_244), .Y(n_422) );
INVx1_ASAP7_75t_L g483 ( .A(n_221), .Y(n_483) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_232), .B(n_236), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_227), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_231), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx1_ASAP7_75t_L g588 ( .A(n_230), .Y(n_588) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_236), .A2(n_261), .B(n_267), .Y(n_260) );
OAI21x1_ASAP7_75t_L g632 ( .A1(n_236), .A2(n_633), .B(n_636), .Y(n_632) );
NOR2xp67_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g500 ( .A(n_240), .Y(n_500) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g526 ( .A(n_243), .B(n_361), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g340 ( .A(n_244), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_244), .B(n_342), .Y(n_363) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_248), .B(n_250), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_248), .B(n_448), .Y(n_472) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NOR2xp67_ASAP7_75t_L g306 ( .A(n_249), .B(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g431 ( .A(n_250), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g341 ( .A(n_251), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g450 ( .A(n_251), .Y(n_450) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_252), .A2(n_260), .B(n_271), .Y(n_259) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_252), .A2(n_260), .B(n_271), .Y(n_312) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2x1_ASAP7_75t_SL g329 ( .A(n_253), .B(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g349 ( .A(n_254), .Y(n_349) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_254), .Y(n_583) );
INVx2_ASAP7_75t_L g618 ( .A(n_254), .Y(n_618) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_272), .Y(n_256) );
AND2x2_ASAP7_75t_L g356 ( .A(n_257), .B(n_314), .Y(n_356) );
OR2x2_ASAP7_75t_L g523 ( .A(n_257), .B(n_354), .Y(n_523) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g336 ( .A(n_258), .B(n_337), .Y(n_336) );
BUFx3_ASAP7_75t_L g368 ( .A(n_258), .Y(n_368) );
AND2x2_ASAP7_75t_L g495 ( .A(n_258), .B(n_273), .Y(n_495) );
AND2x4_ASAP7_75t_L g511 ( .A(n_258), .B(n_408), .Y(n_511) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_259), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_264), .B(n_266), .Y(n_261) );
INVx2_ASAP7_75t_L g328 ( .A(n_266), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_266), .A2(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g672 ( .A(n_266), .Y(n_672) );
INVxp67_ASAP7_75t_L g301 ( .A(n_270), .Y(n_301) );
OR2x2_ASAP7_75t_L g372 ( .A(n_272), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g419 ( .A(n_272), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_289), .Y(n_272) );
AND2x4_ASAP7_75t_L g311 ( .A(n_273), .B(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_273), .Y(n_358) );
INVx1_ASAP7_75t_L g384 ( .A(n_273), .Y(n_384) );
AND2x2_ASAP7_75t_L g427 ( .A(n_273), .B(n_347), .Y(n_427) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g346 ( .A(n_274), .Y(n_346) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_281), .B(n_288), .Y(n_274) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x4_ASAP7_75t_L g388 ( .A(n_289), .B(n_314), .Y(n_388) );
INVx1_ASAP7_75t_L g402 ( .A(n_289), .Y(n_402) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_290), .Y(n_332) );
INVx2_ASAP7_75t_L g355 ( .A(n_290), .Y(n_355) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B(n_303), .Y(n_291) );
OA21x2_ASAP7_75t_L g347 ( .A1(n_293), .A2(n_303), .B(n_348), .Y(n_347) );
O2A1O1Ixp5_ASAP7_75t_L g633 ( .A1(n_297), .A2(n_592), .B(n_634), .C(n_635), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .B(n_302), .Y(n_298) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g469 ( .A(n_307), .B(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g490 ( .A(n_307), .Y(n_490) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_308), .B(n_479), .Y(n_493) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g400 ( .A(n_311), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g463 ( .A(n_311), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g488 ( .A(n_311), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g532 ( .A(n_311), .Y(n_532) );
AND2x2_ASAP7_75t_L g385 ( .A(n_312), .B(n_355), .Y(n_385) );
AND2x4_ASAP7_75t_L g387 ( .A(n_312), .B(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g392 ( .A(n_312), .B(n_345), .Y(n_392) );
AND2x4_ASAP7_75t_L g407 ( .A(n_312), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_332), .Y(n_313) );
INVx2_ASAP7_75t_L g337 ( .A(n_314), .Y(n_337) );
INVx2_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
BUFx2_ASAP7_75t_L g373 ( .A(n_314), .Y(n_373) );
INVx1_ASAP7_75t_L g429 ( .A(n_314), .Y(n_429) );
AND2x2_ASAP7_75t_L g489 ( .A(n_314), .B(n_347), .Y(n_489) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2x1_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
OAI21x1_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_323), .B(n_329), .Y(n_317) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B(n_328), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g369 ( .A(n_332), .B(n_337), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_343), .B(n_350), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_336), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g512 ( .A(n_336), .Y(n_512) );
AND2x2_ASAP7_75t_L g524 ( .A(n_336), .B(n_344), .Y(n_524) );
BUFx2_ASAP7_75t_L g464 ( .A(n_337), .Y(n_464) );
INVx1_ASAP7_75t_L g538 ( .A(n_337), .Y(n_538) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_341), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g413 ( .A(n_341), .Y(n_413) );
INVx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_344), .A2(n_535), .B1(n_537), .B2(n_539), .Y(n_534) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_SL g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OR2x6_ASAP7_75t_L g354 ( .A(n_346), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g408 ( .A(n_346), .Y(n_408) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_348), .A2(n_559), .B(n_568), .Y(n_558) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_357), .B2(n_360), .Y(n_350) );
INVx2_ASAP7_75t_SL g395 ( .A(n_351), .Y(n_395) );
OR2x2_ASAP7_75t_L g424 ( .A(n_351), .B(n_363), .Y(n_424) );
INVx2_ASAP7_75t_L g461 ( .A(n_352), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_353), .B(n_356), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g509 ( .A(n_354), .B(n_359), .Y(n_509) );
OR2x2_ASAP7_75t_L g542 ( .A(n_354), .B(n_368), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g430 ( .A(n_358), .B(n_385), .Y(n_430) );
INVx1_ASAP7_75t_L g406 ( .A(n_359), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_359), .B(n_383), .Y(n_446) );
OR2x2_ASAP7_75t_L g482 ( .A(n_359), .B(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g479 ( .A(n_361), .Y(n_479) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g380 ( .A(n_362), .Y(n_380) );
INVx1_ASAP7_75t_L g432 ( .A(n_363), .Y(n_432) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_363), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_390), .Y(n_364) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx2_ASAP7_75t_L g436 ( .A(n_368), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_368), .B(n_388), .Y(n_441) );
AND2x2_ASAP7_75t_L g454 ( .A(n_369), .B(n_455), .Y(n_454) );
BUFx3_ASAP7_75t_L g514 ( .A(n_369), .Y(n_514) );
INVx1_ASAP7_75t_L g516 ( .A(n_370), .Y(n_516) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g494 ( .A(n_373), .B(n_495), .Y(n_494) );
NAND2x1_ASAP7_75t_L g480 ( .A(n_374), .B(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g507 ( .A(n_375), .Y(n_507) );
OR2x6_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g470 ( .A(n_377), .Y(n_470) );
AND2x2_ASAP7_75t_L g530 ( .A(n_377), .B(n_380), .Y(n_530) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g411 ( .A(n_379), .B(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_379), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_380), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g521 ( .A(n_380), .Y(n_521) );
NAND2x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_386), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_383), .Y(n_484) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI221x1_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B1(n_396), .B2(n_400), .C(n_403), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_393), .A2(n_426), .B1(n_430), .B2(n_431), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_393), .A2(n_434), .B1(n_437), .B2(n_440), .Y(n_433) );
INVxp67_ASAP7_75t_SL g531 ( .A(n_393), .Y(n_531) );
AND2x4_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g471 ( .A(n_398), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_SL g414 ( .A(n_401), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_401), .B(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_409), .B2(n_414), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
AND2x4_ASAP7_75t_L g474 ( .A(n_406), .B(n_419), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_407), .A2(n_417), .B1(n_420), .B2(n_423), .Y(n_416) );
AND2x2_ASAP7_75t_L g497 ( .A(n_407), .B(n_464), .Y(n_497) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_413), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g478 ( .A(n_411), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g499 ( .A(n_411), .Y(n_499) );
AND2x2_ASAP7_75t_L g520 ( .A(n_411), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g537 ( .A(n_411), .B(n_538), .Y(n_537) );
NAND3xp33_ASAP7_75t_SL g415 ( .A(n_416), .B(n_425), .C(n_433), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_422), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g468 ( .A(n_430), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_431), .A2(n_492), .B(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g536 ( .A(n_439), .Y(n_536) );
INVx1_ASAP7_75t_L g452 ( .A(n_440), .Y(n_452) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_501), .Y(n_442) );
NAND3xp33_ASAP7_75t_SL g443 ( .A(n_444), .B(n_458), .C(n_475), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_447), .B(n_451), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_456), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g535 ( .A1(n_455), .A2(n_510), .B1(n_521), .B2(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g543 ( .A(n_455), .Y(n_543) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_465), .B(n_467), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_471), .B2(n_473), .Y(n_467) );
INVx1_ASAP7_75t_L g487 ( .A(n_470), .Y(n_487) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_474), .A2(n_498), .B(n_518), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_484), .B(n_485), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_480), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_481), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g506 ( .A(n_483), .Y(n_506) );
NAND3xp33_ASAP7_75t_SL g485 ( .A(n_486), .B(n_491), .C(n_496), .Y(n_485) );
NAND3xp33_ASAP7_75t_SL g486 ( .A(n_487), .B(n_488), .C(n_490), .Y(n_486) );
AND2x2_ASAP7_75t_L g518 ( .A(n_489), .B(n_511), .Y(n_518) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND3xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .C(n_500), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_527), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_508), .B(n_515), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2x1p5_ASAP7_75t_L g504 ( .A(n_505), .B(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND4xp25_ASAP7_75t_SL g508 ( .A(n_509), .B(n_510), .C(n_512), .D(n_513), .Y(n_508) );
INVx3_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OAI21xp5_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_517), .B(n_519), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_522), .B1(n_524), .B2(n_525), .Y(n_519) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
AOI21xp5_ASAP7_75t_SL g528 ( .A1(n_529), .A2(n_531), .B(n_532), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_530), .A2(n_539), .B1(n_541), .B2(n_543), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_534), .B(n_540), .Y(n_533) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_545), .Y(n_544) );
CKINVDCx10_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
BUFx6f_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND4xp75_ASAP7_75t_L g551 ( .A(n_552), .B(n_743), .C(n_810), .D(n_852), .Y(n_551) );
NOR3x1_ASAP7_75t_L g552 ( .A(n_553), .B(n_696), .C(n_737), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AOI211x1_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_594), .B(n_640), .C(n_680), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_569), .Y(n_555) );
OAI32xp33_ASAP7_75t_L g640 ( .A1(n_556), .A2(n_641), .A3(n_645), .B1(n_648), .B2(n_663), .Y(n_640) );
INVx2_ASAP7_75t_SL g850 ( .A(n_556), .Y(n_850) );
AND2x4_ASAP7_75t_L g867 ( .A(n_556), .B(n_739), .Y(n_867) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g662 ( .A(n_558), .B(n_580), .Y(n_662) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_558), .Y(n_695) );
INVx1_ASAP7_75t_L g701 ( .A(n_558), .Y(n_701) );
INVx1_ASAP7_75t_L g717 ( .A(n_558), .Y(n_717) );
AND2x2_ASAP7_75t_L g725 ( .A(n_558), .B(n_651), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_558), .B(n_580), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_564), .B(n_567), .Y(n_559) );
AND2x4_ASAP7_75t_L g617 ( .A(n_567), .B(n_618), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g679 ( .A1(n_567), .A2(n_661), .B(n_678), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g804 ( .A1(n_569), .A2(n_724), .B(n_805), .C(n_809), .Y(n_804) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g647 ( .A(n_571), .Y(n_647) );
OR2x2_ASAP7_75t_L g715 ( .A(n_571), .B(n_716), .Y(n_715) );
NOR2x1_ASAP7_75t_L g771 ( .A(n_571), .B(n_650), .Y(n_771) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_580), .Y(n_571) );
INVx2_ASAP7_75t_SL g689 ( .A(n_572), .Y(n_689) );
AND2x2_ASAP7_75t_L g702 ( .A(n_572), .B(n_693), .Y(n_702) );
AND2x2_ASAP7_75t_L g711 ( .A(n_572), .B(n_694), .Y(n_711) );
AND2x2_ASAP7_75t_L g728 ( .A(n_572), .B(n_691), .Y(n_728) );
BUFx3_ASAP7_75t_L g756 ( .A(n_572), .Y(n_756) );
AND2x2_ASAP7_75t_L g851 ( .A(n_572), .B(n_690), .Y(n_851) );
OR2x2_ASAP7_75t_L g884 ( .A(n_572), .B(n_701), .Y(n_884) );
AO31x2_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .A3(n_577), .B(n_578), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_576), .B(n_604), .Y(n_603) );
INVx3_ASAP7_75t_L g691 ( .A(n_580), .Y(n_691) );
AND2x2_ASAP7_75t_L g700 ( .A(n_580), .B(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_589), .B(n_593), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_588), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_588), .A2(n_607), .B(n_610), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_592), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_592), .A2(n_654), .B(n_655), .Y(n_653) );
INVxp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_613), .Y(n_595) );
AND2x4_ASAP7_75t_L g721 ( .A(n_596), .B(n_722), .Y(n_721) );
AND2x4_ASAP7_75t_L g741 ( .A(n_596), .B(n_742), .Y(n_741) );
NAND2x1_ASAP7_75t_L g820 ( .A(n_596), .B(n_757), .Y(n_820) );
INVx5_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_SL g646 ( .A(n_597), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g761 ( .A(n_597), .B(n_756), .Y(n_761) );
AND2x4_ASAP7_75t_L g765 ( .A(n_597), .B(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g790 ( .A(n_597), .B(n_666), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_597), .B(n_613), .Y(n_881) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVxp67_ASAP7_75t_L g736 ( .A(n_598), .Y(n_736) );
AO21x1_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_601), .B(n_605), .Y(n_598) );
AO21x2_ASAP7_75t_L g750 ( .A1(n_599), .A2(n_601), .B(n_605), .Y(n_750) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
OAI21x1_ASAP7_75t_SL g605 ( .A1(n_600), .A2(n_606), .B(n_612), .Y(n_605) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g669 ( .A(n_609), .Y(n_669) );
INVx1_ASAP7_75t_L g708 ( .A(n_613), .Y(n_708) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_629), .Y(n_613) );
INVx3_ASAP7_75t_L g705 ( .A(n_614), .Y(n_705) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g643 ( .A(n_615), .Y(n_643) );
OR2x2_ASAP7_75t_L g683 ( .A(n_615), .B(n_667), .Y(n_683) );
AND2x2_ASAP7_75t_L g759 ( .A(n_615), .B(n_631), .Y(n_759) );
AND2x2_ASAP7_75t_L g877 ( .A(n_615), .B(n_630), .Y(n_877) );
NAND2x1p5_ASAP7_75t_L g615 ( .A(n_616), .B(n_624), .Y(n_615) );
NAND2x1_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
AOI21x1_ASAP7_75t_L g624 ( .A1(n_617), .A2(n_625), .B(n_628), .Y(n_624) );
O2A1O1Ixp5_ASAP7_75t_L g652 ( .A1(n_617), .A2(n_653), .B(n_656), .C(n_659), .Y(n_652) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g664 ( .A(n_629), .Y(n_664) );
OR2x2_ASAP7_75t_L g729 ( .A(n_629), .B(n_683), .Y(n_729) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g644 ( .A(n_630), .Y(n_644) );
INVx1_ASAP7_75t_L g685 ( .A(n_630), .Y(n_685) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVxp33_ASAP7_75t_L g723 ( .A(n_631), .Y(n_723) );
OR2x2_ASAP7_75t_L g809 ( .A(n_641), .B(n_803), .Y(n_809) );
INVx1_ASAP7_75t_L g842 ( .A(n_641), .Y(n_842) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
AND2x2_ASAP7_75t_L g766 ( .A(n_642), .B(n_667), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_642), .B(n_707), .Y(n_808) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g666 ( .A(n_643), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g706 ( .A(n_644), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g823 ( .A(n_644), .B(n_750), .Y(n_823) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g815 ( .A(n_646), .B(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g870 ( .A(n_647), .B(n_650), .Y(n_870) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g760 ( .A(n_649), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_662), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_650), .B(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g814 ( .A(n_650), .Y(n_814) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g694 ( .A(n_651), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_651), .B(n_717), .Y(n_716) );
BUFx2_ASAP7_75t_SL g828 ( .A(n_651), .Y(n_828) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
AND2x4_ASAP7_75t_SL g773 ( .A(n_662), .B(n_689), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_662), .B(n_756), .Y(n_799) );
AND2x2_ASAP7_75t_L g827 ( .A(n_662), .B(n_828), .Y(n_827) );
OR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
AND2x2_ASAP7_75t_L g769 ( .A(n_664), .B(n_666), .Y(n_769) );
AND2x2_ASAP7_75t_L g777 ( .A(n_664), .B(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g817 ( .A(n_664), .Y(n_817) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_666), .B(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g707 ( .A(n_667), .Y(n_707) );
INVx2_ASAP7_75t_L g714 ( .A(n_667), .Y(n_714) );
INVx1_ASAP7_75t_L g780 ( .A(n_667), .Y(n_780) );
AND2x2_ASAP7_75t_L g886 ( .A(n_667), .B(n_749), .Y(n_886) );
AO21x2_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_673), .B(n_679), .Y(n_667) );
NOR2xp67_ASAP7_75t_L g670 ( .A(n_669), .B(n_671), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_677), .B(n_678), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
AOI21x1_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B(n_686), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x4_ASAP7_75t_SL g742 ( .A(n_682), .B(n_685), .Y(n_742) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g747 ( .A(n_683), .Y(n_747) );
BUFx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_685), .B(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g838 ( .A(n_685), .Y(n_838) );
OR2x2_ASAP7_75t_L g861 ( .A(n_685), .B(n_808), .Y(n_861) );
OR2x6_ASAP7_75t_L g686 ( .A(n_687), .B(n_692), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_688), .Y(n_854) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
AND2x2_ASAP7_75t_L g833 ( .A(n_689), .B(n_796), .Y(n_833) );
INVx1_ASAP7_75t_L g753 ( .A(n_690), .Y(n_753) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_691), .B(n_694), .Y(n_740) );
INVx1_ASAP7_75t_L g856 ( .A(n_692), .Y(n_856) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g734 ( .A(n_693), .Y(n_734) );
AND2x2_ASAP7_75t_L g786 ( .A(n_693), .B(n_773), .Y(n_786) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2x1_ASAP7_75t_L g696 ( .A(n_697), .B(n_718), .Y(n_696) );
OA222x2_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_703), .B1(n_708), .B2(n_709), .C1(n_712), .C2(n_715), .Y(n_697) );
INVx3_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI21xp33_ASAP7_75t_L g871 ( .A1(n_699), .A2(n_872), .B(n_874), .Y(n_871) );
AND2x4_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
AND2x4_ASAP7_75t_L g710 ( .A(n_700), .B(n_711), .Y(n_710) );
NAND2x1_ASAP7_75t_L g733 ( .A(n_700), .B(n_734), .Y(n_733) );
OAI21xp5_ASAP7_75t_L g818 ( .A1(n_700), .A2(n_819), .B(n_821), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_703), .A2(n_768), .B1(n_770), .B2(n_772), .Y(n_767) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND2x4_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
NAND2x1p5_ASAP7_75t_L g735 ( .A(n_705), .B(n_736), .Y(n_735) );
INVx4_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g731 ( .A(n_711), .B(n_732), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_711), .A2(n_821), .B1(n_888), .B2(n_889), .Y(n_887) );
NOR2xp33_ASAP7_75t_SL g847 ( .A(n_712), .B(n_838), .Y(n_847) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2x1_ASAP7_75t_L g831 ( .A(n_713), .B(n_757), .Y(n_831) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g722 ( .A(n_714), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g782 ( .A(n_714), .B(n_749), .Y(n_782) );
OR2x2_ASAP7_75t_L g803 ( .A(n_714), .B(n_749), .Y(n_803) );
INVx2_ASAP7_75t_L g796 ( .A(n_716), .Y(n_796) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI322xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_724), .A3(n_726), .B1(n_729), .B2(n_730), .C1(n_733), .C2(n_735), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g748 ( .A(n_723), .B(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g858 ( .A(n_724), .B(n_859), .Y(n_858) );
INVx2_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
AND2x4_ASAP7_75t_L g784 ( .A(n_725), .B(n_728), .Y(n_784) );
AO221x1_ASAP7_75t_L g853 ( .A1(n_726), .A2(n_850), .B1(n_854), .B2(n_855), .C(n_857), .Y(n_853) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g839 ( .A(n_728), .B(n_796), .Y(n_839) );
AOI21xp5_ASAP7_75t_SL g763 ( .A1(n_730), .A2(n_758), .B(n_764), .Y(n_763) );
INVx4_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_731), .A2(n_777), .B1(n_847), .B2(n_848), .Y(n_846) );
AND2x2_ASAP7_75t_L g888 ( .A(n_734), .B(n_851), .Y(n_888) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_741), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI21xp5_ASAP7_75t_L g834 ( .A1(n_742), .A2(n_835), .B(n_839), .Y(n_834) );
INVx2_ASAP7_75t_L g844 ( .A(n_742), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_742), .A2(n_864), .B1(n_865), .B2(n_868), .Y(n_863) );
NOR3x1_ASAP7_75t_L g743 ( .A(n_744), .B(n_774), .C(n_797), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_762), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_751), .B1(n_757), .B2(n_760), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g793 ( .A(n_747), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_748), .B(n_793), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_748), .B(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_748), .B(n_891), .Y(n_890) );
INVx2_ASAP7_75t_L g807 ( .A(n_749), .Y(n_807) );
INVx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_750), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_753), .B(n_796), .Y(n_795) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_754), .Y(n_873) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g859 ( .A(n_756), .Y(n_859) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_756), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_757), .B(n_802), .Y(n_801) );
INVx6_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx4_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g885 ( .A(n_759), .B(n_886), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_761), .B(n_827), .Y(n_845) );
NOR2xp67_ASAP7_75t_SL g762 ( .A(n_763), .B(n_767), .Y(n_762) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OAI21xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_783), .B(n_785), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_776), .B(n_781), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g837 ( .A(n_778), .Y(n_837) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g788 ( .A(n_782), .Y(n_788) );
INVxp67_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_787), .B1(n_791), .B2(n_794), .Y(n_785) );
INVx2_ASAP7_75t_L g843 ( .A(n_786), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
INVx2_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
INVxp67_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
AO21x1_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_800), .B(n_804), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVxp67_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g864 ( .A(n_805), .Y(n_864) );
OR2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_808), .Y(n_805) );
OR2x2_ASAP7_75t_L g875 ( .A(n_806), .B(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
BUFx2_ASAP7_75t_SL g830 ( .A(n_807), .Y(n_830) );
OR2x2_ASAP7_75t_L g829 ( .A(n_808), .B(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g891 ( .A(n_808), .Y(n_891) );
NOR2x1_ASAP7_75t_L g810 ( .A(n_811), .B(n_840), .Y(n_810) );
NAND4xp75_ASAP7_75t_L g811 ( .A(n_812), .B(n_818), .C(n_824), .D(n_834), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_815), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_829), .B1(n_831), .B2(n_832), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
OR2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_839), .A2(n_880), .B1(n_882), .B2(n_885), .Y(n_879) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_843), .B1(n_844), .B2(n_845), .C(n_846), .Y(n_840) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
AOI211x1_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_860), .B(n_862), .C(n_878), .Y(n_852) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_SL g862 ( .A(n_863), .B(n_871), .Y(n_862) );
AND2x4_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx2_ASAP7_75t_SL g869 ( .A(n_870), .Y(n_869) );
INVxp67_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
NAND2xp5_ASAP7_75t_SL g878 ( .A(n_879), .B(n_887), .Y(n_878) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
HB1xp67_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVxp67_ASAP7_75t_SL g889 ( .A(n_890), .Y(n_889) );
AOI21xp5_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_911), .B(n_912), .Y(n_893) );
INVxp67_ASAP7_75t_L g927 ( .A(n_894), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_895), .B(n_908), .Y(n_894) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVxp67_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_SL g907 ( .A(n_899), .Y(n_907) );
HB1xp67_ASAP7_75t_L g938 ( .A(n_899), .Y(n_938) );
NOR2x1p5_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
INVx2_ASAP7_75t_L g909 ( .A(n_902), .Y(n_909) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NOR2x1_ASAP7_75t_R g904 ( .A(n_905), .B(n_906), .Y(n_904) );
BUFx6f_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_907), .B(n_920), .Y(n_919) );
BUFx12f_ASAP7_75t_L g932 ( .A(n_907), .Y(n_932) );
NAND2xp5_ASAP7_75t_SL g908 ( .A(n_909), .B(n_910), .Y(n_908) );
NOR2xp33_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
BUFx6f_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
BUFx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
OR2x2_ASAP7_75t_L g935 ( .A(n_921), .B(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g931 ( .A(n_924), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_927), .A2(n_928), .B1(n_933), .B2(n_939), .Y(n_926) );
BUFx10_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
OR2x6_ASAP7_75t_L g929 ( .A(n_930), .B(n_932), .Y(n_929) );
INVx2_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
BUFx6f_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx2_ASAP7_75t_SL g937 ( .A(n_938), .Y(n_937) );
endmodule