module real_aes_349_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_815;
wire n_564;
wire n_638;
wire n_519;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_314;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
XNOR2x1_ASAP7_75t_L g740 ( .A(n_0), .B(n_741), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_1), .A2(n_258), .B1(n_479), .B2(n_480), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_2), .A2(n_215), .B1(n_443), .B2(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_3), .A2(n_266), .B1(n_488), .B2(n_577), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_4), .A2(n_156), .B1(n_398), .B2(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_5), .A2(n_80), .B1(n_400), .B2(n_500), .Y(n_499) );
AO22x2_ASAP7_75t_L g322 ( .A1(n_6), .A2(n_202), .B1(n_312), .B2(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g783 ( .A(n_6), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_7), .A2(n_203), .B1(n_442), .B2(n_443), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_8), .A2(n_259), .B1(n_475), .B2(n_524), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_9), .A2(n_118), .B1(n_341), .B2(n_439), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_10), .A2(n_168), .B1(n_515), .B2(n_652), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_11), .A2(n_182), .B1(n_419), .B2(n_652), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_12), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_13), .A2(n_252), .B1(n_350), .B2(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_14), .A2(n_183), .B1(n_406), .B2(n_408), .Y(n_405) );
AO22x2_ASAP7_75t_L g319 ( .A1(n_15), .A2(n_63), .B1(n_312), .B2(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_15), .B(n_782), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_16), .A2(n_239), .B1(n_433), .B2(n_434), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_17), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_18), .A2(n_282), .B1(n_356), .B2(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_19), .A2(n_92), .B1(n_472), .B2(n_473), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_20), .A2(n_138), .B1(n_406), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_21), .A2(n_187), .B1(n_439), .B2(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_22), .A2(n_235), .B1(n_486), .B2(n_705), .Y(n_704) );
AO222x2_ASAP7_75t_SL g520 ( .A1(n_23), .A2(n_48), .B1(n_163), .B2(n_449), .C1(n_452), .C2(n_521), .Y(n_520) );
AO22x2_ASAP7_75t_L g301 ( .A1(n_24), .A2(n_302), .B1(n_384), .B2(n_385), .Y(n_301) );
INVx1_ASAP7_75t_L g385 ( .A(n_24), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_25), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_26), .A2(n_89), .B1(n_439), .B2(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_27), .A2(n_280), .B1(n_331), .B2(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_28), .A2(n_69), .B1(n_417), .B2(n_419), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_29), .A2(n_157), .B1(n_442), .B2(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_30), .A2(n_211), .B1(n_372), .B2(n_375), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_31), .A2(n_165), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_32), .A2(n_219), .B1(n_326), .B2(n_331), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_33), .B(n_306), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_34), .A2(n_51), .B1(n_510), .B2(n_511), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_35), .A2(n_241), .B1(n_820), .B2(n_821), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_36), .A2(n_285), .B1(n_372), .B2(n_515), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_37), .A2(n_159), .B1(n_482), .B2(n_488), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_38), .A2(n_228), .B1(n_583), .B2(n_584), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_39), .A2(n_142), .B1(n_515), .B2(n_654), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_40), .A2(n_196), .B1(n_402), .B2(n_720), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_41), .A2(n_195), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_42), .A2(n_166), .B1(n_338), .B2(n_340), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_43), .A2(n_221), .B1(n_443), .B2(n_475), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_44), .A2(n_144), .B1(n_479), .B2(n_480), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_45), .A2(n_136), .B1(n_363), .B2(n_402), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_46), .A2(n_122), .B1(n_445), .B2(n_580), .Y(n_579) );
OAI22x1_ASAP7_75t_L g388 ( .A1(n_47), .A2(n_389), .B1(n_390), .B2(n_425), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_47), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_49), .A2(n_77), .B1(n_480), .B2(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_50), .A2(n_201), .B1(n_421), .B2(n_713), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_52), .A2(n_267), .B1(n_338), .B2(n_377), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_53), .A2(n_96), .B1(n_472), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_54), .A2(n_116), .B1(n_442), .B2(n_443), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_55), .A2(n_178), .B1(n_396), .B2(n_723), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_56), .A2(n_263), .B1(n_377), .B2(n_439), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_57), .A2(n_191), .B1(n_356), .B2(n_358), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_58), .A2(n_130), .B1(n_472), .B2(n_526), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_59), .A2(n_169), .B1(n_485), .B2(n_486), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_60), .A2(n_162), .B1(n_408), .B2(n_726), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_61), .A2(n_155), .B1(n_452), .B2(n_521), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_62), .A2(n_274), .B1(n_627), .B2(n_628), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_64), .A2(n_217), .B1(n_452), .B2(n_521), .Y(n_666) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_65), .A2(n_112), .B1(n_475), .B2(n_524), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_66), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_67), .B(n_393), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_68), .A2(n_265), .B1(n_410), .B2(n_414), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_70), .A2(n_236), .B1(n_379), .B2(n_381), .Y(n_378) );
AO222x2_ASAP7_75t_SL g792 ( .A1(n_71), .A2(n_194), .B1(n_220), .B2(n_449), .C1(n_452), .C2(n_521), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_72), .A2(n_120), .B1(n_624), .B2(n_815), .Y(n_814) );
OA22x2_ASAP7_75t_L g683 ( .A1(n_73), .A2(n_684), .B1(n_685), .B2(n_707), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_73), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_74), .A2(n_125), .B1(n_623), .B2(n_624), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_75), .A2(n_200), .B1(n_654), .B2(n_655), .Y(n_816) );
INVx3_ASAP7_75t_L g312 ( .A(n_76), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_78), .A2(n_149), .B1(n_485), .B2(n_486), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_79), .A2(n_227), .B1(n_345), .B2(n_350), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_81), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_82), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_83), .A2(n_245), .B1(n_452), .B2(n_521), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_84), .A2(n_207), .B1(n_482), .B2(n_534), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_85), .A2(n_197), .B1(n_363), .B2(n_367), .Y(n_818) );
OA22x2_ASAP7_75t_L g808 ( .A1(n_86), .A2(n_809), .B1(n_810), .B2(n_824), .Y(n_808) );
INVxp67_ASAP7_75t_L g824 ( .A(n_86), .Y(n_824) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_87), .A2(n_104), .B1(n_204), .B2(n_448), .C1(n_450), .C2(n_453), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_88), .A2(n_212), .B1(n_358), .B2(n_641), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_90), .A2(n_99), .B1(n_345), .B2(n_431), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_91), .B(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_93), .A2(n_255), .B1(n_479), .B2(n_480), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_94), .A2(n_137), .B1(n_446), .B2(n_503), .Y(n_746) );
INVx1_ASAP7_75t_SL g313 ( .A(n_95), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_95), .B(n_134), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_97), .A2(n_150), .B1(n_395), .B2(n_396), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_98), .A2(n_264), .B1(n_718), .B2(n_720), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_100), .A2(n_179), .B1(n_356), .B2(n_505), .Y(n_745) );
INVx2_ASAP7_75t_L g296 ( .A(n_101), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_102), .A2(n_261), .B1(n_350), .B2(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_103), .A2(n_131), .B1(n_398), .B2(n_400), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_105), .A2(n_287), .B1(n_297), .B2(n_785), .C(n_786), .Y(n_286) );
XOR2x2_ASAP7_75t_L g756 ( .A(n_106), .B(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_107), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_108), .A2(n_225), .B1(n_472), .B2(n_473), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_109), .A2(n_139), .B1(n_452), .B2(n_453), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_110), .A2(n_152), .B1(n_485), .B2(n_486), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_111), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_113), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_114), .A2(n_192), .B1(n_479), .B2(n_480), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_115), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_117), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_119), .B(n_646), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_121), .A2(n_256), .B1(n_445), .B2(n_446), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_123), .A2(n_185), .B1(n_446), .B2(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_124), .A2(n_158), .B1(n_514), .B2(n_515), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_126), .A2(n_270), .B1(n_406), .B2(n_408), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_127), .A2(n_206), .B1(n_488), .B2(n_535), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_128), .A2(n_272), .B1(n_731), .B2(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_129), .A2(n_184), .B1(n_479), .B2(n_480), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_132), .A2(n_205), .B1(n_417), .B2(n_729), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_133), .A2(n_146), .B1(n_372), .B2(n_381), .Y(n_813) );
AO22x2_ASAP7_75t_L g315 ( .A1(n_134), .A2(n_214), .B1(n_312), .B2(n_316), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_135), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_140), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_141), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_143), .A2(n_250), .B1(n_363), .B2(n_367), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_145), .A2(n_279), .B1(n_437), .B2(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_147), .A2(n_233), .B1(n_482), .B2(n_488), .Y(n_532) );
XOR2x2_ASAP7_75t_L g493 ( .A(n_148), .B(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_151), .A2(n_284), .B1(n_412), .B2(n_431), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_153), .A2(n_281), .B1(n_503), .B2(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_154), .A2(n_181), .B1(n_654), .B2(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g314 ( .A(n_160), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_161), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_164), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_167), .A2(n_234), .B1(n_338), .B2(n_437), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_170), .A2(n_262), .B1(n_433), .B2(n_511), .Y(n_750) );
AOI222xp33_ASAP7_75t_L g730 ( .A1(n_171), .A2(n_176), .B1(n_275), .B2(n_468), .C1(n_731), .C2(n_732), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_172), .A2(n_268), .B1(n_421), .B2(n_423), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_173), .A2(n_238), .B1(n_760), .B2(n_761), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_174), .A2(n_177), .B1(n_485), .B2(n_486), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_175), .B(n_468), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_180), .A2(n_193), .B1(n_331), .B2(n_648), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_186), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_188), .A2(n_209), .B1(n_485), .B2(n_486), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_189), .A2(n_251), .B1(n_345), .B2(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_190), .A2(n_248), .B1(n_482), .B2(n_488), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_198), .A2(n_230), .B1(n_345), .B2(n_431), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_199), .A2(n_254), .B1(n_534), .B2(n_535), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g471 ( .A1(n_208), .A2(n_216), .B1(n_472), .B2(n_473), .Y(n_471) );
OA22x2_ASAP7_75t_L g610 ( .A1(n_210), .A2(n_611), .B1(n_629), .B2(n_630), .Y(n_610) );
INVx1_ASAP7_75t_L g629 ( .A(n_210), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_213), .A2(n_231), .B1(n_400), .B2(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_218), .B(n_748), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_222), .A2(n_242), .B1(n_402), .B2(n_403), .Y(n_401) );
OAI22x1_ASAP7_75t_L g636 ( .A1(n_223), .A2(n_637), .B1(n_638), .B2(n_658), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_223), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_224), .B(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_226), .A2(n_276), .B1(n_439), .B2(n_482), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_229), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g779 ( .A(n_229), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_232), .Y(n_665) );
XOR2x2_ASAP7_75t_L g708 ( .A(n_237), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g293 ( .A(n_240), .Y(n_293) );
AND2x2_ASAP7_75t_R g807 ( .A(n_240), .B(n_779), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_243), .B(n_448), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_244), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_246), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_247), .B(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_249), .A2(n_278), .B1(n_423), .B2(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_253), .B(n_295), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_257), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_260), .A2(n_283), .B1(n_485), .B2(n_486), .Y(n_802) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_269), .B(n_468), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_271), .A2(n_788), .B1(n_789), .B2(n_803), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_271), .Y(n_803) );
OA22x2_ASAP7_75t_L g426 ( .A1(n_273), .A2(n_427), .B1(n_428), .B2(n_454), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_273), .Y(n_427) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_273), .A2(n_428), .B(n_458), .Y(n_457) );
XNOR2xp5_ASAP7_75t_L g660 ( .A(n_277), .B(n_661), .Y(n_660) );
CKINVDCx6p67_ASAP7_75t_R g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_SL g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g828 ( .A(n_292), .B(n_294), .Y(n_828) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_293), .B(n_779), .Y(n_778) );
AOI21xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_678), .B(n_776), .Y(n_297) );
OR2x2_ASAP7_75t_L g785 ( .A(n_298), .B(n_678), .Y(n_785) );
XNOR2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_461), .Y(n_298) );
OAI22xp33_ASAP7_75t_R g299 ( .A1(n_300), .A2(n_386), .B1(n_387), .B2(n_460), .Y(n_299) );
INVx1_ASAP7_75t_L g460 ( .A(n_300), .Y(n_460) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_SL g384 ( .A(n_302), .Y(n_384) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_353), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_336), .Y(n_303) );
OAI21xp33_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_324), .B(n_325), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_306), .Y(n_393) );
INVx3_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx4_ASAP7_75t_SL g468 ( .A(n_307), .Y(n_468) );
BUFx2_ASAP7_75t_L g497 ( .A(n_307), .Y(n_497) );
INVx3_ASAP7_75t_L g646 ( .A(n_307), .Y(n_646) );
INVx4_ASAP7_75t_SL g748 ( .A(n_307), .Y(n_748) );
INVx6_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_317), .Y(n_308) );
AND2x4_ASAP7_75t_L g360 ( .A(n_309), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g364 ( .A(n_309), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g443 ( .A(n_309), .B(n_361), .Y(n_443) );
AND2x4_ASAP7_75t_L g449 ( .A(n_309), .B(n_317), .Y(n_449) );
AND2x2_ASAP7_75t_L g473 ( .A(n_309), .B(n_365), .Y(n_473) );
AND2x2_ASAP7_75t_L g524 ( .A(n_309), .B(n_361), .Y(n_524) );
AND2x2_ASAP7_75t_L g526 ( .A(n_309), .B(n_365), .Y(n_526) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_315), .Y(n_309) );
AND2x2_ASAP7_75t_L g329 ( .A(n_310), .B(n_330), .Y(n_329) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_310), .Y(n_335) );
INVx2_ASAP7_75t_L g343 ( .A(n_310), .Y(n_343) );
OAI22x1_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B1(n_313), .B2(n_314), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g316 ( .A(n_312), .Y(n_316) );
INVx2_ASAP7_75t_L g320 ( .A(n_312), .Y(n_320) );
INVx1_ASAP7_75t_L g323 ( .A(n_312), .Y(n_323) );
INVx2_ASAP7_75t_L g330 ( .A(n_315), .Y(n_330) );
AND2x2_ASAP7_75t_L g349 ( .A(n_315), .B(n_343), .Y(n_349) );
BUFx2_ASAP7_75t_L g352 ( .A(n_315), .Y(n_352) );
AND2x4_ASAP7_75t_L g339 ( .A(n_317), .B(n_329), .Y(n_339) );
AND2x4_ASAP7_75t_L g374 ( .A(n_317), .B(n_342), .Y(n_374) );
AND2x2_ASAP7_75t_L g380 ( .A(n_317), .B(n_349), .Y(n_380) );
AND2x2_ASAP7_75t_L g485 ( .A(n_317), .B(n_329), .Y(n_485) );
AND2x6_ASAP7_75t_L g488 ( .A(n_317), .B(n_349), .Y(n_488) );
AND2x2_ASAP7_75t_L g534 ( .A(n_317), .B(n_342), .Y(n_534) );
AND2x2_ASAP7_75t_L g705 ( .A(n_317), .B(n_329), .Y(n_705) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_321), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g328 ( .A(n_319), .B(n_321), .Y(n_328) );
AND2x2_ASAP7_75t_L g334 ( .A(n_319), .B(n_322), .Y(n_334) );
INVx1_ASAP7_75t_L g348 ( .A(n_319), .Y(n_348) );
INVxp67_ASAP7_75t_L g361 ( .A(n_321), .Y(n_361) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g347 ( .A(n_322), .B(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_326), .Y(n_548) );
BUFx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g399 ( .A(n_327), .Y(n_399) );
BUFx3_ASAP7_75t_L g616 ( .A(n_327), .Y(n_616) );
BUFx5_ASAP7_75t_L g648 ( .A(n_327), .Y(n_648) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x4_ASAP7_75t_L g341 ( .A(n_328), .B(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g357 ( .A(n_328), .B(n_349), .Y(n_357) );
AND2x2_ASAP7_75t_L g442 ( .A(n_328), .B(n_349), .Y(n_442) );
AND2x4_ASAP7_75t_L g452 ( .A(n_328), .B(n_329), .Y(n_452) );
AND2x2_ASAP7_75t_L g475 ( .A(n_328), .B(n_349), .Y(n_475) );
AND2x2_ASAP7_75t_L g535 ( .A(n_328), .B(n_342), .Y(n_535) );
AND2x2_ASAP7_75t_L g369 ( .A(n_329), .B(n_347), .Y(n_369) );
AND2x4_ASAP7_75t_L g472 ( .A(n_329), .B(n_347), .Y(n_472) );
AND2x4_ASAP7_75t_L g342 ( .A(n_330), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g744 ( .A(n_332), .Y(n_744) );
INVx3_ASAP7_75t_L g766 ( .A(n_332), .Y(n_766) );
INVx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx12f_ASAP7_75t_L g400 ( .A(n_333), .Y(n_400) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x4_ASAP7_75t_L g351 ( .A(n_334), .B(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g377 ( .A(n_334), .B(n_342), .Y(n_377) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_334), .B(n_335), .Y(n_453) );
AND2x4_ASAP7_75t_L g480 ( .A(n_334), .B(n_352), .Y(n_480) );
AND2x4_ASAP7_75t_L g486 ( .A(n_334), .B(n_342), .Y(n_486) );
AND2x2_ASAP7_75t_SL g521 ( .A(n_334), .B(n_335), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_344), .Y(n_336) );
BUFx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx6_ASAP7_75t_L g407 ( .A(n_339), .Y(n_407) );
BUFx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g424 ( .A(n_341), .Y(n_424) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_341), .Y(n_515) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_341), .Y(n_577) );
AND2x4_ASAP7_75t_L g383 ( .A(n_342), .B(n_347), .Y(n_383) );
AND2x6_ASAP7_75t_L g482 ( .A(n_342), .B(n_347), .Y(n_482) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_345), .Y(n_557) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g413 ( .A(n_346), .Y(n_413) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_347), .B(n_349), .Y(n_479) );
AND2x2_ASAP7_75t_L g601 ( .A(n_347), .B(n_349), .Y(n_601) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_348), .Y(n_366) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx5_ASAP7_75t_SL g415 ( .A(n_351), .Y(n_415) );
BUFx2_ASAP7_75t_L g624 ( .A(n_351), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_370), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_362), .Y(n_354) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_357), .Y(n_395) );
BUFx2_ASAP7_75t_L g641 ( .A(n_357), .Y(n_641) );
BUFx2_ASAP7_75t_L g820 ( .A(n_357), .Y(n_820) );
INVx2_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g396 ( .A(n_359), .Y(n_396) );
INVx2_ASAP7_75t_L g505 ( .A(n_359), .Y(n_505) );
INVx2_ASAP7_75t_L g584 ( .A(n_359), .Y(n_584) );
INVx2_ASAP7_75t_L g761 ( .A(n_359), .Y(n_761) );
INVx1_ASAP7_75t_L g821 ( .A(n_359), .Y(n_821) );
INVx6_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx6f_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
BUFx4f_ASAP7_75t_L g403 ( .A(n_364), .Y(n_403) );
BUFx3_ASAP7_75t_L g446 ( .A(n_364), .Y(n_446) );
INVx1_ASAP7_75t_L g581 ( .A(n_364), .Y(n_581) );
INVx2_ASAP7_75t_L g644 ( .A(n_364), .Y(n_644) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx4_ASAP7_75t_L g445 ( .A(n_368), .Y(n_445) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_369), .Y(n_402) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_369), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_378), .Y(n_370) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx4_ASAP7_75t_L g418 ( .A(n_373), .Y(n_418) );
INVx3_ASAP7_75t_L g439 ( .A(n_373), .Y(n_439) );
INVx2_ASAP7_75t_SL g510 ( .A(n_373), .Y(n_510) );
INVx3_ASAP7_75t_SL g627 ( .A(n_373), .Y(n_627) );
INVx8_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_SL g655 ( .A(n_376), .Y(n_655) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_SL g408 ( .A(n_377), .Y(n_408) );
BUFx2_ASAP7_75t_SL g570 ( .A(n_377), .Y(n_570) );
BUFx3_ASAP7_75t_L g754 ( .A(n_377), .Y(n_754) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g422 ( .A(n_380), .Y(n_422) );
BUFx2_ASAP7_75t_L g514 ( .A(n_380), .Y(n_514) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g419 ( .A(n_382), .Y(n_419) );
INVx2_ASAP7_75t_L g434 ( .A(n_382), .Y(n_434) );
INVx2_ASAP7_75t_L g511 ( .A(n_382), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_382), .A2(n_560), .B1(n_561), .B2(n_564), .Y(n_559) );
INVx2_ASAP7_75t_SL g628 ( .A(n_382), .Y(n_628) );
INVx2_ASAP7_75t_L g713 ( .A(n_382), .Y(n_713) );
INVx8_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
OA22x2_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_426), .B1(n_455), .B2(n_456), .Y(n_387) );
INVx1_ASAP7_75t_SL g455 ( .A(n_388), .Y(n_455) );
INVx2_ASAP7_75t_SL g425 ( .A(n_390), .Y(n_425) );
OR2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_404), .Y(n_390) );
NAND4xp25_ASAP7_75t_SL g391 ( .A(n_392), .B(n_394), .C(n_397), .D(n_401), .Y(n_391) );
INVx3_ASAP7_75t_L g546 ( .A(n_393), .Y(n_546) );
BUFx2_ASAP7_75t_L g583 ( .A(n_395), .Y(n_583) );
BUFx4f_ASAP7_75t_SL g723 ( .A(n_395), .Y(n_723) );
BUFx2_ASAP7_75t_L g760 ( .A(n_395), .Y(n_760) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g500 ( .A(n_399), .Y(n_500) );
INVx2_ASAP7_75t_L g552 ( .A(n_400), .Y(n_552) );
BUFx3_ASAP7_75t_L g732 ( .A(n_400), .Y(n_732) );
INVx1_ASAP7_75t_L g692 ( .A(n_402), .Y(n_692) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_409), .C(n_416), .D(n_420), .Y(n_404) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_407), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_566) );
INVx3_ASAP7_75t_L g654 ( .A(n_407), .Y(n_654) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g715 ( .A(n_411), .Y(n_715) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_412), .Y(n_815) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g623 ( .A(n_413), .Y(n_623) );
INVx1_ASAP7_75t_L g772 ( .A(n_413), .Y(n_772) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g431 ( .A(n_415), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_415), .A2(n_555), .B1(n_556), .B2(n_558), .Y(n_554) );
INVx2_ASAP7_75t_L g657 ( .A(n_415), .Y(n_657) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g727 ( .A(n_418), .Y(n_727) );
INVx2_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g433 ( .A(n_422), .Y(n_433) );
INVx2_ASAP7_75t_L g563 ( .A(n_422), .Y(n_563) );
INVx2_ASAP7_75t_L g652 ( .A(n_422), .Y(n_652) );
INVx2_ASAP7_75t_SL g712 ( .A(n_422), .Y(n_712) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g437 ( .A(n_424), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_427), .Y(n_459) );
INVx1_ASAP7_75t_L g454 ( .A(n_428), .Y(n_454) );
NOR2x1_ASAP7_75t_SL g458 ( .A(n_428), .B(n_459), .Y(n_458) );
NAND4xp75_ASAP7_75t_L g428 ( .A(n_429), .B(n_435), .C(n_440), .D(n_447), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_444), .Y(n_440) );
INVxp67_ASAP7_75t_L g696 ( .A(n_442), .Y(n_696) );
INVx2_ASAP7_75t_SL g719 ( .A(n_445), .Y(n_719) );
BUFx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_SL g664 ( .A(n_449), .Y(n_664) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
XNOR2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_588), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_490), .B1(n_491), .B2(n_587), .Y(n_462) );
INVx1_ASAP7_75t_L g587 ( .A(n_463), .Y(n_587) );
XOR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_489), .Y(n_463) );
NAND2x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_476), .Y(n_464) );
NOR2x1_ASAP7_75t_L g465 ( .A(n_466), .B(n_470), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
BUFx2_ASAP7_75t_L g763 ( .A(n_468), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_474), .Y(n_470) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_483), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_481), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
INVx1_ASAP7_75t_L g621 ( .A(n_488), .Y(n_621) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI22x1_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_539), .B1(n_540), .B2(n_586), .Y(n_491) );
INVx2_ASAP7_75t_L g586 ( .A(n_492), .Y(n_586) );
AO22x2_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_517), .B1(n_537), .B2(n_538), .Y(n_492) );
INVx2_ASAP7_75t_L g538 ( .A(n_493), .Y(n_538) );
NAND2x1_ASAP7_75t_SL g494 ( .A(n_495), .B(n_506), .Y(n_494) );
NOR2x1_ASAP7_75t_L g495 ( .A(n_496), .B(n_501), .Y(n_495) );
OAI21xp5_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_498), .B(n_499), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_507), .B(n_512), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
BUFx2_ASAP7_75t_L g574 ( .A(n_510), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_516), .Y(n_512) );
INVx2_ASAP7_75t_L g537 ( .A(n_517), .Y(n_537) );
XOR2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_536), .Y(n_517) );
NAND2x1_ASAP7_75t_L g518 ( .A(n_519), .B(n_527), .Y(n_518) );
NOR2x1_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVxp67_ASAP7_75t_L g698 ( .A(n_524), .Y(n_698) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_531), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
XNOR2x1_ASAP7_75t_L g541 ( .A(n_542), .B(n_585), .Y(n_541) );
NAND4xp75_ASAP7_75t_L g542 ( .A(n_543), .B(n_553), .C(n_565), .D(n_578), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B1(n_547), .B2(n_549), .C(n_550), .Y(n_544) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_559), .Y(n_553) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NOR2x1_ASAP7_75t_L g565 ( .A(n_566), .B(n_571), .Y(n_565) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_575), .B2(n_576), .Y(n_571) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_577), .Y(n_729) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
INVx2_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_581), .A2(n_691), .B1(n_692), .B2(n_693), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_632), .B1(n_633), .B2(n_677), .Y(n_588) );
INVx1_ASAP7_75t_L g677 ( .A(n_589), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_606), .B2(n_631), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
XNOR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_605), .Y(n_592) );
NOR2x1_ASAP7_75t_L g593 ( .A(n_594), .B(n_599), .Y(n_593) );
NAND4xp25_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .C(n_597), .D(n_598), .Y(n_594) );
NAND4xp25_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .C(n_603), .D(n_604), .Y(n_599) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g631 ( .A(n_609), .Y(n_631) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g630 ( .A(n_611), .Y(n_630) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_618), .Y(n_611) );
NAND4xp25_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .C(n_615), .D(n_617), .Y(n_612) );
BUFx6f_ASAP7_75t_SL g731 ( .A(n_616), .Y(n_731) );
NAND4xp25_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .C(n_625), .D(n_626), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
XNOR2x1_ASAP7_75t_L g635 ( .A(n_636), .B(n_659), .Y(n_635) );
INVx2_ASAP7_75t_L g658 ( .A(n_638), .Y(n_658) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_649), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .C(n_645), .D(n_647), .Y(n_639) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g721 ( .A(n_644), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .C(n_653), .D(n_656), .Y(n_649) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_662), .B(n_670), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_667), .Y(n_662) );
OAI21xp5_ASAP7_75t_SL g663 ( .A1(n_664), .A2(n_665), .B(n_666), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_674), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_737), .B2(n_775), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
AO22x2_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_708), .B1(n_733), .B2(n_736), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g735 ( .A(n_683), .Y(n_735) );
INVx1_ASAP7_75t_L g707 ( .A(n_685), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_699), .Y(n_685) );
NOR3xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_690), .C(n_694), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_688), .B(n_689), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_703), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVx2_ASAP7_75t_L g736 ( .A(n_708), .Y(n_736) );
NAND4xp75_ASAP7_75t_L g709 ( .A(n_710), .B(n_716), .C(n_724), .D(n_730), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .Y(n_710) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_722), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_728), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g775 ( .A(n_737), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B1(n_755), .B2(n_756), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_749), .Y(n_741) );
NAND4xp25_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .C(n_746), .D(n_747), .Y(n_742) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .C(n_752), .D(n_753), .Y(n_749) );
INVx5_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NOR2x1_ASAP7_75t_L g757 ( .A(n_758), .B(n_768), .Y(n_757) );
NAND4xp25_ASAP7_75t_L g758 ( .A(n_759), .B(n_762), .C(n_764), .D(n_767), .Y(n_758) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND4xp25_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .C(n_773), .D(n_774), .Y(n_768) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_780), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_778), .B(n_781), .Y(n_827) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
OAI222xp33_ASAP7_75t_R g786 ( .A1(n_787), .A2(n_804), .B1(n_808), .B2(n_824), .C1(n_825), .C2(n_828), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NAND2x1_ASAP7_75t_SL g790 ( .A(n_791), .B(n_796), .Y(n_790) );
NOR2xp67_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
NOR2x1_ASAP7_75t_L g796 ( .A(n_797), .B(n_800), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx2_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
NOR2x1_ASAP7_75t_L g810 ( .A(n_811), .B(n_817), .Y(n_810) );
NAND4xp25_ASAP7_75t_SL g811 ( .A(n_812), .B(n_813), .C(n_814), .D(n_816), .Y(n_811) );
NAND4xp25_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .C(n_822), .D(n_823), .Y(n_817) );
INVx1_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
CKINVDCx6p67_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
endmodule