module fake_jpeg_29414_n_457 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_457);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_457;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_15),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_48),
.B(n_92),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_63),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_60),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_62),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_15),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_67),
.Y(n_101)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_41),
.Y(n_72)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g105 ( 
.A(n_74),
.Y(n_105)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_29),
.B(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_43),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_29),
.B(n_0),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_24),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_99),
.B(n_103),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_51),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_51),
.A2(n_24),
.B(n_40),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_108),
.B(n_38),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_62),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_111),
.B(n_116),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_28),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_133),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_47),
.B(n_28),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_52),
.B(n_25),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_54),
.B(n_25),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_44),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_83),
.B(n_44),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_150),
.Y(n_193)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_94),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_153),
.B(n_161),
.Y(n_216)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_108),
.A2(n_53),
.B1(n_75),
.B2(n_86),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_124),
.B1(n_70),
.B2(n_123),
.Y(n_206)
);

CKINVDCx11_ASAP7_75t_R g159 ( 
.A(n_109),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_170),
.Y(n_204)
);

CKINVDCx12_ASAP7_75t_R g160 ( 
.A(n_109),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_97),
.A2(n_92),
.B1(n_90),
.B2(n_49),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_162),
.A2(n_169),
.B1(n_177),
.B2(n_98),
.Y(n_227)
);

CKINVDCx9p33_ASAP7_75t_R g163 ( 
.A(n_109),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_167),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_21),
.B1(n_57),
.B2(n_65),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_104),
.A2(n_36),
.B1(n_33),
.B2(n_40),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_42),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_189),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_121),
.A2(n_68),
.B1(n_80),
.B2(n_56),
.Y(n_169)
);

CKINVDCx12_ASAP7_75t_R g170 ( 
.A(n_122),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_SL g172 ( 
.A(n_101),
.B(n_35),
.C(n_23),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_178),
.Y(n_209)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

CKINVDCx9p33_ASAP7_75t_R g176 ( 
.A(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_61),
.B1(n_69),
.B2(n_71),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_180),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_129),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_186),
.Y(n_220)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_183),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_100),
.B(n_81),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_164),
.CI(n_162),
.CON(n_207),
.SN(n_207)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_138),
.A2(n_74),
.B1(n_125),
.B2(n_42),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_113),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_102),
.A2(n_107),
.B1(n_142),
.B2(n_96),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_142),
.B1(n_96),
.B2(n_137),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g191 ( 
.A(n_112),
.B(n_23),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_191),
.B(n_35),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_198),
.A2(n_208),
.B1(n_217),
.B2(n_163),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_125),
.B(n_120),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_136),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_210),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_207),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_136),
.B1(n_98),
.B2(n_130),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_130),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_147),
.A2(n_113),
.B1(n_36),
.B2(n_20),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_184),
.A2(n_118),
.B1(n_127),
.B2(n_95),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_34),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_148),
.B(n_105),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_221),
.B(n_38),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_173),
.A2(n_20),
.B1(n_34),
.B2(n_105),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_227),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_167),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_228),
.B(n_31),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_240),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_156),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_230),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_191),
.B1(n_177),
.B2(n_169),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_232),
.A2(n_243),
.B1(n_227),
.B2(n_188),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_157),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_237),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_187),
.B1(n_176),
.B2(n_123),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_236),
.A2(n_212),
.B1(n_199),
.B2(n_222),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_171),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_238),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_239),
.B(n_247),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_186),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_152),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_245),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_242),
.A2(n_258),
.B1(n_199),
.B2(n_193),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_127),
.B1(n_118),
.B2(n_182),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_155),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_189),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_179),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_251),
.Y(n_274)
);

AND2x6_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_105),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_257),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_175),
.Y(n_253)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_254),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_220),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_260),
.Y(n_290)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_206),
.A2(n_149),
.B1(n_74),
.B2(n_77),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_203),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_201),
.B(n_151),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_262),
.A2(n_275),
.B(n_283),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_200),
.C(n_215),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_265),
.C(n_271),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_213),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_264),
.B(n_272),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_195),
.C(n_220),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_234),
.C(n_231),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_225),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_204),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_273),
.B(n_228),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_246),
.A2(n_197),
.B(n_217),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_279),
.A2(n_243),
.B1(n_227),
.B2(n_238),
.Y(n_309)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_241),
.B(n_239),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_282),
.B(n_287),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_246),
.A2(n_208),
.B(n_193),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_228),
.B(n_244),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_255),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_233),
.B1(n_242),
.B2(n_258),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_229),
.B(n_194),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_194),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_245),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_292),
.B(n_300),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_233),
.B1(n_232),
.B2(n_246),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_293),
.A2(n_227),
.B1(n_276),
.B2(n_291),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_266),
.B(n_251),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_294),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_260),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_295),
.B(n_263),
.C(n_265),
.Y(n_333)
);

OR2x4_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_249),
.Y(n_297)
);

OAI31xp33_ASAP7_75t_L g342 ( 
.A1(n_297),
.A2(n_250),
.A3(n_254),
.B(n_214),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_237),
.Y(n_299)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_278),
.Y(n_302)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_303),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_304),
.A2(n_318),
.B(n_319),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_306),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_267),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_270),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_267),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_311),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_290),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_268),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_266),
.B(n_252),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_274),
.B(n_252),
.Y(n_315)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_315),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_261),
.A2(n_256),
.B1(n_259),
.B2(n_196),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_316),
.A2(n_310),
.B(n_278),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_196),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_259),
.B(n_203),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_284),
.A2(n_268),
.B(n_274),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_321),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_323),
.B(n_304),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_284),
.B(n_288),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_324),
.A2(n_332),
.B(n_348),
.Y(n_350)
);

OA21x2_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_269),
.B(n_279),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_328),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_318),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_330),
.A2(n_338),
.B1(n_313),
.B2(n_306),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_320),
.A2(n_290),
.B(n_291),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_336),
.C(n_341),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_273),
.C(n_270),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_307),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_124),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_301),
.B(n_276),
.C(n_224),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_342),
.A2(n_319),
.B(n_296),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_343),
.A2(n_131),
.B(n_110),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_281),
.Y(n_344)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_344),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_310),
.A2(n_277),
.B(n_150),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_347),
.A2(n_349),
.B1(n_340),
.B2(n_300),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_351),
.A2(n_353),
.B1(n_358),
.B2(n_361),
.Y(n_374)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_344),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_369),
.Y(n_375)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_335),
.Y(n_357)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_357),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_349),
.A2(n_308),
.B1(n_311),
.B2(n_296),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_324),
.A2(n_293),
.B1(n_309),
.B2(n_312),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_359),
.A2(n_368),
.B1(n_370),
.B2(n_342),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_303),
.C(n_299),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_363),
.C(n_365),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_347),
.A2(n_298),
.B1(n_294),
.B2(n_292),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_362),
.B(n_334),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_297),
.C(n_277),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_224),
.C(n_214),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_322),
.A2(n_302),
.B1(n_256),
.B2(n_43),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_367),
.A2(n_372),
.B1(n_348),
.B2(n_329),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_328),
.A2(n_302),
.B1(n_254),
.B2(n_250),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_331),
.B(n_183),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_345),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_325),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_322),
.A2(n_330),
.B1(n_346),
.B2(n_326),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_346),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_339),
.C(n_323),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_379),
.C(n_386),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_378),
.A2(n_350),
.B1(n_370),
.B2(n_368),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_334),
.C(n_332),
.Y(n_379)
);

NOR2x1_ASAP7_75t_SL g381 ( 
.A(n_357),
.B(n_327),
.Y(n_381)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_381),
.Y(n_393)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_387),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_384),
.B(n_385),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_326),
.C(n_343),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_325),
.C(n_345),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_388),
.B(n_362),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_372),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_329),
.C(n_327),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_392),
.C(n_350),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_391),
.A2(n_367),
.B1(n_39),
.B2(n_131),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_327),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_380),
.A2(n_352),
.B(n_364),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_394),
.A2(n_385),
.B(n_376),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_396),
.B(n_397),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_353),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_399),
.B(n_404),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_359),
.Y(n_400)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_400),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_401),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_418)
);

XNOR2x1_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_43),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_379),
.B(n_366),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_405),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_376),
.B(n_364),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_29),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_384),
.A2(n_392),
.B(n_390),
.C(n_386),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_407),
.A2(n_377),
.B(n_3),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_408),
.A2(n_39),
.B1(n_73),
.B2(n_50),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_402),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_409),
.Y(n_425)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_411),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_414),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_415),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_110),
.C(n_31),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_416),
.B(n_419),
.C(n_31),
.Y(n_433)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_417),
.A2(n_403),
.B(n_405),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_418),
.A2(n_408),
.B1(n_410),
.B2(n_421),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_31),
.C(n_29),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_394),
.B(n_1),
.Y(n_422)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_422),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_412),
.B(n_395),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_427),
.Y(n_441)
);

AOI21x1_ASAP7_75t_L g428 ( 
.A1(n_420),
.A2(n_407),
.B(n_395),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_428),
.A2(n_431),
.B(n_415),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_430),
.A2(n_433),
.B1(n_427),
.B2(n_429),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_409),
.A2(n_1),
.B(n_6),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_31),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_432),
.B(n_433),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_416),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_440),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_434),
.B(n_411),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_438),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_414),
.C(n_419),
.Y(n_438)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_439),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_441),
.B(n_429),
.C(n_428),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_443),
.B(n_430),
.Y(n_450)
);

INVx11_ASAP7_75t_L g446 ( 
.A(n_442),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_446),
.A2(n_435),
.B(n_436),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_444),
.Y(n_448)
);

AOI322xp5_ASAP7_75t_L g451 ( 
.A1(n_448),
.A2(n_449),
.A3(n_450),
.B1(n_446),
.B2(n_447),
.C1(n_444),
.C2(n_443),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_451),
.B(n_452),
.C(n_7),
.Y(n_453)
);

AOI322xp5_ASAP7_75t_L g452 ( 
.A1(n_450),
.A2(n_445),
.A3(n_7),
.B1(n_9),
.B2(n_10),
.C1(n_12),
.C2(n_6),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_453),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_454),
.A2(n_7),
.B(n_9),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_455),
.A2(n_7),
.B(n_10),
.Y(n_456)
);

FAx1_ASAP7_75t_SL g457 ( 
.A(n_456),
.B(n_12),
.CI(n_453),
.CON(n_457),
.SN(n_457)
);


endmodule