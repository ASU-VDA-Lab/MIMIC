module real_jpeg_10278_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_302, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_302;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_286;
wire n_215;
wire n_166;
wire n_300;
wire n_176;
wire n_221;
wire n_249;
wire n_292;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_295;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_181;
wire n_85;
wire n_102;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx24_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_1),
.A2(n_52),
.B1(n_64),
.B2(n_67),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_2),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_2),
.A2(n_11),
.B(n_33),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_27),
.B1(n_35),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_3),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_95),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_3),
.A2(n_64),
.B1(n_67),
.B2(n_95),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_4),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_4),
.A2(n_36),
.B1(n_64),
.B2(n_67),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_4),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_10),
.A2(n_27),
.B1(n_35),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_10),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_64),
.B1(n_67),
.B2(n_116),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_116),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_116),
.Y(n_236)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_11),
.A2(n_49),
.B(n_59),
.C(n_130),
.D(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_11),
.B(n_49),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_11),
.B(n_47),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_11),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_11),
.A2(n_84),
.B(n_149),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_11),
.A2(n_32),
.B(n_43),
.C(n_180),
.D(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_11),
.B(n_32),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_11),
.B(n_118),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_11),
.A2(n_27),
.B1(n_35),
.B2(n_162),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_13),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_13),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_13),
.A2(n_38),
.B1(n_64),
.B2(n_67),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_55),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_14),
.A2(n_55),
.B1(n_64),
.B2(n_67),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_15),
.A2(n_48),
.B1(n_49),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_15),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_15),
.A2(n_64),
.B1(n_67),
.B2(n_70),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_16),
.A2(n_48),
.B1(n_49),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_16),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_16),
.A2(n_64),
.B1(n_67),
.B2(n_144),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_144),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_16),
.A2(n_27),
.B1(n_35),
.B2(n_144),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_119),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_97),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_20),
.B(n_97),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_72),
.B2(n_73),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_25)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_26),
.A2(n_115),
.B(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_26),
.A2(n_31),
.B1(n_115),
.B2(n_248),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_29),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_27),
.A2(n_29),
.B(n_162),
.C(n_222),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_31),
.A2(n_34),
.B(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_31),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_31),
.A2(n_93),
.B(n_248),
.Y(n_247)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_44),
.B(n_46),
.C(n_47),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_44),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_56),
.B1(n_57),
.B2(n_71),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_42),
.A2(n_53),
.B1(n_200),
.B2(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_42),
.A2(n_236),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_47),
.B1(n_51),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_43),
.A2(n_47),
.B1(n_75),
.B2(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_43),
.B(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_44),
.B(n_49),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_46),
.A2(n_48),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_60),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_53),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_53),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_53),
.A2(n_201),
.B(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_68),
.B(n_69),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_68),
.B1(n_78),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_58),
.A2(n_68),
.B1(n_90),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_58),
.A2(n_68),
.B1(n_143),
.B2(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_58),
.A2(n_178),
.B(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_58),
.A2(n_68),
.B1(n_110),
.B2(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_63),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_59),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_67),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_60),
.B(n_67),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_62),
.A2(n_64),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_67),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_68),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_68),
.A2(n_143),
.B(n_145),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_68),
.B(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_68),
.A2(n_145),
.B(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_74),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_91),
.B(n_92),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_82),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_91),
.B1(n_92),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_83),
.A2(n_89),
.B1(n_91),
.B2(n_283),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B(n_88),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_87),
.B1(n_88),
.B2(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_84),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_84),
.A2(n_87),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_84),
.A2(n_87),
.B1(n_108),
.B2(n_226),
.Y(n_255)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_85),
.A2(n_86),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_85),
.B(n_150),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_85),
.A2(n_86),
.B1(n_191),
.B2(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_86),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_87),
.A2(n_155),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_87),
.B(n_162),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_87),
.A2(n_164),
.B(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_89),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_96),
.A2(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.C(n_104),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_98),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_104),
.A2(n_105),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.C(n_113),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_106),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_107),
.B(n_109),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_111),
.A2(n_113),
.B1(n_114),
.B2(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_111),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_112),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_117),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI321xp33_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_276),
.A3(n_289),
.B1(n_295),
.B2(n_300),
.C(n_302),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_242),
.C(n_272),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_215),
.B(n_241),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_194),
.B(n_214),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_172),
.B(n_193),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_151),
.B(n_171),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_137),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_128),
.B(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_133),
.B1(n_134),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_131),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_147),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_142),
.C(n_147),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_148),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_159),
.B(n_170),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_153),
.B(n_157),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_165),
.B(n_169),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_163),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_173),
.B(n_174),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_185),
.B2(n_192),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_179),
.B1(n_183),
.B2(n_184),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_184),
.C(n_192),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_181),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_189),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_196),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_208),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_210),
.C(n_212),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_203),
.B2(n_207),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_204),
.C(n_205),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_203),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_209),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_210),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_216),
.B(n_217),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_230),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_219),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_229),
.C(n_230),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_224),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_227),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_238),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_234),
.B1(n_235),
.B2(n_237),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_232),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_243),
.A2(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_258),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_244),
.B(n_258),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_254),
.C(n_257),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_249),
.B1(n_250),
.B2(n_252),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_247),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_252),
.C(n_253),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_257),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_256),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_270),
.B2(n_271),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_262),
.C(n_271),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_267),
.C(n_269),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_265),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_274),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_285),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_285),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_282),
.C(n_284),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_278),
.A2(n_279),
.B1(n_282),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_282),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_296),
.B(n_299),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);


endmodule