module fake_aes_7818_n_830 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_830);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_830;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_384;
wire n_434;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_86;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_SL g85 ( .A(n_62), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_61), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_67), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_64), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_5), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_11), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_58), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_14), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_41), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_46), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_56), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_74), .Y(n_96) );
BUFx8_ASAP7_75t_SL g97 ( .A(n_63), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_51), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_80), .Y(n_99) );
BUFx10_ASAP7_75t_L g100 ( .A(n_65), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_59), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_36), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_5), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_38), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_76), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_18), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_23), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_33), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_15), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_57), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_20), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_73), .Y(n_112) );
INVx4_ASAP7_75t_R g113 ( .A(n_68), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_39), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_19), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_49), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_40), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_3), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_60), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_17), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_36), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_18), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_14), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_6), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_30), .Y(n_125) );
AND2x6_ASAP7_75t_L g126 ( .A(n_118), .B(n_45), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_92), .B(n_0), .Y(n_127) );
BUFx12f_ASAP7_75t_L g128 ( .A(n_100), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_85), .B(n_0), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_92), .B(n_1), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_115), .B(n_1), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
BUFx12f_ASAP7_75t_L g133 ( .A(n_100), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_115), .B(n_2), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
INVx5_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_90), .B(n_2), .Y(n_137) );
BUFx12f_ASAP7_75t_L g138 ( .A(n_100), .Y(n_138) );
NOR2xp33_ASAP7_75t_SL g139 ( .A(n_98), .B(n_47), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_115), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_90), .B(n_3), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_87), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_87), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_85), .B(n_4), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_102), .B(n_4), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_122), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
INVx5_ASAP7_75t_L g148 ( .A(n_100), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_129), .A2(n_103), .B1(n_99), .B2(n_123), .Y(n_149) );
NAND2xp33_ASAP7_75t_SL g150 ( .A(n_127), .B(n_99), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_132), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_129), .A2(n_103), .B1(n_124), .B2(n_107), .Y(n_152) );
OAI22xp33_ASAP7_75t_SL g153 ( .A1(n_139), .A2(n_125), .B1(n_89), .B2(n_120), .Y(n_153) );
INVxp33_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
AO22x2_ASAP7_75t_L g155 ( .A1(n_129), .A2(n_121), .B1(n_109), .B2(n_104), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_129), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_148), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_129), .A2(n_108), .B1(n_114), .B2(n_93), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_148), .B(n_100), .Y(n_159) );
INVxp67_ASAP7_75t_SL g160 ( .A(n_140), .Y(n_160) );
OAI22xp33_ASAP7_75t_L g161 ( .A1(n_137), .A2(n_109), .B1(n_121), .B2(n_102), .Y(n_161) );
OA22x2_ASAP7_75t_L g162 ( .A1(n_127), .A2(n_104), .B1(n_118), .B2(n_111), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_148), .B(n_118), .Y(n_163) );
OAI22xp33_ASAP7_75t_L g164 ( .A1(n_137), .A2(n_106), .B1(n_117), .B2(n_122), .Y(n_164) );
AO22x2_ASAP7_75t_L g165 ( .A1(n_129), .A2(n_91), .B1(n_94), .B2(n_119), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_129), .A2(n_98), .B1(n_122), .B2(n_105), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_148), .B(n_122), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_129), .A2(n_122), .B1(n_119), .B2(n_91), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_148), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_144), .A2(n_122), .B1(n_94), .B2(n_116), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_140), .B(n_101), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_128), .Y(n_172) );
OAI22xp33_ASAP7_75t_SL g173 ( .A1(n_139), .A2(n_116), .B1(n_105), .B2(n_101), .Y(n_173) );
OAI22xp33_ASAP7_75t_SL g174 ( .A1(n_139), .A2(n_88), .B1(n_95), .B2(n_96), .Y(n_174) );
NAND2xp33_ASAP7_75t_SL g175 ( .A(n_127), .B(n_122), .Y(n_175) );
INVx8_ASAP7_75t_L g176 ( .A(n_128), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_148), .B(n_110), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_144), .A2(n_112), .B1(n_113), .B2(n_97), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_140), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_148), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_144), .A2(n_113), .B1(n_97), .B2(n_8), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_131), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_137), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_183) );
NAND3x1_ASAP7_75t_L g184 ( .A(n_127), .B(n_7), .C(n_9), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_144), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g186 ( .A1(n_141), .A2(n_10), .B1(n_12), .B2(n_13), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_144), .A2(n_12), .B1(n_13), .B2(n_15), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_148), .B(n_16), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_131), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_148), .B(n_135), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_148), .B(n_16), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_144), .A2(n_17), .B1(n_19), .B2(n_20), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_144), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
BUFx6f_ASAP7_75t_SL g196 ( .A(n_176), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_156), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_191), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_154), .B(n_130), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_191), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
NOR2xp33_ASAP7_75t_SL g203 ( .A(n_176), .B(n_128), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_160), .B(n_130), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_179), .B(n_128), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_155), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_168), .A2(n_147), .B(n_135), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_160), .B(n_130), .Y(n_208) );
XOR2x2_ASAP7_75t_L g209 ( .A(n_149), .B(n_130), .Y(n_209) );
NAND2x1p5_ASAP7_75t_L g210 ( .A(n_185), .B(n_148), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_155), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_165), .B(n_130), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_188), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_150), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_163), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_171), .B(n_148), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_182), .B(n_128), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_176), .Y(n_220) );
BUFx6f_ASAP7_75t_SL g221 ( .A(n_157), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_190), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_167), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_159), .Y(n_224) );
XNOR2xp5_ASAP7_75t_L g225 ( .A(n_181), .B(n_131), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_171), .B(n_148), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_170), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_187), .Y(n_228) );
OR2x2_ASAP7_75t_SL g229 ( .A(n_184), .B(n_141), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_178), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_193), .Y(n_231) );
INVxp67_ASAP7_75t_SL g232 ( .A(n_169), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_152), .B(n_131), .Y(n_233) );
NOR2xp67_ASAP7_75t_L g234 ( .A(n_166), .B(n_133), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_194), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_158), .B(n_133), .Y(n_236) );
XOR2xp5_ASAP7_75t_SL g237 ( .A(n_189), .B(n_131), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_177), .B(n_133), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_172), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_157), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_180), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_192), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_175), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_162), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_162), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_183), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_153), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_183), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_164), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_161), .B(n_134), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_186), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_186), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_173), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_161), .Y(n_254) );
AND2x2_ASAP7_75t_SL g255 ( .A(n_174), .B(n_134), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_199), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_213), .B(n_133), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_213), .B(n_138), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_208), .B(n_138), .Y(n_259) );
INVxp67_ASAP7_75t_SL g260 ( .A(n_212), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_208), .B(n_138), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_199), .Y(n_262) );
NOR2xp67_ASAP7_75t_R g263 ( .A(n_217), .B(n_135), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_196), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_204), .B(n_138), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_204), .B(n_164), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_201), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_204), .B(n_138), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_204), .B(n_134), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_250), .B(n_134), .Y(n_270) );
AND2x2_ASAP7_75t_SL g271 ( .A(n_217), .B(n_134), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_201), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_250), .B(n_135), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_233), .B(n_147), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_221), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_220), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_233), .B(n_147), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_255), .B(n_141), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_255), .B(n_145), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_197), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_197), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_202), .B(n_136), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_220), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_196), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_198), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_202), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_198), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_233), .B(n_147), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_240), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_221), .Y(n_290) );
AND2x2_ASAP7_75t_SL g291 ( .A(n_206), .B(n_132), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_240), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_206), .B(n_136), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_211), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_221), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_211), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_196), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_196), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_233), .B(n_136), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_222), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_195), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_228), .B(n_136), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_228), .B(n_231), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_231), .B(n_136), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_221), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_214), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_256), .B(n_262), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_256), .B(n_222), .Y(n_308) );
NOR2x1_ASAP7_75t_SL g309 ( .A(n_256), .B(n_237), .Y(n_309) );
CKINVDCx8_ASAP7_75t_R g310 ( .A(n_267), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_256), .B(n_235), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_256), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_257), .B(n_235), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_267), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_267), .Y(n_315) );
AND2x2_ASAP7_75t_SL g316 ( .A(n_291), .B(n_203), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_267), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_267), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_256), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_262), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_262), .B(n_254), .Y(n_321) );
OR2x6_ASAP7_75t_L g322 ( .A(n_262), .B(n_210), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_267), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_277), .B(n_209), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_262), .Y(n_325) );
AND2x6_ASAP7_75t_L g326 ( .A(n_262), .B(n_246), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_267), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_277), .B(n_209), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_272), .B(n_254), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_257), .B(n_225), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_272), .Y(n_331) );
OR2x6_ASAP7_75t_L g332 ( .A(n_272), .B(n_210), .Y(n_332) );
BUFx4f_ASAP7_75t_L g333 ( .A(n_275), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_275), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_277), .B(n_237), .Y(n_335) );
NOR2x1_ASAP7_75t_L g336 ( .A(n_275), .B(n_253), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_272), .B(n_216), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_272), .B(n_200), .Y(n_338) );
BUFx12f_ASAP7_75t_L g339 ( .A(n_331), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_312), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_331), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_317), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_307), .B(n_272), .Y(n_344) );
BUFx4f_ASAP7_75t_SL g345 ( .A(n_307), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
INVx1_ASAP7_75t_SL g347 ( .A(n_307), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_326), .Y(n_348) );
CKINVDCx11_ASAP7_75t_R g349 ( .A(n_310), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_312), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_319), .B(n_286), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_313), .A2(n_251), .B1(n_246), .B2(n_248), .Y(n_352) );
BUFx2_ASAP7_75t_SL g353 ( .A(n_319), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_320), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g355 ( .A(n_319), .B(n_286), .Y(n_355) );
BUFx2_ASAP7_75t_SL g356 ( .A(n_310), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_317), .Y(n_358) );
CKINVDCx6p67_ASAP7_75t_R g359 ( .A(n_326), .Y(n_359) );
INVx5_ASAP7_75t_L g360 ( .A(n_322), .Y(n_360) );
BUFx12f_ASAP7_75t_L g361 ( .A(n_326), .Y(n_361) );
INVx4_ASAP7_75t_L g362 ( .A(n_322), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_317), .Y(n_363) );
INVx2_ASAP7_75t_SL g364 ( .A(n_317), .Y(n_364) );
CKINVDCx16_ASAP7_75t_R g365 ( .A(n_322), .Y(n_365) );
INVx8_ASAP7_75t_L g366 ( .A(n_326), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_317), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_354), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_354), .B(n_303), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_352), .B(n_303), .Y(n_371) );
INVx4_ASAP7_75t_L g372 ( .A(n_339), .Y(n_372) );
OAI21xp5_ASAP7_75t_SL g373 ( .A1(n_348), .A2(n_264), .B(n_284), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_340), .Y(n_375) );
BUFx2_ASAP7_75t_SL g376 ( .A(n_360), .Y(n_376) );
BUFx2_ASAP7_75t_R g377 ( .A(n_356), .Y(n_377) );
BUFx10_ASAP7_75t_L g378 ( .A(n_350), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_352), .B(n_303), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_345), .Y(n_380) );
INVx6_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
INVx8_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_350), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_350), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_345), .A2(n_316), .B1(n_332), .B2(n_322), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g386 ( .A1(n_348), .A2(n_264), .B(n_284), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_339), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_343), .B(n_303), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
BUFx8_ASAP7_75t_L g390 ( .A(n_339), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_345), .A2(n_316), .B1(n_332), .B2(n_322), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_341), .A2(n_313), .B1(n_330), .B2(n_324), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_365), .A2(n_335), .B1(n_324), .B2(n_328), .Y(n_393) );
INVx6_ASAP7_75t_L g394 ( .A(n_343), .Y(n_394) );
OAI22xp5_ASAP7_75t_SL g395 ( .A1(n_365), .A2(n_229), .B1(n_215), .B2(n_247), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_349), .Y(n_396) );
CKINVDCx6p67_ASAP7_75t_R g397 ( .A(n_349), .Y(n_397) );
BUFx2_ASAP7_75t_SL g398 ( .A(n_360), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_352), .B(n_303), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_343), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_361), .A2(n_309), .B1(n_316), .B2(n_326), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_343), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_365), .A2(n_332), .B1(n_311), .B2(n_260), .Y(n_403) );
BUFx12f_ASAP7_75t_L g404 ( .A(n_361), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_344), .Y(n_405) );
INVx6_ASAP7_75t_L g406 ( .A(n_343), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_359), .A2(n_332), .B1(n_229), .B2(n_325), .Y(n_407) );
CKINVDCx6p67_ASAP7_75t_R g408 ( .A(n_360), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_341), .A2(n_326), .B1(n_337), .B2(n_308), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_341), .A2(n_361), .B1(n_326), .B2(n_337), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_393), .A2(n_361), .B1(n_362), .B2(n_348), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_368), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g413 ( .A1(n_369), .A2(n_361), .B1(n_366), .B2(n_309), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_388), .B(n_347), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_369), .B(n_344), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_374), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_407), .A2(n_362), .B1(n_348), .B2(n_366), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_375), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_383), .B(n_347), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_400), .B(n_362), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_409), .A2(n_359), .B1(n_360), .B2(n_366), .Y(n_422) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_382), .A2(n_366), .B1(n_360), .B2(n_362), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_382), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_384), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_372), .A2(n_359), .B1(n_360), .B2(n_366), .Y(n_426) );
OAI21xp5_ASAP7_75t_SL g427 ( .A1(n_401), .A2(n_264), .B(n_284), .Y(n_427) );
OAI222xp33_ASAP7_75t_L g428 ( .A1(n_372), .A2(n_362), .B1(n_360), .B2(n_347), .C1(n_332), .C2(n_346), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_395), .A2(n_362), .B1(n_366), .B2(n_360), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_370), .B(n_230), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_408), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g432 ( .A1(n_371), .A2(n_311), .B(n_251), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_392), .A2(n_362), .B1(n_366), .B2(n_360), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_378), .Y(n_434) );
OAI21xp33_ASAP7_75t_L g435 ( .A1(n_409), .A2(n_325), .B(n_320), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_392), .A2(n_366), .B1(n_360), .B2(n_359), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_378), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_379), .A2(n_366), .B1(n_360), .B2(n_252), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_399), .A2(n_326), .B1(n_308), .B2(n_249), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_382), .A2(n_366), .B1(n_360), .B2(n_248), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_389), .B(n_337), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_405), .B(n_342), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_385), .A2(n_353), .B1(n_356), .B2(n_260), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_378), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_376), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_396), .B(n_239), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_396), .B(n_225), .Y(n_447) );
BUFx12f_ASAP7_75t_L g448 ( .A(n_390), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_381), .A2(n_356), .B1(n_353), .B2(n_346), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_400), .B(n_342), .Y(n_450) );
AOI22xp33_ASAP7_75t_SL g451 ( .A1(n_381), .A2(n_353), .B1(n_346), .B2(n_274), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_390), .A2(n_252), .B1(n_255), .B2(n_308), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_402), .B(n_342), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_398), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_408), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_390), .A2(n_279), .B1(n_278), .B2(n_271), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_402), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_397), .A2(n_279), .B1(n_278), .B2(n_271), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_410), .B(n_342), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_397), .B(n_244), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_391), .A2(n_353), .B1(n_260), .B2(n_321), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_403), .A2(n_338), .B1(n_279), .B2(n_278), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_372), .A2(n_271), .B1(n_338), .B2(n_210), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_381), .A2(n_346), .B1(n_333), .B2(n_297), .Y(n_464) );
AOI22xp5_ASAP7_75t_SL g465 ( .A1(n_387), .A2(n_346), .B1(n_297), .B2(n_298), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_410), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_394), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_404), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_394), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_373), .A2(n_271), .B1(n_274), .B2(n_288), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_394), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_406), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_406), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_406), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_380), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_377), .A2(n_329), .B1(n_321), .B2(n_271), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_386), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_409), .A2(n_329), .B1(n_271), .B2(n_346), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_408), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_393), .A2(n_336), .B1(n_291), .B2(n_346), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_388), .B(n_342), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_415), .B(n_244), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_412), .B(n_245), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_412), .B(n_245), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_470), .A2(n_300), .B1(n_274), .B2(n_288), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_478), .A2(n_126), .B1(n_291), .B2(n_300), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_460), .B(n_145), .C(n_142), .Y(n_487) );
OAI211xp5_ASAP7_75t_SL g488 ( .A1(n_447), .A2(n_145), .B(n_253), .C(n_273), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_476), .A2(n_126), .B1(n_291), .B2(n_300), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_425), .B(n_274), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_459), .B(n_367), .Y(n_491) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_435), .A2(n_364), .B(n_318), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_476), .A2(n_126), .B1(n_288), .B2(n_274), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_470), .A2(n_351), .B1(n_355), .B2(n_273), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_477), .A2(n_126), .B1(n_288), .B2(n_266), .Y(n_495) );
OAI221xp5_ASAP7_75t_SL g496 ( .A1(n_477), .A2(n_427), .B1(n_439), .B2(n_458), .C(n_452), .Y(n_496) );
OAI211xp5_ASAP7_75t_L g497 ( .A1(n_427), .A2(n_298), .B(n_297), .C(n_266), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_466), .A2(n_126), .B1(n_288), .B2(n_266), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_466), .A2(n_126), .B1(n_333), .B2(n_270), .Y(n_499) );
AOI22xp33_ASAP7_75t_SL g500 ( .A1(n_431), .A2(n_357), .B1(n_363), .B2(n_298), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_422), .A2(n_126), .B1(n_333), .B2(n_270), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_465), .B(n_142), .C(n_146), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_425), .B(n_367), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_439), .A2(n_351), .B1(n_355), .B2(n_364), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_429), .A2(n_351), .B1(n_355), .B2(n_364), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_433), .A2(n_126), .B1(n_294), .B2(n_299), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_411), .A2(n_126), .B1(n_294), .B2(n_299), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_459), .B(n_367), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_479), .A2(n_357), .B1(n_363), .B2(n_367), .Y(n_509) );
OAI222xp33_ASAP7_75t_L g510 ( .A1(n_465), .A2(n_364), .B1(n_334), .B2(n_351), .C1(n_355), .C2(n_367), .Y(n_510) );
OAI222xp33_ASAP7_75t_L g511 ( .A1(n_424), .A2(n_334), .B1(n_351), .B2(n_355), .C1(n_367), .C2(n_363), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_456), .A2(n_126), .B1(n_299), .B2(n_357), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_434), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_462), .A2(n_351), .B1(n_355), .B2(n_273), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_416), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_420), .B(n_126), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_420), .B(n_126), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_448), .A2(n_363), .B1(n_357), .B2(n_334), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_416), .B(n_358), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_461), .A2(n_299), .B1(n_267), .B2(n_304), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_416), .B(n_358), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_448), .A2(n_334), .B1(n_358), .B2(n_258), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_463), .A2(n_267), .B1(n_302), .B2(n_304), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_480), .A2(n_267), .B1(n_302), .B2(n_304), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_443), .A2(n_267), .B1(n_302), .B2(n_304), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_443), .A2(n_267), .B1(n_302), .B2(n_304), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_436), .A2(n_302), .B1(n_236), .B2(n_257), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_462), .A2(n_358), .B1(n_306), .B2(n_327), .Y(n_528) );
INVxp33_ASAP7_75t_L g529 ( .A(n_446), .Y(n_529) );
AOI222xp33_ASAP7_75t_L g530 ( .A1(n_448), .A2(n_269), .B1(n_257), .B2(n_258), .C1(n_259), .C2(n_261), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_423), .A2(n_358), .B1(n_306), .B2(n_327), .Y(n_531) );
INVx4_ASAP7_75t_L g532 ( .A(n_418), .Y(n_532) );
NOR3xp33_ASAP7_75t_SL g533 ( .A(n_430), .B(n_243), .C(n_219), .Y(n_533) );
OAI22xp33_ASAP7_75t_L g534 ( .A1(n_418), .A2(n_358), .B1(n_327), .B2(n_283), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_438), .A2(n_258), .B1(n_257), .B2(n_358), .Y(n_535) );
AO22x1_ASAP7_75t_L g536 ( .A1(n_418), .A2(n_358), .B1(n_295), .B2(n_275), .Y(n_536) );
OAI21xp33_ASAP7_75t_L g537 ( .A1(n_435), .A2(n_132), .B(n_143), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_432), .A2(n_258), .B1(n_358), .B2(n_280), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_417), .A2(n_287), .B1(n_280), .B2(n_234), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_455), .A2(n_287), .B1(n_280), .B2(n_234), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_455), .A2(n_280), .B1(n_287), .B2(n_281), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_445), .A2(n_280), .B1(n_287), .B2(n_281), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_445), .A2(n_454), .B1(n_451), .B2(n_414), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_454), .A2(n_287), .B1(n_285), .B2(n_281), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_414), .A2(n_287), .B1(n_285), .B2(n_281), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_419), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_424), .A2(n_261), .B1(n_259), .B2(n_306), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_434), .B(n_142), .C(n_146), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_419), .B(n_142), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_421), .A2(n_285), .B1(n_269), .B2(n_327), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_413), .A2(n_327), .B1(n_283), .B2(n_276), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_419), .B(n_21), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_421), .A2(n_269), .B1(n_323), .B2(n_315), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_440), .A2(n_306), .B1(n_318), .B2(n_296), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_481), .B(n_22), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_457), .B(n_146), .Y(n_556) );
OAI22xp33_ASAP7_75t_SL g557 ( .A1(n_437), .A2(n_295), .B1(n_275), .B2(n_290), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_442), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_467), .A2(n_323), .B1(n_314), .B2(n_315), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_467), .A2(n_323), .B1(n_314), .B2(n_315), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_481), .B(n_24), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_450), .B(n_142), .Y(n_562) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_437), .A2(n_261), .B1(n_259), .B2(n_295), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_442), .B(n_24), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_473), .A2(n_314), .B1(n_242), .B2(n_296), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_473), .A2(n_314), .B1(n_242), .B2(n_296), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_464), .A2(n_261), .B1(n_259), .B2(n_306), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_441), .B(n_25), .Y(n_568) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_437), .B(n_142), .C(n_146), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_457), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_496), .A2(n_449), .B1(n_444), .B2(n_426), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_502), .B(n_444), .C(n_469), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_558), .B(n_469), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_558), .B(n_444), .Y(n_574) );
NAND4xp25_ASAP7_75t_L g575 ( .A(n_543), .B(n_475), .C(n_472), .D(n_469), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_562), .B(n_471), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_502), .B(n_471), .C(n_475), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_493), .B(n_475), .C(n_472), .D(n_471), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_562), .B(n_450), .Y(n_579) );
OAI221xp5_ASAP7_75t_SL g580 ( .A1(n_497), .A2(n_472), .B1(n_474), .B2(n_457), .C(n_453), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_487), .B(n_142), .C(n_143), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_546), .B(n_453), .Y(n_582) );
OAI21xp33_ASAP7_75t_L g583 ( .A1(n_529), .A2(n_143), .B(n_142), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_491), .B(n_474), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_532), .A2(n_474), .B1(n_428), .B2(n_283), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_570), .B(n_25), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_532), .B(n_142), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_570), .B(n_26), .Y(n_588) );
OAI21xp5_ASAP7_75t_SL g589 ( .A1(n_522), .A2(n_143), .B(n_261), .Y(n_589) );
OA21x2_ASAP7_75t_L g590 ( .A1(n_510), .A2(n_318), .B(n_243), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_487), .A2(n_142), .B1(n_216), .B2(n_259), .C(n_223), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_513), .B(n_26), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_491), .B(n_27), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_532), .B(n_142), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_515), .B(n_27), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_533), .B(n_136), .C(n_282), .Y(n_596) );
OAI221xp5_ASAP7_75t_L g597 ( .A1(n_488), .A2(n_223), .B1(n_276), .B2(n_207), .C(n_268), .Y(n_597) );
OAI21xp5_ASAP7_75t_SL g598 ( .A1(n_518), .A2(n_305), .B(n_295), .Y(n_598) );
NOR3xp33_ASAP7_75t_L g599 ( .A(n_568), .B(n_561), .C(n_555), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_515), .B(n_28), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_508), .B(n_29), .Y(n_601) );
AOI22xp33_ASAP7_75t_SL g602 ( .A1(n_494), .A2(n_305), .B1(n_275), .B2(n_290), .Y(n_602) );
OAI211xp5_ASAP7_75t_SL g603 ( .A1(n_530), .A2(n_227), .B(n_224), .C(n_282), .Y(n_603) );
NOR2xp33_ASAP7_75t_SL g604 ( .A(n_511), .B(n_275), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_495), .B(n_136), .C(n_293), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_567), .A2(n_305), .B1(n_295), .B2(n_290), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_508), .B(n_30), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_519), .B(n_31), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_552), .B(n_136), .C(n_282), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_564), .B(n_32), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_503), .B(n_32), .Y(n_611) );
NOR2xp33_ASAP7_75t_R g612 ( .A(n_501), .B(n_33), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_485), .A2(n_286), .B1(n_296), .B2(n_265), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_549), .B(n_34), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g615 ( .A(n_557), .B(n_305), .C(n_290), .Y(n_615) );
INVxp67_ASAP7_75t_SL g616 ( .A(n_521), .Y(n_616) );
NAND4xp25_ASAP7_75t_L g617 ( .A(n_489), .B(n_265), .C(n_268), .D(n_205), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_567), .A2(n_305), .B1(n_295), .B2(n_290), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_482), .B(n_34), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_500), .A2(n_305), .B(n_295), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_549), .B(n_35), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_514), .B(n_35), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_486), .A2(n_268), .B1(n_265), .B2(n_295), .C(n_290), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_504), .B(n_37), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_485), .A2(n_305), .B1(n_290), .B2(n_301), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_514), .B(n_37), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_494), .B(n_38), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_490), .B(n_39), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_505), .B(n_40), .Y(n_629) );
OA21x2_ASAP7_75t_L g630 ( .A1(n_537), .A2(n_301), .B(n_214), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_520), .B(n_41), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_516), .B(n_42), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_509), .B(n_531), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_556), .B(n_42), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_517), .B(n_43), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_563), .A2(n_136), .B1(n_224), .B2(n_289), .C(n_292), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_556), .B(n_43), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_537), .A2(n_44), .B(n_286), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_525), .B(n_44), .Y(n_639) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_551), .A2(n_547), .B(n_507), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_526), .B(n_263), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_556), .B(n_48), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_498), .A2(n_136), .B1(n_218), .B2(n_226), .C(n_292), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g644 ( .A1(n_557), .A2(n_136), .B(n_218), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g645 ( .A(n_512), .B(n_238), .C(n_289), .D(n_292), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_534), .B(n_286), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_483), .B(n_484), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_527), .A2(n_292), .B1(n_289), .B2(n_195), .C(n_286), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_545), .B(n_263), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_556), .B(n_50), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_528), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_499), .A2(n_292), .B1(n_289), .B2(n_286), .C(n_263), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_538), .A2(n_286), .B1(n_292), .B2(n_289), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_506), .B(n_289), .C(n_241), .D(n_53), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_536), .B(n_286), .C(n_52), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_535), .A2(n_524), .B1(n_523), .B2(n_547), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_544), .B(n_286), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_542), .B(n_286), .Y(n_658) );
OAI21xp5_ASAP7_75t_SL g659 ( .A1(n_550), .A2(n_54), .B(n_55), .Y(n_659) );
OAI21xp33_ASAP7_75t_SL g660 ( .A1(n_633), .A2(n_539), .B(n_553), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g661 ( .A(n_610), .B(n_536), .C(n_569), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_616), .B(n_582), .Y(n_662) );
AO21x2_ASAP7_75t_L g663 ( .A1(n_592), .A2(n_569), .B(n_548), .Y(n_663) );
NOR2xp33_ASAP7_75t_R g664 ( .A(n_604), .B(n_541), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_574), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_633), .B(n_548), .C(n_540), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_573), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_610), .B(n_589), .C(n_619), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_599), .B(n_560), .C(n_559), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_593), .B(n_492), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_601), .B(n_492), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_584), .B(n_492), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_577), .B(n_566), .C(n_565), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_640), .B(n_554), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_608), .B(n_66), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_617), .A2(n_241), .B1(n_69), .B2(n_70), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_579), .Y(n_677) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_572), .B(n_71), .C(n_72), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_607), .B(n_75), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_576), .B(n_77), .Y(n_680) );
NOR2xp33_ASAP7_75t_SL g681 ( .A(n_580), .B(n_78), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_651), .B(n_79), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_647), .B(n_624), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_586), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_587), .B(n_81), .C(n_82), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_588), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_575), .B(n_595), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_600), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_594), .B(n_629), .C(n_620), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_659), .B(n_611), .C(n_628), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_590), .A2(n_83), .B1(n_84), .B2(n_232), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_634), .B(n_590), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_603), .A2(n_656), .B1(n_612), .B2(n_645), .Y(n_693) );
NAND4xp75_ASAP7_75t_L g694 ( .A(n_627), .B(n_626), .C(n_622), .D(n_634), .Y(n_694) );
NAND4xp75_ASAP7_75t_L g695 ( .A(n_590), .B(n_637), .C(n_614), .D(n_650), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_602), .B(n_585), .C(n_578), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_642), .B(n_621), .Y(n_697) );
OA21x2_ASAP7_75t_L g698 ( .A1(n_646), .A2(n_655), .B(n_598), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_646), .Y(n_699) );
NAND3xp33_ASAP7_75t_SL g700 ( .A(n_615), .B(n_612), .C(n_638), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_597), .B(n_583), .C(n_631), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_632), .B(n_635), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_656), .B(n_641), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_654), .A2(n_649), .B1(n_636), .B2(n_630), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_630), .A2(n_625), .B1(n_644), .B2(n_639), .Y(n_705) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_630), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_581), .B(n_653), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_658), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_609), .B(n_657), .Y(n_709) );
NAND4xp75_ASAP7_75t_L g710 ( .A(n_652), .B(n_591), .C(n_643), .D(n_618), .Y(n_710) );
BUFx3_ASAP7_75t_L g711 ( .A(n_648), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_605), .A2(n_623), .B1(n_606), .B2(n_596), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_613), .B(n_616), .Y(n_713) );
NAND3xp33_ASAP7_75t_SL g714 ( .A(n_659), .B(n_620), .C(n_354), .Y(n_714) );
OAI211xp5_ASAP7_75t_SL g715 ( .A1(n_640), .A2(n_533), .B(n_633), .C(n_599), .Y(n_715) );
NAND3xp33_ASAP7_75t_L g716 ( .A(n_633), .B(n_599), .C(n_571), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_616), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_616), .B(n_573), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_610), .B(n_529), .Y(n_719) );
INVx3_ASAP7_75t_L g720 ( .A(n_590), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_633), .B(n_599), .C(n_571), .Y(n_721) );
NAND2xp33_ASAP7_75t_R g722 ( .A(n_590), .B(n_468), .Y(n_722) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_604), .A2(n_354), .B1(n_369), .B2(n_448), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_677), .B(n_662), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_695), .A2(n_723), .B1(n_721), .B2(n_716), .Y(n_725) );
XNOR2x2_ASAP7_75t_L g726 ( .A(n_714), .B(n_674), .Y(n_726) );
NOR4xp75_ASAP7_75t_L g727 ( .A(n_714), .B(n_700), .C(n_694), .D(n_710), .Y(n_727) );
OA22x2_ASAP7_75t_L g728 ( .A1(n_703), .A2(n_692), .B1(n_683), .B2(n_684), .Y(n_728) );
NAND4xp25_ASAP7_75t_L g729 ( .A(n_715), .B(n_693), .C(n_668), .D(n_696), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_667), .B(n_718), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_715), .B(n_719), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_672), .B(n_671), .Y(n_732) );
INVx2_ASAP7_75t_SL g733 ( .A(n_720), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_670), .B(n_720), .Y(n_734) );
XOR2x2_ASAP7_75t_L g735 ( .A(n_668), .B(n_700), .Y(n_735) );
NOR4xp25_ASAP7_75t_L g736 ( .A(n_660), .B(n_686), .C(n_688), .D(n_693), .Y(n_736) );
XNOR2x2_ASAP7_75t_L g737 ( .A(n_689), .B(n_666), .Y(n_737) );
XNOR2x2_ASAP7_75t_L g738 ( .A(n_687), .B(n_669), .Y(n_738) );
NOR2x1_ASAP7_75t_L g739 ( .A(n_698), .B(n_678), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_713), .Y(n_740) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_722), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_699), .B(n_697), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_708), .B(n_663), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_706), .B(n_663), .Y(n_744) );
INVxp67_ASAP7_75t_L g745 ( .A(n_702), .Y(n_745) );
AOI211xp5_ASAP7_75t_SL g746 ( .A1(n_681), .A2(n_704), .B(n_661), .C(n_690), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_706), .B(n_705), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_705), .B(n_711), .Y(n_748) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_682), .Y(n_749) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_661), .Y(n_750) );
NAND3xp33_ASAP7_75t_SL g751 ( .A(n_723), .B(n_664), .C(n_691), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_709), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_707), .Y(n_753) );
NAND4xp75_ASAP7_75t_SL g754 ( .A(n_679), .B(n_680), .C(n_704), .D(n_691), .Y(n_754) );
INVx1_ASAP7_75t_SL g755 ( .A(n_675), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_701), .B(n_690), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_701), .B(n_673), .Y(n_757) );
AND2x4_ASAP7_75t_SL g758 ( .A(n_676), .B(n_712), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_685), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_717), .Y(n_760) );
AND4x1_ASAP7_75t_L g761 ( .A(n_716), .B(n_721), .C(n_681), .D(n_693), .Y(n_761) );
INVx2_ASAP7_75t_SL g762 ( .A(n_665), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_760), .Y(n_763) );
XNOR2x1_ASAP7_75t_L g764 ( .A(n_735), .B(n_726), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_730), .Y(n_765) );
INVxp67_ASAP7_75t_L g766 ( .A(n_731), .Y(n_766) );
INVx1_ASAP7_75t_SL g767 ( .A(n_755), .Y(n_767) );
OR2x2_ASAP7_75t_L g768 ( .A(n_752), .B(n_753), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_762), .Y(n_769) );
NOR2xp33_ASAP7_75t_SL g770 ( .A(n_751), .B(n_741), .Y(n_770) );
INVx1_ASAP7_75t_SL g771 ( .A(n_752), .Y(n_771) );
INVx2_ASAP7_75t_SL g772 ( .A(n_728), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_734), .B(n_732), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_730), .Y(n_774) );
AO22x1_ASAP7_75t_L g775 ( .A1(n_750), .A2(n_747), .B1(n_748), .B2(n_725), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_728), .B(n_736), .Y(n_776) );
INVxp67_ASAP7_75t_L g777 ( .A(n_753), .Y(n_777) );
XOR2x2_ASAP7_75t_L g778 ( .A(n_735), .B(n_727), .Y(n_778) );
OR2x2_ASAP7_75t_L g779 ( .A(n_732), .B(n_740), .Y(n_779) );
INVx2_ASAP7_75t_SL g780 ( .A(n_728), .Y(n_780) );
INVx1_ASAP7_75t_SL g781 ( .A(n_748), .Y(n_781) );
AO22x2_ASAP7_75t_L g782 ( .A1(n_747), .A2(n_740), .B1(n_754), .B2(n_744), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_733), .Y(n_783) );
BUFx2_ASAP7_75t_L g784 ( .A(n_782), .Y(n_784) );
OAI22x1_ASAP7_75t_L g785 ( .A1(n_776), .A2(n_761), .B1(n_738), .B2(n_739), .Y(n_785) );
CKINVDCx16_ASAP7_75t_R g786 ( .A(n_770), .Y(n_786) );
XNOR2x1_ASAP7_75t_L g787 ( .A(n_764), .B(n_726), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_765), .Y(n_788) );
OA22x2_ASAP7_75t_L g789 ( .A1(n_772), .A2(n_757), .B1(n_756), .B2(n_758), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_781), .B(n_724), .Y(n_790) );
AOI22x1_ASAP7_75t_L g791 ( .A1(n_782), .A2(n_746), .B1(n_738), .B2(n_737), .Y(n_791) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_771), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_772), .A2(n_739), .B1(n_745), .B2(n_758), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_763), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_780), .A2(n_733), .B1(n_742), .B2(n_743), .Y(n_795) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_766), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_774), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_768), .Y(n_798) );
INVx1_ASAP7_75t_SL g799 ( .A(n_792), .Y(n_799) );
AOI322xp5_ASAP7_75t_L g800 ( .A1(n_784), .A2(n_786), .A3(n_796), .B1(n_780), .B2(n_787), .C1(n_764), .C2(n_790), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_798), .Y(n_801) );
BUFx2_ASAP7_75t_L g802 ( .A(n_784), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_794), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_788), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_794), .Y(n_805) );
OAI322xp33_ASAP7_75t_L g806 ( .A1(n_787), .A2(n_737), .A3(n_777), .B1(n_768), .B2(n_778), .C1(n_775), .C2(n_767), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_799), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_802), .A2(n_789), .B1(n_778), .B2(n_729), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_806), .A2(n_785), .B1(n_775), .B2(n_793), .C(n_782), .Y(n_809) );
BUFx2_ASAP7_75t_L g810 ( .A(n_801), .Y(n_810) );
AND4x1_ASAP7_75t_L g811 ( .A(n_800), .B(n_789), .C(n_785), .D(n_791), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_807), .Y(n_812) );
O2A1O1Ixp33_ASAP7_75t_L g813 ( .A1(n_809), .A2(n_802), .B(n_801), .C(n_795), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_810), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_812), .A2(n_808), .B1(n_789), .B2(n_782), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_814), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_816), .Y(n_817) );
NOR2xp67_ASAP7_75t_L g818 ( .A(n_815), .B(n_804), .Y(n_818) );
NOR2x1_ASAP7_75t_L g819 ( .A(n_817), .B(n_813), .Y(n_819) );
AO22x2_ASAP7_75t_L g820 ( .A1(n_818), .A2(n_811), .B1(n_805), .B2(n_803), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_820), .Y(n_821) );
INVx1_ASAP7_75t_SL g822 ( .A(n_819), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_821), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_823), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_824), .A2(n_822), .B1(n_797), .B2(n_805), .Y(n_825) );
OR2x2_ASAP7_75t_L g826 ( .A(n_825), .B(n_803), .Y(n_826) );
AOI22xp5_ASAP7_75t_SL g827 ( .A1(n_826), .A2(n_773), .B1(n_759), .B2(n_749), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_827), .Y(n_828) );
AOI221xp5_ASAP7_75t_L g829 ( .A1(n_828), .A2(n_791), .B1(n_773), .B2(n_783), .C(n_744), .Y(n_829) );
AOI211xp5_ASAP7_75t_L g830 ( .A1(n_829), .A2(n_779), .B(n_783), .C(n_769), .Y(n_830) );
endmodule