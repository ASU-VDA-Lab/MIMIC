module real_jpeg_22094_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_276, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_276;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_253;
wire n_96;
wire n_269;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_0),
.A2(n_3),
.B1(n_18),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_54),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_0),
.A2(n_5),
.B1(n_54),
.B2(n_65),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_3),
.B1(n_18),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_1),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_1),
.A2(n_5),
.B1(n_30),
.B2(n_65),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_2),
.A2(n_3),
.B1(n_18),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_5),
.B1(n_50),
.B2(n_65),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_50),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_2),
.A2(n_23),
.B(n_27),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_2),
.B(n_28),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_2),
.A2(n_5),
.B(n_10),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_2),
.B(n_37),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_SL g165 ( 
.A1(n_2),
.A2(n_40),
.B(n_41),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_3),
.A2(n_7),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_3),
.A2(n_24),
.B(n_50),
.C(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_4),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_10),
.B1(n_63),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_7),
.B1(n_19),
.B2(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_5),
.B(n_94),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_7),
.A2(n_19),
.B1(n_39),
.B2(n_40),
.Y(n_220)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_9),
.A2(n_18),
.B(n_22),
.C(n_25),
.Y(n_21)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_9),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_69),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_67),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_31),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_31),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_17),
.A2(n_25),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_20),
.A2(n_28),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_21),
.B(n_25),
.Y(n_239)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_38),
.B(n_41),
.C(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_41),
.Y(n_45)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_27),
.A2(n_42),
.B(n_50),
.C(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_28),
.A2(n_48),
.B(n_53),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_32),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_32),
.B(n_273),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_46),
.CI(n_51),
.CON(n_32),
.SN(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_37),
.B1(n_43),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_36),
.B(n_99),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_37),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_38),
.A2(n_44),
.B1(n_99),
.B2(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_38),
.A2(n_252),
.B(n_253),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_40),
.A2(n_50),
.B(n_63),
.C(n_141),
.Y(n_140)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_44),
.B(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_50),
.B(n_87),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_50),
.B(n_64),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.C(n_58),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_52),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_52),
.B(n_108),
.C(n_109),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_52),
.A2(n_96),
.B1(n_107),
.B2(n_120),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_52),
.B(n_96),
.C(n_215),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_52),
.A2(n_107),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_55),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_56),
.A2(n_58),
.B1(n_250),
.B2(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_56),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_57),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_58),
.A2(n_250),
.B1(n_251),
.B2(n_254),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_58),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_66),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_61),
.A2(n_64),
.B1(n_81),
.B2(n_84),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_61),
.A2(n_64),
.B1(n_66),
.B2(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_64),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_65),
.B(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_272),
.B(n_274),
.Y(n_69)
);

OAI321xp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_245),
.A3(n_265),
.B1(n_270),
.B2(n_271),
.C(n_276),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_228),
.B(n_244),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_209),
.B(n_227),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_130),
.B(n_190),
.C(n_208),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_115),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_75),
.B(n_115),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_103),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_95),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_77),
.B(n_95),
.C(n_103),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_85),
.B2(n_86),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_79),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_78),
.A2(n_79),
.B1(n_96),
.B2(n_120),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_78),
.B(n_86),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_79),
.B(n_140),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_79),
.B(n_96),
.C(n_163),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_83),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_83),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_89),
.Y(n_86)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_87),
.B(n_93),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_87),
.A2(n_88),
.B1(n_93),
.B2(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_114),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_90),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_93),
.B1(n_94),
.B2(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_102),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_100),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_98),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_117),
.B1(n_118),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_102),
.A2(n_117),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_102),
.B(n_202),
.C(n_204),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_102),
.A2(n_117),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_102),
.A2(n_117),
.B1(n_259),
.B2(n_263),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_105),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_125),
.C(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_105),
.A2(n_108),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_105),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_105),
.B(n_234),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_147),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_123),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_155),
.C(n_158),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.C(n_124),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_116),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_117),
.B(n_250),
.C(n_254),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_117),
.B(n_263),
.C(n_264),
.Y(n_273)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_124),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_137),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_189),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_184),
.B(n_188),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_172),
.B(n_183),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_160),
.B(n_171),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_150),
.B(n_159),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_142),
.B(n_149),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_138),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B(n_148),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_152),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_158),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_158),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_175),
.C(n_182),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_162),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_170),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_166),
.B1(n_167),
.B2(n_169),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_164),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_169),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_173),
.B(n_174),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_181),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_186),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_191),
.B(n_192),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_206),
.B2(n_207),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_200),
.B2(n_201),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_201),
.C(n_207),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_206),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_211),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_226),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_217),
.B2(n_218),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_218),
.C(n_226),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_223),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_223),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_238),
.B(n_241),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_230),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_242),
.B2(n_243),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_236),
.C(n_243),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_247),
.C(n_255),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_247),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_238),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_257),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_251),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_255),
.A2(n_256),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_264),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_259),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_268),
.Y(n_269)
);


endmodule