module fake_jpeg_21457_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_68),
.Y(n_76)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_41),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_56),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_41),
.B1(n_42),
.B2(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_77),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

AO22x1_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_63),
.B1(n_2),
.B2(n_1),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_1),
.Y(n_94)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_82),
.A2(n_42),
.B1(n_58),
.B2(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_4),
.B1(n_5),
.B2(n_11),
.Y(n_106)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_91),
.Y(n_99)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_92),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_55),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_3),
.Y(n_100)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_57),
.B1(n_50),
.B2(n_61),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_19),
.B(n_22),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_101),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_53),
.B1(n_45),
.B2(n_6),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_106),
.B(n_17),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_107),
.B(n_38),
.Y(n_110)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_112),
.C(n_114),
.Y(n_117)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_26),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_97),
.B(n_115),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_118),
.B(n_111),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_107),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_110),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_120),
.Y(n_124)
);

OAI21x1_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_117),
.B(n_30),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_102),
.B1(n_105),
.B2(n_108),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_33),
.Y(n_129)
);


endmodule