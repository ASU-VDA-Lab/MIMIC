module fake_jpeg_2802_n_91 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_25),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_43),
.Y(n_47)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_26),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_43),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_41),
.B(n_1),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_36),
.B1(n_35),
.B2(n_24),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_30),
.Y(n_59)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_14),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_54),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_28),
.B1(n_38),
.B2(n_29),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_28),
.B1(n_30),
.B2(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_0),
.C(n_1),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_55),
.B1(n_57),
.B2(n_56),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_74),
.B1(n_7),
.B2(n_10),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_8),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_15),
.C(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_5),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_6),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_3),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_79),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_5),
.Y(n_76)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_83),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_69),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_68),
.C(n_71),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_89),
.A2(n_84),
.B(n_76),
.C(n_80),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_81),
.Y(n_91)
);


endmodule