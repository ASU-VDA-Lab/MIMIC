module fake_netlist_1_1948_n_19 (n_1, n_2, n_0, n_19);
input n_1;
input n_2;
input n_0;
output n_19;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_3;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_6;
wire n_4;
wire n_7;
INVx1_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
INVx3_ASAP7_75t_SL g6 ( .A(n_5), .Y(n_6) );
OAI21x1_ASAP7_75t_L g7 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_7) );
OAI21x1_ASAP7_75t_SL g8 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_8) );
BUFx6f_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
AND2x4_ASAP7_75t_L g11 ( .A(n_10), .B(n_7), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_9), .B(n_8), .Y(n_13) );
NAND3x1_ASAP7_75t_L g14 ( .A(n_11), .B(n_3), .C(n_2), .Y(n_14) );
OAI211xp5_ASAP7_75t_L g15 ( .A1(n_13), .A2(n_12), .B(n_6), .C(n_2), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
AOI22xp33_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_0), .B1(n_11), .B2(n_15), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
AO21x2_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_11), .B(n_17), .Y(n_19) );
endmodule