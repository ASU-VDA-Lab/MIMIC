module fake_netlist_1_5408_n_511 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_511);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_511;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g74 ( .A(n_61), .Y(n_74) );
HB1xp67_ASAP7_75t_L g75 ( .A(n_49), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_51), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_2), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_20), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_59), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_52), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_6), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_0), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_23), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_64), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_7), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_11), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_45), .Y(n_87) );
BUFx6f_ASAP7_75t_SL g88 ( .A(n_46), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_29), .Y(n_89) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_58), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_36), .Y(n_91) );
BUFx3_ASAP7_75t_L g92 ( .A(n_18), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_15), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_72), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_42), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_5), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_63), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_50), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_1), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_22), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_11), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_28), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_31), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_15), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_17), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_26), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_16), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_5), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_71), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_30), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_24), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_101), .B(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_78), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_78), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_95), .Y(n_116) );
BUFx8_ASAP7_75t_L g117 ( .A(n_88), .Y(n_117) );
AND2x4_ASAP7_75t_L g118 ( .A(n_81), .B(n_1), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_86), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_86), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_120) );
CKINVDCx8_ASAP7_75t_R g121 ( .A(n_98), .Y(n_121) );
AND2x2_ASAP7_75t_SL g122 ( .A(n_75), .B(n_73), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_97), .Y(n_124) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_83), .A2(n_39), .B(n_69), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_95), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_81), .B(n_3), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_82), .B(n_4), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_90), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_118), .Y(n_134) );
INVx1_ASAP7_75t_SL g135 ( .A(n_119), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_118), .Y(n_136) );
INVx4_ASAP7_75t_L g137 ( .A(n_118), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_118), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_114), .B(n_82), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_129), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_125), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_114), .B(n_85), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_129), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_115), .B(n_76), .Y(n_145) );
OR2x2_ASAP7_75t_L g146 ( .A(n_113), .B(n_104), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_115), .B(n_79), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_123), .B(n_85), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g150 ( .A(n_113), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_123), .B(n_91), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_126), .B(n_131), .Y(n_152) );
INVx2_ASAP7_75t_SL g153 ( .A(n_117), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_124), .B(n_74), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_125), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_126), .B(n_97), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_137), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_153), .B(n_117), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_134), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_141), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_156), .A2(n_122), .B1(n_130), .B2(n_128), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_153), .B(n_117), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_156), .B(n_131), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_156), .B(n_117), .Y(n_164) );
INVx1_ASAP7_75t_SL g165 ( .A(n_135), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_154), .B(n_121), .Y(n_166) );
AO22x1_ASAP7_75t_L g167 ( .A1(n_134), .A2(n_74), .B1(n_122), .B2(n_87), .Y(n_167) );
AND2x6_ASAP7_75t_SL g168 ( .A(n_139), .B(n_128), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_136), .A2(n_122), .B1(n_130), .B2(n_99), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_136), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_153), .B(n_121), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_135), .B(n_107), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_137), .B(n_100), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g179 ( .A1(n_146), .A2(n_120), .B1(n_104), .B2(n_96), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_152), .B(n_116), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_152), .B(n_127), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_137), .A2(n_77), .B1(n_110), .B2(n_108), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_149), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_139), .B(n_127), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_139), .B(n_112), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_165), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_159), .A2(n_142), .B(n_155), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_165), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_163), .A2(n_146), .B(n_151), .C(n_145), .Y(n_190) );
OR2x6_ASAP7_75t_L g191 ( .A(n_174), .B(n_146), .Y(n_191) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_157), .B(n_143), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_164), .B(n_143), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
OAI21xp33_ASAP7_75t_L g195 ( .A1(n_161), .A2(n_147), .B(n_151), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_172), .B(n_143), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_157), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_159), .A2(n_147), .B(n_145), .C(n_148), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_170), .A2(n_142), .B(n_155), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_163), .B(n_148), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_166), .B(n_148), .Y(n_201) );
CKINVDCx11_ASAP7_75t_R g202 ( .A(n_168), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_SL g203 ( .A1(n_183), .A2(n_149), .B(n_132), .C(n_129), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_186), .A2(n_149), .B(n_112), .C(n_80), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_170), .A2(n_142), .B(n_155), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_181), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_177), .A2(n_142), .B(n_155), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_169), .A2(n_120), .B1(n_149), .B2(n_142), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_185), .B(n_142), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g212 ( .A1(n_185), .A2(n_93), .B1(n_142), .B2(n_89), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_175), .B(n_177), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_175), .B(n_109), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_168), .B(n_111), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_207), .B(n_167), .Y(n_216) );
AO31x2_ASAP7_75t_L g217 ( .A1(n_198), .A2(n_180), .A3(n_186), .B(n_133), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_201), .A2(n_182), .B1(n_181), .B2(n_180), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_211), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_188), .A2(n_208), .B(n_199), .Y(n_220) );
INVx8_ASAP7_75t_L g221 ( .A(n_191), .Y(n_221) );
AO31x2_ASAP7_75t_L g222 ( .A1(n_210), .A2(n_133), .A3(n_182), .B(n_94), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_206), .A2(n_184), .B(n_175), .Y(n_223) );
NOR2xp67_ASAP7_75t_L g224 ( .A(n_189), .B(n_175), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_213), .A2(n_184), .B(n_160), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_187), .B(n_171), .Y(n_226) );
OAI221xp5_ASAP7_75t_L g227 ( .A1(n_215), .A2(n_179), .B1(n_173), .B2(n_162), .C(n_158), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_196), .B(n_190), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_209), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_192), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_192), .Y(n_231) );
INVx6_ASAP7_75t_L g232 ( .A(n_204), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_191), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_197), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_195), .A2(n_179), .B1(n_167), .B2(n_176), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_193), .A2(n_176), .B(n_160), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_197), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_204), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_204), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_205), .A2(n_176), .B(n_160), .C(n_106), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_227), .A2(n_202), .B1(n_191), .B2(n_210), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_221), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_229), .Y(n_243) );
OAI221xp5_ASAP7_75t_L g244 ( .A1(n_228), .A2(n_194), .B1(n_200), .B2(n_203), .C(n_214), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_218), .A2(n_212), .B(n_125), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_229), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_219), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_231), .B(n_93), .Y(n_248) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_220), .A2(n_133), .B(n_103), .Y(n_249) );
AOI22xp33_ASAP7_75t_SL g250 ( .A1(n_221), .A2(n_88), .B1(n_92), .B2(n_105), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_223), .A2(n_125), .B(n_102), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_231), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_236), .A2(n_144), .B(n_141), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_219), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_234), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_230), .B(n_92), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_222), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_233), .A2(n_235), .B1(n_216), .B2(n_221), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_225), .A2(n_132), .B(n_144), .Y(n_259) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_233), .A2(n_93), .B1(n_105), .B2(n_90), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_234), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_254), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_257), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_254), .B(n_217), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_247), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_247), .Y(n_266) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_257), .A2(n_240), .B(n_224), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_259), .A2(n_239), .B(n_237), .Y(n_268) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_245), .A2(n_224), .B(n_222), .Y(n_269) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_252), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_243), .B(n_217), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_243), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_246), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_241), .A2(n_221), .B1(n_226), .B2(n_230), .Y(n_274) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_251), .A2(n_222), .B(n_237), .Y(n_275) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_259), .A2(n_222), .B(n_217), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_246), .B(n_217), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_258), .A2(n_226), .B1(n_93), .B2(n_232), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_252), .B(n_217), .Y(n_279) );
OR2x6_ASAP7_75t_L g280 ( .A(n_252), .B(n_232), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_244), .B(n_226), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_263), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_273), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_263), .Y(n_284) );
AO21x2_ASAP7_75t_L g285 ( .A1(n_269), .A2(n_248), .B(n_260), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_279), .B(n_222), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_281), .A2(n_226), .B1(n_250), .B2(n_256), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_263), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_280), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_279), .B(n_261), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_265), .B(n_261), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_271), .B(n_249), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_264), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_270), .Y(n_294) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_269), .A2(n_256), .B(n_255), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_265), .B(n_255), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_273), .B(n_256), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_264), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_270), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_271), .B(n_249), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_264), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_266), .B(n_256), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_271), .B(n_249), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_277), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_277), .B(n_249), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_277), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_279), .B(n_273), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_262), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_307), .B(n_276), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_282), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_304), .B(n_262), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_304), .B(n_276), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_308), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_306), .B(n_266), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_284), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_307), .B(n_276), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_294), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_307), .B(n_276), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_304), .B(n_276), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_308), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_294), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_282), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_284), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_293), .B(n_269), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_293), .B(n_269), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_291), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_291), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_306), .B(n_272), .Y(n_328) );
INVx2_ASAP7_75t_SL g329 ( .A(n_299), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_293), .B(n_272), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_298), .B(n_269), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_298), .B(n_275), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_298), .B(n_281), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_301), .B(n_275), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_282), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_296), .Y(n_337) );
NAND4xp25_ASAP7_75t_L g338 ( .A(n_287), .B(n_278), .C(n_274), .D(n_286), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_299), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_297), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_301), .B(n_275), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_301), .B(n_275), .Y(n_342) );
NOR2xp67_ASAP7_75t_L g343 ( .A(n_286), .B(n_274), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_297), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_290), .B(n_278), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_288), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_290), .B(n_280), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_286), .B(n_275), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_317), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_320), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_326), .B(n_286), .Y(n_352) );
INVx3_ASAP7_75t_L g353 ( .A(n_348), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_335), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_344), .B(n_290), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_313), .B(n_290), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_311), .B(n_283), .Y(n_357) );
AOI211xp5_ASAP7_75t_L g358 ( .A1(n_338), .A2(n_289), .B(n_303), .C(n_300), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_326), .B(n_303), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_328), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_327), .B(n_303), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_309), .B(n_292), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_328), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_327), .B(n_302), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_330), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_334), .B(n_302), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_334), .B(n_300), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_340), .B(n_300), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_340), .B(n_292), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_330), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_314), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_335), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_337), .B(n_292), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_337), .Y(n_374) );
AND3x2_ASAP7_75t_L g375 ( .A(n_317), .B(n_305), .C(n_288), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_348), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_329), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_315), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_309), .B(n_305), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_315), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_329), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_316), .B(n_295), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_323), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_316), .B(n_283), .Y(n_384) );
INVx2_ASAP7_75t_SL g385 ( .A(n_339), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_323), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_311), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_318), .B(n_295), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_333), .Y(n_389) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_339), .B(n_289), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_318), .B(n_349), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_349), .B(n_295), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_321), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_324), .B(n_295), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_345), .B(n_289), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_347), .B(n_267), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_312), .B(n_319), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_332), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_381), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_382), .B(n_324), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_377), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_358), .A2(n_343), .B1(n_325), .B2(n_342), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_391), .B(n_343), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_375), .B(n_332), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_391), .B(n_325), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_350), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_389), .B(n_342), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_379), .B(n_341), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_382), .B(n_341), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_388), .B(n_312), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_351), .Y(n_412) );
NAND4xp25_ASAP7_75t_SL g413 ( .A(n_392), .B(n_331), .C(n_319), .D(n_310), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_379), .B(n_331), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_362), .B(n_336), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_355), .A2(n_336), .B1(n_322), .B2(n_310), .Y(n_416) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_377), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_378), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_380), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_383), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_374), .Y(n_422) );
OA211x2_ASAP7_75t_L g423 ( .A1(n_375), .A2(n_6), .B(n_7), .C(n_8), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_360), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_363), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_388), .B(n_346), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_385), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_365), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_385), .B(n_322), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_371), .B(n_9), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_362), .B(n_348), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_356), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_370), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_368), .B(n_346), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_394), .B(n_285), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_352), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_397), .B(n_267), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_398), .B(n_267), .Y(n_440) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_353), .B(n_242), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_422), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_411), .B(n_394), .Y(n_443) );
OAI21xp33_ASAP7_75t_L g444 ( .A1(n_413), .A2(n_392), .B(n_367), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_402), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_431), .A2(n_364), .B1(n_366), .B2(n_395), .C(n_361), .Y(n_446) );
INVxp33_ASAP7_75t_L g447 ( .A(n_405), .Y(n_447) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_399), .B(n_395), .C(n_364), .Y(n_448) );
OAI211xp5_ASAP7_75t_L g449 ( .A1(n_403), .A2(n_366), .B(n_359), .C(n_373), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_418), .Y(n_450) );
OAI22xp33_ASAP7_75t_L g451 ( .A1(n_405), .A2(n_390), .B1(n_384), .B2(n_353), .Y(n_451) );
OAI322xp33_ASAP7_75t_L g452 ( .A1(n_433), .A2(n_396), .A3(n_354), .B1(n_372), .B2(n_357), .C1(n_369), .C2(n_390), .Y(n_452) );
AOI21xp33_ASAP7_75t_L g453 ( .A1(n_430), .A2(n_90), .B(n_10), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_412), .B(n_372), .C(n_354), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_427), .B(n_353), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_438), .B(n_376), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_417), .A2(n_242), .B(n_376), .C(n_90), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_411), .B(n_285), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_402), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_436), .B(n_285), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_423), .A2(n_280), .B1(n_285), .B2(n_267), .Y(n_461) );
OAI21xp33_ASAP7_75t_L g462 ( .A1(n_437), .A2(n_132), .B(n_280), .Y(n_462) );
OAI222xp33_ASAP7_75t_L g463 ( .A1(n_404), .A2(n_280), .B1(n_238), .B2(n_239), .C1(n_267), .C2(n_14), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_432), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_428), .B(n_268), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_435), .Y(n_466) );
AOI21xp33_ASAP7_75t_SL g467 ( .A1(n_441), .A2(n_9), .B(n_10), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_419), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_441), .A2(n_280), .B(n_268), .Y(n_469) );
NAND2x1_ASAP7_75t_SL g470 ( .A(n_447), .B(n_407), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_442), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_450), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_444), .A2(n_424), .B1(n_425), .B2(n_434), .C(n_416), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_452), .A2(n_416), .B1(n_437), .B2(n_408), .C(n_400), .Y(n_474) );
NOR3xp33_ASAP7_75t_L g475 ( .A(n_453), .B(n_429), .C(n_401), .Y(n_475) );
XNOR2xp5_ASAP7_75t_L g476 ( .A(n_448), .B(n_415), .Y(n_476) );
AOI211xp5_ASAP7_75t_L g477 ( .A1(n_451), .A2(n_439), .B(n_440), .C(n_426), .Y(n_477) );
AOI322xp5_ASAP7_75t_L g478 ( .A1(n_446), .A2(n_410), .A3(n_400), .B1(n_409), .B2(n_406), .C1(n_426), .C2(n_420), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_468), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_449), .B(n_410), .Y(n_480) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_445), .A2(n_414), .B1(n_421), .B2(n_239), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_453), .A2(n_88), .B1(n_253), .B2(n_238), .C(n_13), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_467), .A2(n_12), .B(n_13), .C(n_14), .Y(n_483) );
OAI21xp33_ASAP7_75t_L g484 ( .A1(n_458), .A2(n_268), .B(n_144), .Y(n_484) );
AOI322xp5_ASAP7_75t_L g485 ( .A1(n_443), .A2(n_12), .A3(n_140), .B1(n_21), .B2(n_25), .C1(n_27), .C2(n_32), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_443), .B(n_19), .Y(n_486) );
AOI322xp5_ASAP7_75t_L g487 ( .A1(n_480), .A2(n_466), .A3(n_464), .B1(n_459), .B2(n_455), .C1(n_460), .C2(n_462), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_SL g488 ( .A1(n_486), .A2(n_469), .B(n_461), .C(n_465), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_483), .A2(n_457), .B(n_463), .C(n_456), .Y(n_489) );
AOI211xp5_ASAP7_75t_SL g490 ( .A1(n_482), .A2(n_454), .B(n_34), .C(n_35), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_478), .B(n_33), .Y(n_491) );
NAND4xp75_ASAP7_75t_L g492 ( .A(n_474), .B(n_232), .C(n_38), .D(n_40), .Y(n_492) );
NAND4xp25_ASAP7_75t_L g493 ( .A(n_473), .B(n_140), .C(n_41), .D(n_43), .Y(n_493) );
OAI211xp5_ASAP7_75t_SL g494 ( .A1(n_477), .A2(n_37), .B(n_44), .C(n_47), .Y(n_494) );
AOI211xp5_ASAP7_75t_SL g495 ( .A1(n_481), .A2(n_48), .B(n_53), .C(n_54), .Y(n_495) );
NOR3xp33_ASAP7_75t_L g496 ( .A(n_491), .B(n_486), .C(n_475), .Y(n_496) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_488), .A2(n_484), .B(n_476), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_487), .B(n_479), .Y(n_498) );
OAI211xp5_ASAP7_75t_L g499 ( .A1(n_489), .A2(n_470), .B(n_485), .C(n_471), .Y(n_499) );
OAI211xp5_ASAP7_75t_SL g500 ( .A1(n_490), .A2(n_472), .B(n_56), .C(n_57), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_496), .B(n_492), .Y(n_501) );
AOI211xp5_ASAP7_75t_SL g502 ( .A1(n_499), .A2(n_494), .B(n_493), .C(n_495), .Y(n_502) );
NAND4xp75_ASAP7_75t_L g503 ( .A(n_498), .B(n_55), .C(n_60), .D(n_62), .Y(n_503) );
XNOR2x1_ASAP7_75t_L g504 ( .A(n_501), .B(n_497), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_503), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_504), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_506), .A2(n_505), .B1(n_500), .B2(n_502), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_507), .B(n_65), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_508), .B(n_66), .Y(n_509) );
NAND2x1_ASAP7_75t_L g510 ( .A(n_509), .B(n_232), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_510), .A2(n_67), .B1(n_68), .B2(n_70), .Y(n_511) );
endmodule