module real_aes_8016_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_316;
wire n_532;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_404;
wire n_147;
wire n_288;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g502 ( .A1(n_0), .A2(n_166), .B(n_503), .C(n_506), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_1), .B(n_498), .Y(n_507) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
INVx1_ASAP7_75t_L g164 ( .A(n_3), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_4), .B(n_167), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_5), .A2(n_466), .B(n_542), .Y(n_541) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_6), .A2(n_174), .B(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_7), .A2(n_36), .B1(n_154), .B2(n_202), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_8), .B(n_174), .Y(n_182) );
AND2x6_ASAP7_75t_L g169 ( .A(n_9), .B(n_170), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_10), .A2(n_169), .B(n_471), .C(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_11), .B(n_37), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_11), .B(n_37), .Y(n_122) );
INVx1_ASAP7_75t_L g148 ( .A(n_12), .Y(n_148) );
INVx1_ASAP7_75t_L g145 ( .A(n_13), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_14), .B(n_150), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_15), .B(n_167), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_16), .B(n_141), .Y(n_248) );
AO32x2_ASAP7_75t_L g218 ( .A1(n_17), .A2(n_140), .A3(n_174), .B1(n_193), .B2(n_219), .Y(n_218) );
AOI222xp33_ASAP7_75t_SL g124 ( .A1(n_18), .A2(n_40), .B1(n_125), .B2(n_744), .C1(n_745), .C2(n_747), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_19), .B(n_154), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_20), .B(n_141), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_21), .A2(n_54), .B1(n_154), .B2(n_202), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g204 ( .A1(n_22), .A2(n_80), .B1(n_150), .B2(n_154), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_23), .B(n_154), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_24), .A2(n_193), .B(n_471), .C(n_489), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_25), .A2(n_193), .B(n_471), .C(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_26), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_27), .B(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_28), .A2(n_466), .B(n_500), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_29), .A2(n_101), .B1(n_111), .B2(n_757), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_30), .B(n_195), .Y(n_236) );
INVx2_ASAP7_75t_L g152 ( .A(n_31), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_32), .A2(n_469), .B(n_473), .C(n_479), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_33), .B(n_154), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_34), .B(n_195), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_35), .B(n_213), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_38), .B(n_487), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_39), .Y(n_519) );
INVx1_ASAP7_75t_L g744 ( .A(n_40), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_41), .B(n_167), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_42), .B(n_466), .Y(n_522) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_43), .A2(n_128), .B1(n_129), .B2(n_450), .Y(n_127) );
INVx1_ASAP7_75t_L g450 ( .A(n_43), .Y(n_450) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_43), .A2(n_45), .B1(n_450), .B2(n_756), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_44), .A2(n_469), .B(n_479), .C(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_45), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_46), .B(n_154), .Y(n_177) );
INVx1_ASAP7_75t_L g504 ( .A(n_47), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_48), .A2(n_89), .B1(n_202), .B2(n_203), .Y(n_201) );
INVx1_ASAP7_75t_L g535 ( .A(n_49), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_50), .B(n_154), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_51), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_52), .B(n_466), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_53), .B(n_162), .Y(n_181) );
AOI22xp33_ASAP7_75t_SL g246 ( .A1(n_55), .A2(n_59), .B1(n_150), .B2(n_154), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_56), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_57), .B(n_154), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_58), .B(n_154), .Y(n_210) );
INVx1_ASAP7_75t_L g170 ( .A(n_60), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_61), .B(n_466), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_62), .B(n_498), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_63), .A2(n_156), .B(n_162), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_64), .B(n_154), .Y(n_165) );
INVx1_ASAP7_75t_L g144 ( .A(n_65), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_66), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_67), .B(n_167), .Y(n_477) );
AO32x2_ASAP7_75t_L g199 ( .A1(n_68), .A2(n_174), .A3(n_193), .B1(n_200), .B2(n_205), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_69), .B(n_168), .Y(n_516) );
INVx1_ASAP7_75t_L g189 ( .A(n_70), .Y(n_189) );
INVx1_ASAP7_75t_L g231 ( .A(n_71), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g501 ( .A(n_72), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_73), .B(n_476), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_74), .A2(n_471), .B(n_479), .C(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_75), .B(n_150), .Y(n_232) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_76), .Y(n_543) );
INVx1_ASAP7_75t_L g110 ( .A(n_77), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_78), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_79), .B(n_475), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_81), .B(n_202), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_82), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_83), .B(n_150), .Y(n_235) );
INVx2_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_85), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_86), .B(n_192), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_87), .B(n_150), .Y(n_178) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_88), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g119 ( .A(n_88), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g453 ( .A(n_88), .B(n_121), .Y(n_453) );
INVx2_ASAP7_75t_L g457 ( .A(n_88), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_90), .A2(n_99), .B1(n_150), .B2(n_151), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_91), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g474 ( .A(n_92), .Y(n_474) );
INVxp67_ASAP7_75t_L g546 ( .A(n_93), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_94), .B(n_150), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_95), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g512 ( .A(n_96), .Y(n_512) );
INVx1_ASAP7_75t_L g570 ( .A(n_97), .Y(n_570) );
AND2x2_ASAP7_75t_L g537 ( .A(n_98), .B(n_195), .Y(n_537) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_103), .Y(n_757) );
CKINVDCx12_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g121 ( .A(n_107), .B(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_124), .B1(n_750), .B2(n_752), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g751 ( .A(n_116), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_117), .A2(n_119), .B(n_753), .Y(n_752) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_123), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NOR2x2_ASAP7_75t_L g749 ( .A(n_120), .B(n_457), .Y(n_749) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g456 ( .A(n_121), .B(n_457), .Y(n_456) );
OAI22x1_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_451), .B1(n_454), .B2(n_458), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_127), .A2(n_451), .B1(n_456), .B2(n_746), .Y(n_745) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_128), .A2(n_129), .B1(n_754), .B2(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_130), .B(n_416), .Y(n_129) );
NOR3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_320), .C(n_404), .Y(n_130) );
NAND4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_263), .C(n_285), .D(n_301), .Y(n_131) );
AOI221xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_196), .B1(n_222), .B2(n_241), .C(n_249), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_172), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_135), .B(n_241), .Y(n_275) );
NAND4xp25_ASAP7_75t_L g315 ( .A(n_135), .B(n_303), .C(n_316), .D(n_318), .Y(n_315) );
INVxp67_ASAP7_75t_L g432 ( .A(n_135), .Y(n_432) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g314 ( .A(n_136), .B(n_252), .Y(n_314) );
AND2x2_ASAP7_75t_L g338 ( .A(n_136), .B(n_172), .Y(n_338) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g305 ( .A(n_137), .B(n_240), .Y(n_305) );
AND2x2_ASAP7_75t_L g345 ( .A(n_137), .B(n_326), .Y(n_345) );
AND2x2_ASAP7_75t_L g362 ( .A(n_137), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_137), .B(n_173), .Y(n_386) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g239 ( .A(n_138), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g257 ( .A(n_138), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g269 ( .A(n_138), .B(n_173), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_138), .B(n_183), .Y(n_291) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_146), .B(n_171), .Y(n_138) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_139), .A2(n_184), .B(n_194), .Y(n_183) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_140), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_142), .B(n_143), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_160), .B(n_169), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_153), .C(n_156), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_149), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_149), .A2(n_525), .B(n_526), .Y(n_524) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g155 ( .A(n_152), .Y(n_155) );
INVx1_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
INVx3_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_154), .Y(n_572) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_155), .Y(n_203) );
AND2x6_ASAP7_75t_L g471 ( .A(n_155), .B(n_472), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g569 ( .A1(n_156), .A2(n_570), .B(n_571), .C(n_572), .Y(n_569) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_157), .A2(n_234), .B(n_235), .Y(n_233) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g476 ( .A(n_158), .Y(n_476) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g168 ( .A(n_159), .Y(n_168) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
INVx1_ASAP7_75t_L g213 ( .A(n_159), .Y(n_213) );
AND2x2_ASAP7_75t_L g467 ( .A(n_159), .B(n_163), .Y(n_467) );
INVx1_ASAP7_75t_L g472 ( .A(n_159), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_164), .B(n_165), .C(n_166), .Y(n_160) );
O2A1O1Ixp5_ASAP7_75t_L g188 ( .A1(n_161), .A2(n_189), .B(n_190), .C(n_191), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_161), .A2(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_166), .A2(n_180), .B(n_181), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_166), .A2(n_192), .B1(n_220), .B2(n_221), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_166), .A2(n_192), .B1(n_245), .B2(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_167), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_167), .A2(n_186), .B(n_187), .Y(n_185) );
O2A1O1Ixp5_ASAP7_75t_SL g229 ( .A1(n_167), .A2(n_230), .B(n_231), .C(n_232), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_167), .B(n_546), .Y(n_545) );
INVx5_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_168), .A2(n_192), .B1(n_201), .B2(n_204), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g175 ( .A1(n_169), .A2(n_176), .B(n_179), .Y(n_175) );
BUFx3_ASAP7_75t_L g193 ( .A(n_169), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_169), .A2(n_209), .B(n_214), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_169), .A2(n_229), .B(n_233), .Y(n_228) );
AND2x4_ASAP7_75t_L g466 ( .A(n_169), .B(n_467), .Y(n_466) );
INVx4_ASAP7_75t_SL g480 ( .A(n_169), .Y(n_480) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_169), .B(n_467), .Y(n_513) );
AND2x2_ASAP7_75t_L g272 ( .A(n_172), .B(n_273), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_172), .A2(n_322), .B1(n_325), .B2(n_327), .C(n_331), .Y(n_321) );
AND2x2_ASAP7_75t_L g380 ( .A(n_172), .B(n_345), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_172), .B(n_362), .Y(n_414) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_183), .Y(n_172) );
INVx3_ASAP7_75t_L g240 ( .A(n_173), .Y(n_240) );
AND2x2_ASAP7_75t_L g289 ( .A(n_173), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g343 ( .A(n_173), .B(n_258), .Y(n_343) );
AND2x2_ASAP7_75t_L g401 ( .A(n_173), .B(n_402), .Y(n_401) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_182), .Y(n_173) );
INVx4_ASAP7_75t_L g243 ( .A(n_174), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_174), .A2(n_522), .B(n_523), .Y(n_521) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_174), .Y(n_540) );
AND2x2_ASAP7_75t_L g241 ( .A(n_183), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
INVx1_ASAP7_75t_L g313 ( .A(n_183), .Y(n_313) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_183), .Y(n_319) );
AND2x2_ASAP7_75t_L g364 ( .A(n_183), .B(n_240), .Y(n_364) );
OR2x2_ASAP7_75t_L g403 ( .A(n_183), .B(n_242), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_188), .B(n_193), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_191), .A2(n_215), .B(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx4_ASAP7_75t_L g505 ( .A(n_192), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g262 ( .A(n_193), .B(n_243), .C(n_244), .Y(n_262) );
INVx2_ASAP7_75t_L g205 ( .A(n_195), .Y(n_205) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_195), .A2(n_208), .B(n_217), .Y(n_207) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_195), .A2(n_228), .B(n_236), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_195), .A2(n_465), .B(n_468), .Y(n_464) );
INVx1_ASAP7_75t_L g495 ( .A(n_195), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_195), .A2(n_532), .B(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_196), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_206), .Y(n_196) );
AND2x2_ASAP7_75t_L g399 ( .A(n_197), .B(n_396), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_197), .B(n_381), .Y(n_431) );
BUFx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g330 ( .A(n_198), .B(n_254), .Y(n_330) );
AND2x2_ASAP7_75t_L g379 ( .A(n_198), .B(n_225), .Y(n_379) );
INVx1_ASAP7_75t_L g425 ( .A(n_198), .Y(n_425) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_199), .Y(n_238) );
AND2x2_ASAP7_75t_L g280 ( .A(n_199), .B(n_254), .Y(n_280) );
INVx1_ASAP7_75t_L g297 ( .A(n_199), .Y(n_297) );
AND2x2_ASAP7_75t_L g303 ( .A(n_199), .B(n_218), .Y(n_303) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_203), .Y(n_478) );
INVx2_ASAP7_75t_L g506 ( .A(n_203), .Y(n_506) );
INVx1_ASAP7_75t_L g492 ( .A(n_205), .Y(n_492) );
AND2x2_ASAP7_75t_L g371 ( .A(n_206), .B(n_279), .Y(n_371) );
INVx2_ASAP7_75t_L g436 ( .A(n_206), .Y(n_436) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_218), .Y(n_206) );
AND2x2_ASAP7_75t_L g253 ( .A(n_207), .B(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g266 ( .A(n_207), .B(n_226), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_207), .B(n_225), .Y(n_294) );
INVx1_ASAP7_75t_L g300 ( .A(n_207), .Y(n_300) );
INVx1_ASAP7_75t_L g317 ( .A(n_207), .Y(n_317) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_207), .Y(n_329) );
INVx2_ASAP7_75t_L g397 ( .A(n_207), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g254 ( .A(n_218), .Y(n_254) );
BUFx2_ASAP7_75t_L g351 ( .A(n_218), .Y(n_351) );
AND2x2_ASAP7_75t_L g396 ( .A(n_218), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_237), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_224), .B(n_333), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_224), .A2(n_395), .B(n_409), .Y(n_419) );
AND2x2_ASAP7_75t_L g444 ( .A(n_224), .B(n_330), .Y(n_444) );
BUFx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g366 ( .A(n_226), .Y(n_366) );
AND2x2_ASAP7_75t_L g395 ( .A(n_226), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_227), .Y(n_279) );
INVx2_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_227), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_L g252 ( .A(n_238), .Y(n_252) );
OR2x2_ASAP7_75t_L g265 ( .A(n_238), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g333 ( .A(n_238), .B(n_329), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_238), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g434 ( .A(n_238), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_238), .B(n_371), .Y(n_446) );
AND2x2_ASAP7_75t_L g325 ( .A(n_239), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g348 ( .A(n_239), .B(n_241), .Y(n_348) );
INVx2_ASAP7_75t_L g260 ( .A(n_240), .Y(n_260) );
AND2x2_ASAP7_75t_L g288 ( .A(n_240), .B(n_261), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_240), .B(n_313), .Y(n_369) );
AND2x2_ASAP7_75t_L g283 ( .A(n_241), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g430 ( .A(n_241), .Y(n_430) );
AND2x2_ASAP7_75t_L g442 ( .A(n_241), .B(n_305), .Y(n_442) );
AND2x2_ASAP7_75t_L g268 ( .A(n_242), .B(n_258), .Y(n_268) );
INVx1_ASAP7_75t_L g363 ( .A(n_242), .Y(n_363) );
AO21x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_247), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_243), .B(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g498 ( .A(n_243), .Y(n_498) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_243), .A2(n_511), .B(n_518), .Y(n_510) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_243), .A2(n_567), .B(n_574), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_243), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g261 ( .A(n_248), .B(n_262), .Y(n_261) );
INVxp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_255), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_252), .B(n_299), .Y(n_308) );
OR2x2_ASAP7_75t_L g440 ( .A(n_252), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g357 ( .A(n_253), .B(n_298), .Y(n_357) );
AND2x2_ASAP7_75t_L g365 ( .A(n_253), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g424 ( .A(n_253), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g448 ( .A(n_253), .B(n_295), .Y(n_448) );
NOR2xp67_ASAP7_75t_L g406 ( .A(n_254), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g435 ( .A(n_254), .B(n_298), .Y(n_435) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2x1p5_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
AND2x2_ASAP7_75t_L g287 ( .A(n_257), .B(n_288), .Y(n_287) );
INVxp67_ASAP7_75t_L g449 ( .A(n_257), .Y(n_449) );
NOR2x1_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g284 ( .A(n_260), .Y(n_284) );
AND2x2_ASAP7_75t_L g335 ( .A(n_260), .B(n_268), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_260), .B(n_403), .Y(n_429) );
INVx2_ASAP7_75t_L g274 ( .A(n_261), .Y(n_274) );
INVx3_ASAP7_75t_L g326 ( .A(n_261), .Y(n_326) );
OR2x2_ASAP7_75t_L g354 ( .A(n_261), .B(n_355), .Y(n_354) );
AOI311xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_267), .A3(n_269), .B(n_270), .C(n_281), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g301 ( .A1(n_264), .A2(n_302), .B(n_304), .C(n_306), .Y(n_301) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_SL g286 ( .A(n_266), .Y(n_286) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g304 ( .A(n_268), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_268), .B(n_284), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_268), .B(n_269), .Y(n_437) );
AND2x2_ASAP7_75t_L g359 ( .A(n_269), .B(n_273), .Y(n_359) );
AOI21xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_275), .B(n_276), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g417 ( .A(n_273), .B(n_305), .Y(n_417) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_274), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g311 ( .A(n_274), .Y(n_311) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
AND2x2_ASAP7_75t_L g302 ( .A(n_278), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g347 ( .A(n_280), .Y(n_347) );
AND2x4_ASAP7_75t_L g409 ( .A(n_280), .B(n_378), .Y(n_409) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AOI222xp33_ASAP7_75t_L g360 ( .A1(n_283), .A2(n_349), .B1(n_361), .B2(n_365), .C1(n_367), .C2(n_371), .Y(n_360) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_289), .C(n_292), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_286), .B(n_330), .Y(n_353) );
INVx1_ASAP7_75t_L g375 ( .A(n_288), .Y(n_375) );
INVx1_ASAP7_75t_L g309 ( .A(n_290), .Y(n_309) );
OR2x2_ASAP7_75t_L g374 ( .A(n_291), .B(n_375), .Y(n_374) );
OAI21xp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_295), .B(n_299), .Y(n_292) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_293), .B(n_311), .C(n_312), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_293), .A2(n_330), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_297), .Y(n_350) );
AND2x2_ASAP7_75t_SL g316 ( .A(n_298), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g407 ( .A(n_298), .Y(n_407) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_298), .Y(n_423) );
INVx2_ASAP7_75t_L g381 ( .A(n_299), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_303), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g355 ( .A(n_305), .Y(n_355) );
OAI221xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B1(n_310), .B2(n_314), .C(n_315), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_309), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g443 ( .A(n_309), .Y(n_443) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g324 ( .A(n_316), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_316), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g382 ( .A(n_316), .B(n_330), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_316), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g415 ( .A(n_316), .B(n_350), .Y(n_415) );
BUFx3_ASAP7_75t_L g378 ( .A(n_317), .Y(n_378) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND5xp2_ASAP7_75t_L g320 ( .A(n_321), .B(n_339), .C(n_360), .D(n_372), .E(n_387), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI32xp33_ASAP7_75t_L g412 ( .A1(n_324), .A2(n_351), .A3(n_367), .B1(n_413), .B2(n_415), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_326), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g336 ( .A(n_330), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B1(n_336), .B2(n_337), .Y(n_331) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_346), .B1(n_348), .B2(n_349), .C(n_352), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g411 ( .A(n_343), .B(n_362), .Y(n_411) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_348), .A2(n_409), .B1(n_427), .B2(n_432), .C(n_433), .Y(n_426) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx2_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_356), .B2(n_358), .Y(n_352) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
INVx1_ASAP7_75t_L g370 ( .A(n_362), .Y(n_370) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
AOI222xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_376), .B1(n_380), .B2(n_381), .C1(n_382), .C2(n_383), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_381), .A2(n_428), .B1(n_430), .B2(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B(n_393), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI21xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_398), .B(n_400), .Y(n_393) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g441 ( .A(n_396), .Y(n_441) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
A2O1A1Ixp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_408), .B(n_410), .C(n_412), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B(n_420), .C(n_445), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g421 ( .A(n_417), .Y(n_421) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI211xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B(n_426), .C(n_438), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B(n_437), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_449), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g746 ( .A(n_458), .Y(n_746) );
OR3x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_658), .C(n_701), .Y(n_458) );
NAND5xp2_ASAP7_75t_L g459 ( .A(n_460), .B(n_585), .C(n_615), .D(n_632), .E(n_647), .Y(n_459) );
AOI221xp5_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_508), .B1(n_548), .B2(n_554), .C(n_558), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_483), .Y(n_461) );
OR2x2_ASAP7_75t_L g563 ( .A(n_462), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g602 ( .A(n_462), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g620 ( .A(n_462), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_462), .B(n_556), .Y(n_637) );
OR2x2_ASAP7_75t_L g649 ( .A(n_462), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_462), .B(n_608), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_462), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_462), .B(n_586), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_462), .B(n_594), .Y(n_700) );
AND2x2_ASAP7_75t_L g732 ( .A(n_462), .B(n_496), .Y(n_732) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_462), .Y(n_740) );
INVx5_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_463), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g560 ( .A(n_463), .B(n_538), .Y(n_560) );
BUFx2_ASAP7_75t_L g582 ( .A(n_463), .Y(n_582) );
AND2x2_ASAP7_75t_L g611 ( .A(n_463), .B(n_484), .Y(n_611) );
AND2x2_ASAP7_75t_L g666 ( .A(n_463), .B(n_564), .Y(n_666) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_481), .Y(n_463) );
BUFx2_ASAP7_75t_L g487 ( .A(n_466), .Y(n_487) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_SL g500 ( .A1(n_470), .A2(n_480), .B(n_501), .C(n_502), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_470), .A2(n_480), .B(n_543), .C(n_544), .Y(n_542) );
INVx5_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_477), .C(n_478), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_475), .A2(n_478), .B(n_535), .C(n_536), .Y(n_534) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_483), .B(n_620), .Y(n_629) );
OAI32xp33_ASAP7_75t_L g643 ( .A1(n_483), .A2(n_579), .A3(n_644), .B1(n_645), .B2(n_646), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_483), .B(n_645), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_483), .B(n_563), .Y(n_686) );
INVx1_ASAP7_75t_SL g715 ( .A(n_483), .Y(n_715) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_483), .B(n_510), .C(n_666), .D(n_725), .Y(n_724) );
AND2x4_ASAP7_75t_L g483 ( .A(n_484), .B(n_496), .Y(n_483) );
INVx5_ASAP7_75t_L g557 ( .A(n_484), .Y(n_557) );
AND2x2_ASAP7_75t_L g586 ( .A(n_484), .B(n_497), .Y(n_586) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_484), .Y(n_665) );
AND2x2_ASAP7_75t_L g735 ( .A(n_484), .B(n_682), .Y(n_735) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_493), .Y(n_484) );
AOI21xp5_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_488), .B(n_492), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
AND2x4_ASAP7_75t_L g608 ( .A(n_496), .B(n_557), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_496), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g642 ( .A(n_496), .B(n_564), .Y(n_642) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g556 ( .A(n_497), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g594 ( .A(n_497), .B(n_566), .Y(n_594) );
AND2x2_ASAP7_75t_L g603 ( .A(n_497), .B(n_565), .Y(n_603) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_507), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_508), .A2(n_672), .B1(n_674), .B2(n_676), .C1(n_679), .C2(n_680), .Y(n_671) );
AND2x4_ASAP7_75t_L g508 ( .A(n_509), .B(n_527), .Y(n_508) );
AND2x2_ASAP7_75t_L g604 ( .A(n_509), .B(n_605), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_509), .B(n_582), .C(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
INVx5_ASAP7_75t_SL g553 ( .A(n_510), .Y(n_553) );
OAI322xp33_ASAP7_75t_L g558 ( .A1(n_510), .A2(n_559), .A3(n_561), .B1(n_562), .B2(n_576), .C1(n_579), .C2(n_581), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_510), .B(n_551), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_510), .B(n_539), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_514), .Y(n_511) );
INVx2_ASAP7_75t_L g551 ( .A(n_520), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_520), .B(n_529), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_527), .B(n_589), .Y(n_644) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g623 ( .A(n_528), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .Y(n_528) );
OR2x2_ASAP7_75t_L g552 ( .A(n_529), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_529), .B(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g591 ( .A(n_529), .B(n_539), .Y(n_591) );
AND2x2_ASAP7_75t_L g614 ( .A(n_529), .B(n_551), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_529), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_529), .B(n_589), .Y(n_630) );
AND2x2_ASAP7_75t_L g638 ( .A(n_529), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_529), .B(n_598), .Y(n_688) );
INVx5_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g578 ( .A(n_530), .B(n_553), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_530), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g605 ( .A(n_530), .B(n_539), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_530), .B(n_652), .Y(n_693) );
OR2x2_ASAP7_75t_L g709 ( .A(n_530), .B(n_653), .Y(n_709) );
AND2x2_ASAP7_75t_SL g716 ( .A(n_530), .B(n_670), .Y(n_716) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_530), .Y(n_723) );
OR2x6_ASAP7_75t_L g530 ( .A(n_531), .B(n_537), .Y(n_530) );
AND2x2_ASAP7_75t_L g577 ( .A(n_538), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g627 ( .A(n_538), .B(n_551), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_538), .B(n_553), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_538), .B(n_589), .Y(n_711) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_539), .B(n_553), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_539), .B(n_551), .Y(n_599) );
OR2x2_ASAP7_75t_L g653 ( .A(n_539), .B(n_551), .Y(n_653) );
AND2x2_ASAP7_75t_L g670 ( .A(n_539), .B(n_550), .Y(n_670) );
INVxp67_ASAP7_75t_L g692 ( .A(n_539), .Y(n_692) );
AND2x2_ASAP7_75t_L g719 ( .A(n_539), .B(n_589), .Y(n_719) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_539), .Y(n_726) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B(n_547), .Y(n_539) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_550), .B(n_600), .Y(n_673) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g589 ( .A(n_551), .B(n_553), .Y(n_589) );
OR2x2_ASAP7_75t_L g656 ( .A(n_551), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g600 ( .A(n_552), .Y(n_600) );
OR2x2_ASAP7_75t_L g661 ( .A(n_552), .B(n_653), .Y(n_661) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g561 ( .A(n_556), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_556), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g562 ( .A(n_557), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_557), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_557), .B(n_564), .Y(n_596) );
INVx2_ASAP7_75t_L g641 ( .A(n_557), .Y(n_641) );
AND2x2_ASAP7_75t_L g654 ( .A(n_557), .B(n_594), .Y(n_654) );
AND2x2_ASAP7_75t_L g679 ( .A(n_557), .B(n_603), .Y(n_679) );
INVx1_ASAP7_75t_L g631 ( .A(n_562), .Y(n_631) );
INVx2_ASAP7_75t_SL g618 ( .A(n_563), .Y(n_618) );
INVx1_ASAP7_75t_L g621 ( .A(n_564), .Y(n_621) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_565), .Y(n_584) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g682 ( .A(n_566), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_573), .Y(n_567) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g651 ( .A(n_578), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g657 ( .A(n_578), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_578), .A2(n_660), .B1(n_662), .B2(n_667), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_578), .B(n_670), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_579), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g613 ( .A(n_580), .Y(n_613) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
OR2x2_ASAP7_75t_L g595 ( .A(n_582), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_582), .B(n_586), .Y(n_646) );
AND2x2_ASAP7_75t_L g669 ( .A(n_582), .B(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g645 ( .A(n_584), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_592), .C(n_606), .Y(n_585) );
INVx1_ASAP7_75t_L g609 ( .A(n_586), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g717 ( .A1(n_586), .A2(n_718), .B1(n_720), .B2(n_721), .C(n_724), .Y(n_717) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g736 ( .A(n_589), .Y(n_736) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g685 ( .A(n_591), .B(n_624), .Y(n_685) );
A2O1A1Ixp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B(n_597), .C(n_601), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
OAI32xp33_ASAP7_75t_L g710 ( .A1(n_599), .A2(n_600), .A3(n_663), .B1(n_700), .B2(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
AND2x2_ASAP7_75t_L g742 ( .A(n_602), .B(n_641), .Y(n_742) );
AND2x2_ASAP7_75t_L g689 ( .A(n_603), .B(n_641), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_603), .B(n_611), .Y(n_707) );
AOI31xp33_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_609), .A3(n_610), .B(n_612), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_608), .B(n_620), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_608), .B(n_618), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_608), .A2(n_638), .B1(n_728), .B2(n_731), .C(n_733), .Y(n_727) );
CKINVDCx16_ASAP7_75t_R g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g633 ( .A(n_613), .B(n_634), .Y(n_633) );
AOI222xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_622), .B1(n_625), .B2(n_628), .C1(n_630), .C2(n_631), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g698 ( .A(n_617), .Y(n_698) );
INVx1_ASAP7_75t_L g720 ( .A(n_620), .Y(n_720) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_623), .A2(n_734), .B1(n_736), .B2(n_737), .Y(n_733) );
INVx1_ASAP7_75t_L g639 ( .A(n_624), .Y(n_639) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .B1(n_638), .B2(n_640), .C(n_643), .Y(n_632) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g677 ( .A(n_635), .B(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g729 ( .A(n_635), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g704 ( .A(n_640), .Y(n_704) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g668 ( .A(n_641), .Y(n_668) );
INVx1_ASAP7_75t_L g650 ( .A(n_642), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_645), .B(n_732), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B1(n_654), .B2(n_655), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g741 ( .A(n_654), .Y(n_741) );
INVxp33_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_656), .B(n_700), .Y(n_699) );
OAI32xp33_ASAP7_75t_L g690 ( .A1(n_657), .A2(n_691), .A3(n_692), .B1(n_693), .B2(n_694), .Y(n_690) );
NAND4xp25_ASAP7_75t_L g658 ( .A(n_659), .B(n_671), .C(n_683), .D(n_695), .Y(n_658) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
NAND2xp33_ASAP7_75t_SL g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_666), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
CKINVDCx16_ASAP7_75t_R g676 ( .A(n_677), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_680), .A2(n_696), .B1(n_713), .B2(n_716), .C(n_717), .Y(n_712) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g731 ( .A(n_682), .B(n_732), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B1(n_687), .B2(n_689), .C(n_690), .Y(n_683) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_692), .B(n_723), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g701 ( .A(n_702), .B(n_712), .C(n_727), .D(n_738), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_706), .B(n_708), .C(n_710), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g743 ( .A(n_730), .Y(n_743) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OAI21xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_742), .B(n_743), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
endmodule