module fake_netlist_6_2104_n_72 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_72);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_72;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_70;
wire n_18;
wire n_21;
wire n_24;
wire n_71;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_69;
wire n_20;
wire n_50;
wire n_64;
wire n_30;
wire n_49;
wire n_43;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_65;
wire n_31;
wire n_48;
wire n_25;
wire n_40;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_2),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_0),
.A2(n_1),
.B1(n_15),
.B2(n_8),
.Y(n_21)
);

AND2x4_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_17),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_1),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_2),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_16),
.C(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_21),
.B1(n_20),
.B2(n_26),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_21),
.B1(n_20),
.B2(n_29),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_23),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_19),
.B(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

AO21x1_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_22),
.B(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_31),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_30),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_52),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_44),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVxp67_ASAP7_75t_SL g60 ( 
.A(n_56),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_54),
.B(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_59),
.B(n_57),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_61),
.B(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_62),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

AND3x2_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_49),
.C(n_48),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_67),
.B1(n_59),
.B2(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_59),
.B1(n_18),
.B2(n_23),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_69),
.B1(n_18),
.B2(n_45),
.Y(n_71)
);

OR2x6_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_45),
.Y(n_72)
);


endmodule