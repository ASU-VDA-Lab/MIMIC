module fake_jpeg_1082_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_12),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_41),
.Y(n_107)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_45),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_23),
.A2(n_6),
.B(n_13),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_18),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_62),
.Y(n_90)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_13),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_14),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

CKINVDCx6p67_ASAP7_75t_R g102 ( 
.A(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_14),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_18),
.B1(n_38),
.B2(n_39),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_74),
.A2(n_93),
.B1(n_101),
.B2(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_30),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_34),
.B1(n_19),
.B2(n_28),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_95),
.B1(n_34),
.B2(n_28),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_22),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_22),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_84),
.Y(n_132)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_43),
.A2(n_24),
.B(n_27),
.C(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_100),
.Y(n_113)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_39),
.B1(n_24),
.B2(n_19),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_35),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_96),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_57),
.A2(n_60),
.B1(n_58),
.B2(n_34),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_8),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_45),
.A2(n_24),
.B(n_27),
.C(n_31),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_39),
.B1(n_21),
.B2(n_32),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_41),
.A2(n_34),
.B1(n_36),
.B2(n_28),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g105 ( 
.A(n_62),
.B(n_36),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_20),
.Y(n_110)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_36),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_117),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_131),
.C(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_114),
.A2(n_118),
.B1(n_134),
.B2(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_20),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_35),
.B1(n_32),
.B2(n_31),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

AO22x1_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_33),
.B1(n_37),
.B2(n_25),
.Y(n_122)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_0),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_124),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_126),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_0),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_71),
.B(n_33),
.C(n_37),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_73),
.C(n_87),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_80),
.A2(n_33),
.B1(n_25),
.B2(n_37),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_72),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_33),
.B1(n_25),
.B2(n_3),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_141),
.B1(n_98),
.B2(n_2),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_33),
.B1(n_2),
.B2(n_3),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_104),
.B(n_11),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_143),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_93),
.A2(n_33),
.B1(n_11),
.B2(n_10),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_70),
.C(n_69),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_156),
.C(n_158),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_160),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_120),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_103),
.B(n_92),
.C(n_97),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_153),
.A2(n_178),
.B(n_115),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_73),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_154),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_76),
.C(n_87),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_109),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_85),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_85),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_8),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_170),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_70),
.B1(n_69),
.B2(n_68),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_173),
.B1(n_134),
.B2(n_114),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_113),
.A2(n_88),
.B1(n_68),
.B2(n_98),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_174),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_72),
.C(n_88),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_116),
.C(n_5),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_126),
.A2(n_8),
.B(n_3),
.C(n_4),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_122),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_177),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_122),
.A2(n_1),
.B(n_4),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_179),
.B(n_209),
.Y(n_218)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_166),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_199),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_210),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_144),
.B1(n_118),
.B2(n_142),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_192),
.B1(n_202),
.B2(n_161),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_112),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_190),
.Y(n_223)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_112),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_123),
.B1(n_130),
.B2(n_128),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_127),
.B1(n_135),
.B2(n_137),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_194),
.A2(n_152),
.B1(n_161),
.B2(n_169),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_201),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_131),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_203),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_198),
.A2(n_154),
.B(n_170),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_4),
.A3(n_5),
.B1(n_138),
.B2(n_121),
.C1(n_116),
.C2(n_72),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_5),
.B1(n_171),
.B2(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_5),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_149),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_177),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_148),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_205),
.B(n_145),
.Y(n_214)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_154),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_208),
.B(n_156),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_147),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_153),
.B1(n_178),
.B2(n_152),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_226),
.B(n_231),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_224),
.B1(n_230),
.B2(n_197),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_235),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_195),
.C(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_159),
.B(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_184),
.B(n_165),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_233),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_165),
.B1(n_151),
.B2(n_160),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_147),
.B(n_177),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_187),
.A2(n_151),
.B(n_162),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_234),
.B(n_218),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_185),
.Y(n_235)
);

AOI322xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_193),
.A3(n_190),
.B1(n_179),
.B2(n_204),
.C1(n_181),
.C2(n_196),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_241),
.A3(n_222),
.B1(n_189),
.B2(n_225),
.C1(n_212),
.C2(n_216),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_217),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_SL g241 ( 
.A(n_215),
.B(n_200),
.C(n_208),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_181),
.A3(n_200),
.B1(n_186),
.B2(n_210),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_221),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_211),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_248),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_250),
.C(n_212),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_183),
.B1(n_210),
.B2(n_209),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_230),
.B1(n_223),
.B2(n_227),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_201),
.C(n_207),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_235),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_251),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_231),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_252),
.A2(n_234),
.B1(n_215),
.B2(n_233),
.Y(n_258)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_219),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_260),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_262),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_268),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_223),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_247),
.B1(n_240),
.B2(n_244),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_244),
.B(n_226),
.CI(n_232),
.CON(n_262),
.SN(n_262)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_232),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_248),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_256),
.C(n_259),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_276),
.C(n_277),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_281),
.B1(n_253),
.B2(n_243),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_279),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_252),
.C(n_237),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_237),
.C(n_249),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_269),
.A2(n_254),
.B1(n_239),
.B2(n_242),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_238),
.C(n_262),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_263),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_264),
.B1(n_261),
.B2(n_254),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_284),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_273),
.A2(n_264),
.B1(n_257),
.B2(n_262),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_276),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_255),
.C(n_228),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_289),
.Y(n_295)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_189),
.B1(n_224),
.B2(n_243),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_294),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_285),
.Y(n_294)
);

AOI31xp67_ASAP7_75t_SL g296 ( 
.A1(n_286),
.A2(n_271),
.A3(n_280),
.B(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_296),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_290),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_300),
.B(n_283),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_283),
.B(n_284),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_302),
.C(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_293),
.C(n_292),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_303),
.A2(n_304),
.B(n_270),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_282),
.B(n_278),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_278),
.Y(n_307)
);


endmodule