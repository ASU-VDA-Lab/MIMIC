module fake_netlist_1_7713_n_746 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_746);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_746;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_33), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_7), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_62), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_21), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_45), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_66), .Y(n_86) );
INVxp33_ASAP7_75t_L g87 ( .A(n_75), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
INVx2_ASAP7_75t_SL g89 ( .A(n_59), .Y(n_89) );
BUFx5_ASAP7_75t_L g90 ( .A(n_13), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_11), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_67), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_76), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_34), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_26), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_42), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_44), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_8), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_17), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_15), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_37), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_20), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_12), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_41), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_32), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_54), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_16), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_65), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_18), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_9), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_6), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_64), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_27), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_18), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_7), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_68), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_43), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_51), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_3), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_25), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_28), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_17), .Y(n_122) );
INVx2_ASAP7_75t_SL g123 ( .A(n_4), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_61), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_80), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_5), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_30), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_12), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_13), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_16), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_47), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_131), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_131), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_90), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_90), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_131), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_90), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_114), .B(n_0), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_131), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_90), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_122), .B(n_0), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_99), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
NAND2xp33_ASAP7_75t_SL g145 ( .A(n_87), .B(n_1), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_99), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_90), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_131), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_90), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_107), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_85), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_85), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_104), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_86), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_107), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_104), .Y(n_156) );
BUFx12f_ASAP7_75t_L g157 ( .A(n_81), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_105), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_105), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_107), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_111), .B(n_1), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_123), .B(n_2), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_107), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_89), .B(n_2), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_86), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_93), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_107), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_118), .Y(n_168) );
NAND2xp33_ASAP7_75t_SL g169 ( .A(n_123), .B(n_3), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_118), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_95), .Y(n_171) );
NAND2x1_ASAP7_75t_L g172 ( .A(n_91), .B(n_4), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_127), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_89), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_91), .B(n_5), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_98), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_127), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_174), .B(n_98), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_162), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_175), .B(n_95), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_170), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_143), .B(n_81), .Y(n_183) );
INVx4_ASAP7_75t_SL g184 ( .A(n_174), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_170), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_170), .Y(n_186) );
NAND2xp33_ASAP7_75t_SL g187 ( .A(n_161), .B(n_97), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_143), .B(n_100), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_170), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_174), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_175), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_151), .B(n_152), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_146), .B(n_100), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_176), .B(n_130), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_151), .B(n_108), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_132), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_132), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_140), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_152), .B(n_83), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_154), .B(n_130), .Y(n_200) );
INVx2_ASAP7_75t_SL g201 ( .A(n_157), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_154), .B(n_88), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_132), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_161), .B(n_166), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_140), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_165), .B(n_102), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_165), .B(n_106), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_171), .B(n_129), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_157), .B(n_97), .Y(n_210) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_164), .B(n_112), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_170), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_157), .B(n_101), .Y(n_213) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_171), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_138), .B(n_128), .C(n_126), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_140), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_177), .B(n_113), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_170), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_134), .Y(n_219) );
OR2x2_ASAP7_75t_L g220 ( .A(n_142), .B(n_115), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_134), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_145), .A2(n_103), .B1(n_82), .B2(n_109), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_132), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_153), .B(n_101), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_160), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_160), .Y(n_226) );
BUFx4f_ASAP7_75t_L g227 ( .A(n_135), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_177), .B(n_116), .Y(n_228) );
INVxp67_ASAP7_75t_SL g229 ( .A(n_153), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_160), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_169), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_153), .B(n_117), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_135), .Y(n_233) );
INVx1_ASAP7_75t_SL g234 ( .A(n_156), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_172), .A2(n_103), .B1(n_110), .B2(n_119), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_156), .B(n_120), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_156), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_160), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_137), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_132), .Y(n_240) );
BUFx8_ASAP7_75t_SL g241 ( .A(n_158), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_137), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_160), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_158), .B(n_125), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_141), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_158), .B(n_125), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_172), .B(n_112), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_180), .B(n_84), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_214), .B(n_147), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_214), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_229), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_181), .A2(n_147), .B1(n_141), .B2(n_144), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_181), .A2(n_144), .B1(n_149), .B2(n_168), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_194), .B(n_177), .Y(n_255) );
NAND2x1p5_ASAP7_75t_L g256 ( .A(n_200), .B(n_96), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_194), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_218), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_224), .B(n_194), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_190), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_182), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_182), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_179), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_181), .A2(n_149), .B1(n_168), .B2(n_173), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_218), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_234), .B(n_173), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_190), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_192), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_200), .Y(n_269) );
INVx2_ASAP7_75t_SL g270 ( .A(n_200), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_181), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_185), .Y(n_272) );
INVx6_ASAP7_75t_L g273 ( .A(n_184), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_179), .Y(n_274) );
INVx5_ASAP7_75t_L g275 ( .A(n_198), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_241), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_185), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_237), .B(n_173), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_188), .B(n_159), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_216), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_181), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_246), .Y(n_282) );
INVx5_ASAP7_75t_L g283 ( .A(n_198), .Y(n_283) );
NAND3xp33_ASAP7_75t_SL g284 ( .A(n_222), .B(n_121), .C(n_124), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_193), .A2(n_92), .B1(n_94), .B2(n_159), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_241), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_195), .B(n_168), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_246), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_195), .B(n_159), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_216), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_179), .Y(n_291) );
BUFx8_ASAP7_75t_L g292 ( .A(n_201), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_244), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_183), .B(n_96), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_209), .B(n_150), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_186), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_211), .A2(n_150), .B1(n_155), .B2(n_133), .Y(n_297) );
BUFx12f_ASAP7_75t_L g298 ( .A(n_188), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_186), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_187), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_231), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_193), .B(n_150), .Y(n_302) );
BUFx4f_ASAP7_75t_L g303 ( .A(n_247), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_189), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_187), .B(n_6), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_228), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_232), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_191), .B(n_150), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_189), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_210), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_199), .A2(n_155), .B(n_133), .C(n_148), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_220), .B(n_8), .Y(n_312) );
AND2x4_ASAP7_75t_SL g313 ( .A(n_213), .B(n_155), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_209), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_205), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_209), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_235), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_247), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_211), .B(n_155), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_247), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_202), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_212), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_298), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_275), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_275), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_321), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_275), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_249), .A2(n_227), .B(n_206), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_SL g329 ( .A1(n_311), .A2(n_212), .B(n_217), .C(n_236), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_268), .B(n_199), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_268), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_291), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_275), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_291), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_292), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_275), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_321), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_283), .Y(n_339) );
HAxp5_ASAP7_75t_L g340 ( .A(n_317), .B(n_215), .CON(n_340), .SN(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_292), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_291), .Y(n_342) );
INVx4_ASAP7_75t_L g343 ( .A(n_283), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_266), .A2(n_227), .B(n_245), .Y(n_344) );
INVx6_ASAP7_75t_L g345 ( .A(n_292), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_263), .Y(n_346) );
INVx5_ASAP7_75t_SL g347 ( .A(n_255), .Y(n_347) );
AO31x2_ASAP7_75t_L g348 ( .A1(n_294), .A2(n_236), .A3(n_217), .B(n_203), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_306), .A2(n_207), .B(n_208), .C(n_203), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_274), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_316), .A2(n_207), .B1(n_208), .B2(n_239), .Y(n_351) );
NOR2xp33_ASAP7_75t_SL g352 ( .A(n_303), .B(n_242), .Y(n_352) );
AO22x1_ASAP7_75t_L g353 ( .A1(n_286), .A2(n_184), .B1(n_10), .B2(n_11), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_306), .B(n_184), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_283), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_283), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_283), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_320), .B(n_219), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_269), .Y(n_359) );
CKINVDCx11_ASAP7_75t_R g360 ( .A(n_315), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_321), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_258), .Y(n_362) );
BUFx4f_ASAP7_75t_SL g363 ( .A(n_300), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_258), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_286), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_258), .Y(n_366) );
AOI21xp33_ASAP7_75t_L g367 ( .A1(n_257), .A2(n_233), .B(n_221), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_269), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_312), .B(n_9), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_307), .B(n_10), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_278), .A2(n_226), .B(n_225), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_280), .A2(n_226), .B(n_225), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_257), .A2(n_133), .B1(n_136), .B2(n_148), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_270), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_307), .B(n_14), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_258), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g377 ( .A1(n_259), .A2(n_136), .B1(n_139), .B2(n_148), .C(n_167), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_270), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_312), .B(n_14), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_258), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_336), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_326), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_331), .B(n_318), .Y(n_383) );
OR2x6_ASAP7_75t_L g384 ( .A(n_345), .B(n_271), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_360), .A2(n_317), .B1(n_300), .B2(n_310), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_379), .A2(n_284), .B1(n_256), .B2(n_314), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_330), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_379), .A2(n_256), .B1(n_314), .B2(n_303), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_345), .A2(n_276), .B1(n_303), .B2(n_305), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_346), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_344), .A2(n_280), .B(n_290), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_360), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_350), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_326), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_338), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_341), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_369), .B(n_255), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_338), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_339), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_339), .Y(n_400) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_324), .B(n_334), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_349), .B(n_255), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_363), .A2(n_305), .B1(n_319), .B2(n_301), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_361), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_363), .A2(n_319), .B1(n_301), .B2(n_250), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_351), .A2(n_256), .B1(n_271), .B2(n_281), .Y(n_407) );
AND2x6_ASAP7_75t_L g408 ( .A(n_347), .B(n_281), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_349), .B(n_293), .Y(n_409) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_324), .B(n_318), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_358), .A2(n_320), .B1(n_318), .B2(n_254), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_365), .A2(n_248), .B1(n_279), .B2(n_293), .C(n_285), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_348), .B(n_279), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_370), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_339), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_347), .B(n_282), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_386), .A2(n_345), .B1(n_352), .B2(n_365), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_386), .A2(n_388), .B1(n_387), .B2(n_403), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_392), .A2(n_375), .B1(n_333), .B2(n_378), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_387), .A2(n_358), .B1(n_347), .B2(n_378), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_382), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_413), .A2(n_358), .B1(n_288), .B2(n_282), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_392), .A2(n_359), .B1(n_374), .B2(n_368), .Y(n_423) );
OAI21xp5_ASAP7_75t_L g424 ( .A1(n_414), .A2(n_367), .B(n_297), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_413), .B(n_348), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_404), .A2(n_288), .B1(n_282), .B2(n_264), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_412), .B(n_348), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_390), .Y(n_428) );
OAI22xp33_ASAP7_75t_L g429 ( .A1(n_384), .A2(n_288), .B1(n_334), .B2(n_343), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_409), .B(n_348), .Y(n_430) );
AOI222xp33_ASAP7_75t_L g431 ( .A1(n_409), .A2(n_353), .B1(n_302), .B2(n_308), .C1(n_340), .C2(n_289), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g432 ( .A1(n_384), .A2(n_343), .B1(n_334), .B2(n_324), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_414), .A2(n_354), .B1(n_313), .B2(n_335), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_389), .A2(n_323), .B1(n_354), .B2(n_356), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_390), .B(n_287), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_393), .A2(n_391), .B(n_328), .C(n_397), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_393), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_385), .A2(n_308), .B1(n_329), .B2(n_332), .C(n_342), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_397), .A2(n_383), .B1(n_381), .B2(n_406), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_396), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_382), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_383), .A2(n_313), .B1(n_343), .B2(n_325), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_410), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_394), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_383), .A2(n_329), .B1(n_340), .B2(n_251), .C(n_377), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_421), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_425), .B(n_398), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_431), .A2(n_383), .B1(n_402), .B2(n_411), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_418), .A2(n_407), .B1(n_402), .B2(n_401), .Y(n_450) );
OAI211xp5_ASAP7_75t_SL g451 ( .A1(n_439), .A2(n_416), .B(n_295), .C(n_373), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_425), .B(n_399), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_421), .Y(n_453) );
INVx5_ASAP7_75t_L g454 ( .A(n_444), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_428), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_428), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_427), .B(n_394), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_443), .B(n_399), .Y(n_458) );
OAI222xp33_ASAP7_75t_L g459 ( .A1(n_434), .A2(n_384), .B1(n_410), .B2(n_400), .C1(n_415), .C2(n_395), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_437), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_430), .B(n_400), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_430), .B(n_395), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_441), .B(n_405), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_441), .B(n_405), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_444), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_445), .B(n_415), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_419), .A2(n_253), .B1(n_252), .B2(n_290), .C(n_136), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_436), .A2(n_401), .B(n_362), .Y(n_468) );
INVx4_ASAP7_75t_L g469 ( .A(n_444), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_445), .B(n_410), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_437), .Y(n_471) );
OAI31xp33_ASAP7_75t_L g472 ( .A1(n_417), .A2(n_325), .A3(n_355), .B(n_337), .Y(n_472) );
AOI33xp33_ASAP7_75t_L g473 ( .A1(n_423), .A2(n_139), .A3(n_230), .B1(n_238), .B2(n_15), .B3(n_19), .Y(n_473) );
OAI221xp5_ASAP7_75t_SL g474 ( .A1(n_435), .A2(n_384), .B1(n_327), .B2(n_356), .C(n_337), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_435), .B(n_366), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_424), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_426), .A2(n_384), .B1(n_408), .B2(n_327), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_422), .A2(n_139), .B1(n_357), .B2(n_167), .C(n_163), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_438), .A2(n_408), .B1(n_357), .B2(n_339), .Y(n_481) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_436), .A2(n_371), .B(n_380), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_429), .Y(n_483) );
OAI33xp33_ASAP7_75t_L g484 ( .A1(n_446), .A2(n_19), .A3(n_380), .B1(n_376), .B2(n_366), .B3(n_238), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_448), .B(n_440), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_448), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_451), .A2(n_433), .B1(n_442), .B2(n_163), .C(n_167), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_452), .B(n_376), .Y(n_488) );
NAND4xp25_ASAP7_75t_L g489 ( .A(n_449), .B(n_372), .C(n_355), .D(n_357), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_451), .A2(n_160), .B1(n_163), .B2(n_167), .C(n_267), .Y(n_490) );
OAI33xp33_ASAP7_75t_L g491 ( .A1(n_455), .A2(n_230), .A3(n_163), .B1(n_167), .B2(n_296), .B3(n_277), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_471), .Y(n_492) );
AOI211xp5_ASAP7_75t_SL g493 ( .A1(n_474), .A2(n_267), .B(n_408), .C(n_24), .Y(n_493) );
BUFx3_ASAP7_75t_L g494 ( .A(n_454), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_447), .Y(n_495) );
OAI211xp5_ASAP7_75t_L g496 ( .A1(n_475), .A2(n_163), .B(n_167), .C(n_267), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_475), .A2(n_408), .B1(n_364), .B2(n_362), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_452), .B(n_364), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_447), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_447), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_478), .A2(n_408), .B1(n_364), .B2(n_362), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_471), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_462), .B(n_364), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_462), .B(n_362), .Y(n_504) );
OAI31xp33_ASAP7_75t_L g505 ( .A1(n_474), .A2(n_260), .A3(n_408), .B(n_304), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_453), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_476), .B(n_455), .Y(n_508) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_473), .B(n_163), .C(n_243), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_456), .B(n_408), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_461), .B(n_260), .Y(n_511) );
INVx5_ASAP7_75t_L g512 ( .A(n_469), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_469), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_476), .B(n_265), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g515 ( .A(n_484), .B(n_322), .C(n_304), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_471), .B(n_22), .Y(n_516) );
OAI31xp33_ASAP7_75t_L g517 ( .A1(n_459), .A2(n_450), .A3(n_472), .B(n_478), .Y(n_517) );
OAI33xp33_ASAP7_75t_L g518 ( .A1(n_456), .A2(n_322), .A3(n_299), .B1(n_296), .B2(n_277), .B3(n_262), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_460), .B(n_23), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_461), .B(n_29), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_460), .Y(n_521) );
OAI31xp33_ASAP7_75t_SL g522 ( .A1(n_450), .A2(n_31), .A3(n_36), .B(n_38), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_458), .B(n_265), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_463), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_469), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_463), .B(n_464), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_464), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_457), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_457), .B(n_39), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_454), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_470), .B(n_40), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_469), .B(n_46), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_470), .B(n_48), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_477), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_472), .B(n_243), .C(n_178), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g536 ( .A1(n_449), .A2(n_273), .B1(n_50), .B2(n_52), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_466), .B(n_49), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_477), .Y(n_538) );
NAND2xp67_ASAP7_75t_L g539 ( .A(n_485), .B(n_458), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_517), .B(n_480), .C(n_468), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_526), .B(n_466), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_486), .B(n_477), .Y(n_542) );
INVxp67_ASAP7_75t_SL g543 ( .A(n_506), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_521), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_508), .B(n_454), .Y(n_545) );
INVxp67_ASAP7_75t_L g546 ( .A(n_525), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_507), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_526), .B(n_483), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_492), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_507), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_524), .B(n_483), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_492), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_517), .A2(n_484), .B1(n_481), .B2(n_479), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_527), .B(n_465), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_535), .A2(n_468), .B(n_459), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_527), .B(n_465), .Y(n_556) );
INVxp67_ASAP7_75t_SL g557 ( .A(n_495), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_502), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_525), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_512), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_528), .B(n_465), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_502), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_528), .B(n_488), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_488), .B(n_465), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_495), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_498), .B(n_454), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_498), .B(n_454), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_520), .B(n_454), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_499), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_512), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_512), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_509), .A2(n_467), .B1(n_480), .B2(n_479), .C(n_482), .Y(n_572) );
OAI33xp33_ASAP7_75t_L g573 ( .A1(n_536), .A2(n_482), .A3(n_454), .B1(n_467), .B2(n_56), .B3(n_57), .Y(n_573) );
AND2x2_ASAP7_75t_SL g574 ( .A(n_522), .B(n_482), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_499), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_503), .B(n_482), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_511), .B(n_53), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_504), .B(n_55), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_512), .B(n_58), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_509), .B(n_243), .C(n_223), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_500), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_512), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_512), .B(n_265), .Y(n_583) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_535), .B(n_243), .Y(n_584) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_513), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_534), .Y(n_586) );
AND2x2_ASAP7_75t_SL g587 ( .A(n_532), .B(n_60), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_504), .B(n_63), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_534), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_511), .B(n_69), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_520), .B(n_70), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_523), .B(n_71), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_538), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g594 ( .A1(n_493), .A2(n_261), .B(n_262), .C(n_299), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_504), .B(n_72), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_538), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_489), .B(n_73), .Y(n_597) );
NAND4xp25_ASAP7_75t_L g598 ( .A(n_487), .B(n_261), .C(n_77), .D(n_78), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_541), .B(n_513), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_539), .B(n_536), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_576), .B(n_504), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_543), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_548), .B(n_543), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_547), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_553), .B(n_505), .C(n_510), .Y(n_605) );
XOR2xp5_ASAP7_75t_L g606 ( .A(n_582), .B(n_533), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_557), .B(n_513), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_551), .B(n_530), .Y(n_608) );
AOI211xp5_ASAP7_75t_L g609 ( .A1(n_540), .A2(n_505), .B(n_532), .C(n_496), .Y(n_609) );
INVx2_ASAP7_75t_SL g610 ( .A(n_560), .Y(n_610) );
NAND2xp33_ASAP7_75t_SL g611 ( .A(n_571), .B(n_530), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_549), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_557), .B(n_516), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_570), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_563), .B(n_519), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_552), .Y(n_616) );
INVx2_ASAP7_75t_SL g617 ( .A(n_585), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_562), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_558), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_544), .B(n_516), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_550), .B(n_519), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_586), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_567), .B(n_494), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_553), .B(n_490), .C(n_501), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_542), .B(n_514), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g626 ( .A(n_597), .B(n_497), .C(n_529), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_589), .Y(n_627) );
OAI31xp33_ASAP7_75t_SL g628 ( .A1(n_584), .A2(n_532), .A3(n_533), .B(n_531), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_587), .A2(n_491), .B(n_518), .Y(n_629) );
INVxp67_ASAP7_75t_L g630 ( .A(n_585), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_561), .B(n_529), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_546), .B(n_537), .Y(n_632) );
OAI21x1_ASAP7_75t_SL g633 ( .A1(n_555), .A2(n_494), .B(n_532), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_565), .B(n_531), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_593), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_569), .B(n_537), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_596), .B(n_515), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_554), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_575), .B(n_74), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_546), .B(n_79), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_559), .B(n_178), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g642 ( .A1(n_597), .A2(n_178), .B(n_196), .C(n_197), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_587), .A2(n_273), .B1(n_265), .B2(n_197), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_556), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_559), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_581), .B(n_178), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_564), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_566), .B(n_545), .Y(n_648) );
AND2x2_ASAP7_75t_SL g649 ( .A(n_574), .B(n_196), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_568), .B(n_196), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_579), .Y(n_651) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_643), .B(n_579), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_603), .B(n_577), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_649), .B(n_574), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_602), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_638), .B(n_572), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_612), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_601), .B(n_555), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_644), .B(n_578), .Y(n_659) );
XOR2x2_ASAP7_75t_L g660 ( .A(n_606), .B(n_591), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_616), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_611), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_600), .A2(n_590), .B1(n_598), .B2(n_594), .C(n_592), .Y(n_663) );
AOI21xp33_ASAP7_75t_L g664 ( .A1(n_600), .A2(n_594), .B(n_595), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_599), .B(n_583), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_647), .B(n_588), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_623), .B(n_580), .Y(n_667) );
XNOR2xp5_ASAP7_75t_L g668 ( .A(n_648), .B(n_573), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_628), .A2(n_573), .B(n_265), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_604), .B(n_196), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_645), .B(n_197), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_618), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_605), .A2(n_197), .B1(n_204), .B2(n_223), .C(n_240), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_622), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_627), .Y(n_675) );
INVxp67_ASAP7_75t_L g676 ( .A(n_604), .Y(n_676) );
AOI222xp33_ASAP7_75t_L g677 ( .A1(n_649), .A2(n_204), .B1(n_223), .B2(n_240), .C1(n_273), .C2(n_272), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_610), .B(n_204), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_611), .Y(n_679) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_624), .A2(n_223), .B1(n_240), .B2(n_273), .C1(n_272), .C2(n_309), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_626), .A2(n_240), .B1(n_272), .B2(n_309), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_635), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_625), .B(n_272), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g684 ( .A1(n_637), .A2(n_309), .B(n_633), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_607), .B(n_309), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_617), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_608), .B(n_309), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_609), .A2(n_630), .B1(n_632), .B2(n_617), .C(n_651), .Y(n_688) );
AOI211xp5_ASAP7_75t_SL g689 ( .A1(n_632), .A2(n_642), .B(n_629), .C(n_607), .Y(n_689) );
OAI221xp5_ASAP7_75t_SL g690 ( .A1(n_615), .A2(n_634), .B1(n_636), .B2(n_651), .C(n_631), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_636), .B(n_634), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_619), .Y(n_692) );
BUFx2_ASAP7_75t_L g693 ( .A(n_614), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_620), .B(n_613), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_620), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_621), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_613), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_640), .B(n_621), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_641), .Y(n_699) );
INVxp67_ASAP7_75t_L g700 ( .A(n_646), .Y(n_700) );
INVx2_ASAP7_75t_SL g701 ( .A(n_650), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_639), .A2(n_628), .B(n_649), .Y(n_702) );
INVxp67_ASAP7_75t_L g703 ( .A(n_604), .Y(n_703) );
OAI21xp5_ASAP7_75t_L g704 ( .A1(n_649), .A2(n_587), .B(n_605), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_628), .B(n_602), .C(n_609), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_602), .Y(n_706) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_643), .B(n_584), .Y(n_707) );
OAI322xp33_ASAP7_75t_L g708 ( .A1(n_688), .A2(n_705), .A3(n_656), .B1(n_668), .B2(n_703), .C1(n_676), .C2(n_654), .Y(n_708) );
OAI31xp33_ASAP7_75t_L g709 ( .A1(n_679), .A2(n_654), .A3(n_702), .B(n_689), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_704), .B(n_669), .C(n_703), .Y(n_710) );
OAI21xp33_ASAP7_75t_L g711 ( .A1(n_658), .A2(n_690), .B(n_660), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_664), .A2(n_663), .B(n_676), .C(n_693), .Y(n_712) );
AND2x4_ASAP7_75t_L g713 ( .A(n_662), .B(n_652), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_655), .B(n_706), .Y(n_714) );
OAI211xp5_ASAP7_75t_SL g715 ( .A1(n_686), .A2(n_680), .B(n_684), .C(n_707), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_682), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_670), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_662), .A2(n_660), .B(n_673), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_690), .B(n_681), .C(n_686), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_672), .Y(n_720) );
AOI322xp5_ASAP7_75t_L g721 ( .A1(n_658), .A2(n_691), .A3(n_695), .B1(n_694), .B2(n_696), .C1(n_697), .C2(n_698), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_692), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_708), .A2(n_661), .B1(n_675), .B2(n_657), .C(n_674), .Y(n_723) );
AOI221xp5_ASAP7_75t_SL g724 ( .A1(n_711), .A2(n_700), .B1(n_699), .B2(n_666), .C(n_659), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_714), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_714), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_717), .Y(n_727) );
OAI211xp5_ASAP7_75t_SL g728 ( .A1(n_709), .A2(n_677), .B(n_681), .C(n_700), .Y(n_728) );
NOR2x1p5_ASAP7_75t_L g729 ( .A(n_713), .B(n_653), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g730 ( .A(n_718), .B(n_678), .C(n_671), .Y(n_730) );
NOR2xp67_ASAP7_75t_L g731 ( .A(n_713), .B(n_665), .Y(n_731) );
INVx1_ASAP7_75t_SL g732 ( .A(n_725), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_731), .A2(n_718), .B1(n_710), .B2(n_719), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_726), .Y(n_734) );
NAND4xp25_ASAP7_75t_SL g735 ( .A(n_724), .B(n_712), .C(n_721), .D(n_716), .Y(n_735) );
OAI211xp5_ASAP7_75t_SL g736 ( .A1(n_723), .A2(n_720), .B(n_687), .C(n_683), .Y(n_736) );
XNOR2x1_ASAP7_75t_L g737 ( .A(n_733), .B(n_729), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_734), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_732), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_737), .A2(n_730), .B1(n_727), .B2(n_735), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_739), .A2(n_724), .B1(n_736), .B2(n_728), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_741), .Y(n_742) );
OAI22x1_ASAP7_75t_L g743 ( .A1(n_740), .A2(n_738), .B1(n_722), .B2(n_715), .Y(n_743) );
XNOR2xp5_ASAP7_75t_L g744 ( .A(n_743), .B(n_667), .Y(n_744) );
INVxp67_ASAP7_75t_L g745 ( .A(n_744), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_745), .A2(n_742), .B1(n_685), .B2(n_701), .Y(n_746) );
endmodule