module real_aes_2811_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_498;
wire n_481;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_0), .A2(n_116), .B1(n_366), .B2(n_393), .Y(n_573) );
AOI222xp33_ASAP7_75t_L g422 ( .A1(n_1), .A2(n_109), .B1(n_139), .B2(n_341), .C1(n_423), .C2(n_424), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_2), .A2(n_212), .B1(n_366), .B2(n_393), .Y(n_663) );
OAI22x1_ASAP7_75t_L g581 ( .A1(n_3), .A2(n_582), .B1(n_583), .B2(n_613), .Y(n_581) );
INVx1_ASAP7_75t_L g613 ( .A(n_3), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_4), .A2(n_104), .B1(n_417), .B2(n_421), .Y(n_416) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_5), .A2(n_166), .B1(n_249), .B2(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g623 ( .A(n_5), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_6), .A2(n_142), .B1(n_324), .B2(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_7), .A2(n_13), .B1(n_421), .B2(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_8), .A2(n_151), .B1(n_421), .B2(n_645), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_9), .A2(n_53), .B1(n_338), .B2(n_339), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_10), .A2(n_123), .B1(n_243), .B2(n_326), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_11), .A2(n_106), .B1(n_368), .B2(n_369), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_12), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_14), .B(n_464), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_15), .A2(n_98), .B1(n_636), .B2(n_637), .Y(n_635) );
AO22x2_ASAP7_75t_L g248 ( .A1(n_16), .A2(n_51), .B1(n_249), .B2(n_250), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_16), .B(n_622), .Y(n_621) );
AO222x2_ASAP7_75t_L g384 ( .A1(n_17), .A2(n_50), .B1(n_184), .B2(n_351), .C1(n_361), .C2(n_385), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_18), .A2(n_210), .B1(n_297), .B2(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_19), .A2(n_185), .B1(n_366), .B2(n_393), .Y(n_392) );
AO222x2_ASAP7_75t_SL g657 ( .A1(n_20), .A2(n_39), .B1(n_133), .B2(n_351), .C1(n_353), .C2(n_354), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_21), .A2(n_66), .B1(n_339), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_22), .A2(n_169), .B1(n_304), .B2(n_306), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_23), .A2(n_211), .B1(n_375), .B2(n_376), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_24), .A2(n_120), .B1(n_385), .B2(n_568), .Y(n_567) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_25), .A2(n_115), .B1(n_264), .B2(n_595), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_26), .A2(n_138), .B1(n_375), .B2(n_376), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_27), .A2(n_126), .B1(n_361), .B2(n_570), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_28), .A2(n_188), .B1(n_243), .B2(n_441), .Y(n_646) );
INVx1_ASAP7_75t_L g465 ( .A(n_29), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_30), .A2(n_192), .B1(n_299), .B2(n_338), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_31), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g388 ( .A1(n_32), .A2(n_194), .B1(n_353), .B2(n_389), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_33), .A2(n_170), .B1(n_263), .B2(n_324), .Y(n_405) );
AOI222xp33_ASAP7_75t_L g340 ( .A1(n_34), .A2(n_140), .B1(n_200), .B2(n_292), .C1(n_341), .C2(n_343), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_35), .A2(n_97), .B1(n_368), .B2(n_369), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_36), .A2(n_82), .B1(n_372), .B2(n_373), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_37), .B(n_454), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_38), .A2(n_156), .B1(n_360), .B2(n_361), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_40), .A2(n_91), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_41), .A2(n_84), .B1(n_357), .B2(n_360), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_42), .A2(n_80), .B1(n_357), .B2(n_358), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_43), .A2(n_218), .B1(n_311), .B2(n_336), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_44), .A2(n_627), .B1(n_647), .B2(n_648), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_44), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_45), .A2(n_61), .B1(n_608), .B2(n_609), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_46), .A2(n_198), .B1(n_311), .B2(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_47), .A2(n_180), .B1(n_389), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_48), .A2(n_124), .B1(n_326), .B2(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_49), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_52), .A2(n_108), .B1(n_263), .B2(n_324), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_54), .A2(n_95), .B1(n_443), .B2(n_444), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_55), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_56), .A2(n_147), .B1(n_368), .B2(n_375), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_57), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g396 ( .A1(n_58), .A2(n_203), .B1(n_373), .B2(n_376), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_59), .A2(n_162), .B1(n_407), .B2(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_60), .A2(n_99), .B1(n_357), .B2(n_358), .Y(n_356) );
INVx3_ASAP7_75t_L g249 ( .A(n_62), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_63), .A2(n_130), .B1(n_369), .B2(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_64), .A2(n_137), .B1(n_297), .B2(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_65), .A2(n_167), .B1(n_263), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_67), .A2(n_103), .B1(n_373), .B2(n_398), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_68), .A2(n_86), .B1(n_326), .B2(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_69), .A2(n_101), .B1(n_297), .B2(n_299), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_70), .A2(n_160), .B1(n_332), .B2(n_408), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_71), .A2(n_121), .B1(n_373), .B2(n_398), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_72), .A2(n_161), .B1(n_336), .B2(n_449), .Y(n_448) );
OA22x2_ASAP7_75t_L g434 ( .A1(n_73), .A2(n_435), .B1(n_436), .B2(n_455), .Y(n_434) );
INVxp67_ASAP7_75t_L g455 ( .A(n_73), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_74), .Y(n_603) );
INVx1_ASAP7_75t_L g344 ( .A(n_75), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_76), .A2(n_152), .B1(n_365), .B2(n_366), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_77), .Y(n_604) );
INVx1_ASAP7_75t_SL g258 ( .A(n_78), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_78), .B(n_107), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_79), .A2(n_144), .B1(n_286), .B2(n_288), .Y(n_285) );
INVx2_ASAP7_75t_L g229 ( .A(n_81), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_83), .A2(n_195), .B1(n_267), .B2(n_518), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_85), .A2(n_93), .B1(n_336), .B2(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_87), .A2(n_219), .B1(n_277), .B2(n_493), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_88), .A2(n_163), .B1(n_332), .B2(n_333), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_89), .A2(n_165), .B1(n_286), .B2(n_443), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_90), .A2(n_110), .B1(n_277), .B2(n_281), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_92), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_94), .B(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_96), .A2(n_187), .B1(n_491), .B2(n_553), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_100), .Y(n_578) );
OA22x2_ASAP7_75t_L g458 ( .A1(n_102), .A2(n_459), .B1(n_460), .B2(n_500), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_102), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_105), .A2(n_112), .B1(n_243), .B2(n_441), .Y(n_440) );
AO22x2_ASAP7_75t_L g261 ( .A1(n_107), .A2(n_174), .B1(n_249), .B2(n_262), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_111), .A2(n_176), .B1(n_407), .B2(n_408), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_113), .A2(n_131), .B1(n_311), .B2(n_313), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_114), .A2(n_193), .B1(n_333), .B2(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_117), .A2(n_186), .B1(n_368), .B2(n_369), .Y(n_666) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_118), .A2(n_197), .B1(n_590), .B2(n_592), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g586 ( .A1(n_119), .A2(n_150), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_122), .A2(n_135), .B1(n_336), .B2(n_449), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_125), .A2(n_201), .B1(n_243), .B2(n_263), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_127), .A2(n_183), .B1(n_297), .B2(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g259 ( .A(n_128), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_129), .A2(n_190), .B1(n_353), .B2(n_354), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_132), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_134), .A2(n_178), .B1(n_267), .B2(n_271), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_136), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_141), .A2(n_177), .B1(n_547), .B2(n_548), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_143), .A2(n_172), .B1(n_286), .B2(n_329), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_145), .Y(n_484) );
INVx1_ASAP7_75t_L g534 ( .A(n_146), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_148), .A2(n_158), .B1(n_304), .B2(n_306), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_149), .B(n_471), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_153), .Y(n_498) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_154), .A2(n_223), .B(n_232), .C(n_625), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_155), .A2(n_196), .B1(n_491), .B2(n_558), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_157), .A2(n_171), .B1(n_304), .B2(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_159), .A2(n_181), .B1(n_361), .B2(n_570), .Y(n_569) );
CKINVDCx16_ASAP7_75t_R g377 ( .A(n_164), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_168), .A2(n_191), .B1(n_311), .B2(n_336), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_173), .A2(n_381), .B1(n_382), .B2(n_399), .Y(n_380) );
INVx1_ASAP7_75t_L g399 ( .A(n_173), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g492 ( .A1(n_175), .A2(n_221), .B1(n_493), .B2(n_494), .C(n_496), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_179), .A2(n_217), .B1(n_353), .B2(n_389), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_182), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g619 ( .A(n_182), .Y(n_619) );
INVx1_ASAP7_75t_L g226 ( .A(n_189), .Y(n_226) );
AND2x2_ASAP7_75t_R g650 ( .A(n_189), .B(n_619), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_199), .A2(n_214), .B1(n_412), .B2(n_477), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_202), .A2(n_215), .B1(n_304), .B2(n_343), .Y(n_508) );
OA22x2_ASAP7_75t_L g401 ( .A1(n_204), .A2(n_402), .B1(n_403), .B2(n_425), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_204), .Y(n_402) );
INVxp67_ASAP7_75t_L g231 ( .A(n_205), .Y(n_231) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_206), .A2(n_240), .B1(n_317), .B2(n_318), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_206), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_207), .B(n_292), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_208), .A2(n_220), .B1(n_311), .B2(n_313), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_209), .B(n_351), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_213), .Y(n_469) );
XNOR2x1_ASAP7_75t_L g502 ( .A(n_216), .B(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2x1_ASAP7_75t_R g224 ( .A(n_225), .B(n_227), .Y(n_224) );
OR2x2_ASAP7_75t_L g674 ( .A(n_225), .B(n_228), .Y(n_674) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_226), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_527), .B1(n_614), .B2(n_615), .C(n_616), .Y(n_232) );
INVx1_ASAP7_75t_L g615 ( .A(n_233), .Y(n_615) );
XNOR2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_430), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_378), .B1(n_428), .B2(n_429), .Y(n_234) );
INVx1_ASAP7_75t_L g428 ( .A(n_235), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B1(n_345), .B2(n_346), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OAI22xp5_ASAP7_75t_SL g237 ( .A1(n_238), .A2(n_239), .B1(n_319), .B2(n_320), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_SL g318 ( .A(n_240), .Y(n_318) );
NOR2x1_ASAP7_75t_L g240 ( .A(n_241), .B(n_290), .Y(n_240) );
NAND4xp25_ASAP7_75t_L g241 ( .A(n_242), .B(n_266), .C(n_276), .D(n_285), .Y(n_241) );
INVx2_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_SL g415 ( .A(n_244), .Y(n_415) );
INVx4_ASAP7_75t_L g488 ( .A(n_244), .Y(n_488) );
INVx3_ASAP7_75t_SL g558 ( .A(n_244), .Y(n_558) );
INVx2_ASAP7_75t_L g587 ( .A(n_244), .Y(n_587) );
INVx8_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_254), .Y(n_245) );
AND2x2_ASAP7_75t_L g269 ( .A(n_246), .B(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g279 ( .A(n_246), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g294 ( .A(n_246), .B(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g351 ( .A(n_246), .B(n_295), .Y(n_351) );
AND2x6_ASAP7_75t_L g368 ( .A(n_246), .B(n_270), .Y(n_368) );
AND2x2_ASAP7_75t_L g372 ( .A(n_246), .B(n_280), .Y(n_372) );
AND2x2_ASAP7_75t_L g375 ( .A(n_246), .B(n_254), .Y(n_375) );
AND2x2_ASAP7_75t_L g398 ( .A(n_246), .B(n_280), .Y(n_398) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_251), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g265 ( .A(n_248), .B(n_251), .Y(n_265) );
INVx1_ASAP7_75t_L g275 ( .A(n_248), .Y(n_275) );
AND2x2_ASAP7_75t_L g284 ( .A(n_248), .B(n_252), .Y(n_284) );
INVx2_ASAP7_75t_L g250 ( .A(n_249), .Y(n_250) );
INVx1_ASAP7_75t_L g253 ( .A(n_249), .Y(n_253) );
OAI22x1_ASAP7_75t_L g256 ( .A1(n_249), .A2(n_257), .B1(n_258), .B2(n_259), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_249), .Y(n_257) );
INVx1_ASAP7_75t_L g262 ( .A(n_249), .Y(n_262) );
INVxp67_ASAP7_75t_L g302 ( .A(n_251), .Y(n_302) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g274 ( .A(n_252), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g264 ( .A(n_254), .B(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g273 ( .A(n_254), .B(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g283 ( .A(n_254), .B(n_284), .Y(n_283) );
AND2x6_ASAP7_75t_L g369 ( .A(n_254), .B(n_274), .Y(n_369) );
AND2x4_ASAP7_75t_L g373 ( .A(n_254), .B(n_284), .Y(n_373) );
AND2x2_ASAP7_75t_L g376 ( .A(n_254), .B(n_265), .Y(n_376) );
AND2x4_ASAP7_75t_L g254 ( .A(n_255), .B(n_260), .Y(n_254) );
AND2x2_ASAP7_75t_L g270 ( .A(n_255), .B(n_261), .Y(n_270) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g280 ( .A(n_256), .B(n_260), .Y(n_280) );
AND2x2_ASAP7_75t_L g295 ( .A(n_256), .B(n_261), .Y(n_295) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_256), .Y(n_309) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx2_ASAP7_75t_L g289 ( .A(n_261), .Y(n_289) );
BUFx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_264), .Y(n_439) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_264), .Y(n_491) );
INVx2_ASAP7_75t_L g638 ( .A(n_264), .Y(n_638) );
AND2x4_ASAP7_75t_L g298 ( .A(n_265), .B(n_270), .Y(n_298) );
AND2x2_ASAP7_75t_L g305 ( .A(n_265), .B(n_280), .Y(n_305) );
AND2x4_ASAP7_75t_L g353 ( .A(n_265), .B(n_280), .Y(n_353) );
AND2x2_ASAP7_75t_L g360 ( .A(n_265), .B(n_270), .Y(n_360) );
AND2x2_ASAP7_75t_L g570 ( .A(n_265), .B(n_270), .Y(n_570) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g324 ( .A(n_268), .Y(n_324) );
INVx3_ASAP7_75t_L g556 ( .A(n_268), .Y(n_556) );
INVx2_ASAP7_75t_L g636 ( .A(n_268), .Y(n_636) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g495 ( .A(n_269), .Y(n_495) );
BUFx2_ASAP7_75t_L g595 ( .A(n_269), .Y(n_595) );
AND2x2_ASAP7_75t_L g287 ( .A(n_270), .B(n_274), .Y(n_287) );
AND2x2_ASAP7_75t_L g365 ( .A(n_270), .B(n_274), .Y(n_365) );
AND2x2_ASAP7_75t_SL g393 ( .A(n_270), .B(n_274), .Y(n_393) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g326 ( .A(n_272), .Y(n_326) );
INVx2_ASAP7_75t_L g441 ( .A(n_272), .Y(n_441) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_272), .Y(n_499) );
INVx2_ASAP7_75t_SL g518 ( .A(n_272), .Y(n_518) );
INVx2_ASAP7_75t_SL g588 ( .A(n_272), .Y(n_588) );
INVx8_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g312 ( .A(n_274), .B(n_280), .Y(n_312) );
AND2x4_ASAP7_75t_L g357 ( .A(n_274), .B(n_280), .Y(n_357) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_275), .Y(n_316) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g332 ( .A(n_278), .Y(n_332) );
INVx3_ASAP7_75t_L g407 ( .A(n_278), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_278), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_496) );
INVx1_ASAP7_75t_SL g597 ( .A(n_278), .Y(n_597) );
INVx6_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
BUFx3_ASAP7_75t_L g553 ( .A(n_279), .Y(n_553) );
INVx2_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_SL g446 ( .A(n_282), .Y(n_446) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx3_ASAP7_75t_L g333 ( .A(n_283), .Y(n_333) );
BUFx3_ASAP7_75t_L g408 ( .A(n_283), .Y(n_408) );
BUFx2_ASAP7_75t_SL g493 ( .A(n_283), .Y(n_493) );
AND2x4_ASAP7_75t_L g288 ( .A(n_284), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g308 ( .A(n_284), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_284), .B(n_309), .Y(n_354) );
AND2x4_ASAP7_75t_L g366 ( .A(n_284), .B(n_289), .Y(n_366) );
AND2x2_ASAP7_75t_SL g389 ( .A(n_284), .B(n_309), .Y(n_389) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g420 ( .A(n_287), .Y(n_420) );
BUFx3_ASAP7_75t_L g645 ( .A(n_287), .Y(n_645) );
INVx5_ASAP7_75t_SL g330 ( .A(n_288), .Y(n_330) );
BUFx2_ASAP7_75t_L g443 ( .A(n_288), .Y(n_443) );
NAND4xp25_ASAP7_75t_SL g290 ( .A(n_291), .B(n_296), .C(n_303), .D(n_310), .Y(n_290) );
INVx1_ASAP7_75t_L g506 ( .A(n_292), .Y(n_506) );
INVx4_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
INVx3_ASAP7_75t_L g423 ( .A(n_293), .Y(n_423) );
INVx3_ASAP7_75t_L g454 ( .A(n_293), .Y(n_454) );
INVx4_ASAP7_75t_SL g464 ( .A(n_293), .Y(n_464) );
BUFx2_ASAP7_75t_L g602 ( .A(n_293), .Y(n_602) );
INVx6_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g301 ( .A(n_295), .B(n_302), .Y(n_301) );
AND2x4_ASAP7_75t_L g314 ( .A(n_295), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g358 ( .A(n_295), .B(n_315), .Y(n_358) );
AND2x2_ASAP7_75t_L g361 ( .A(n_295), .B(n_302), .Y(n_361) );
AND2x2_ASAP7_75t_L g385 ( .A(n_295), .B(n_315), .Y(n_385) );
BUFx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_L g338 ( .A(n_298), .Y(n_338) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_298), .Y(n_477) );
BUFx2_ASAP7_75t_L g547 ( .A(n_298), .Y(n_547) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g339 ( .A(n_300), .Y(n_339) );
INVx2_ASAP7_75t_L g412 ( .A(n_300), .Y(n_412) );
INVx2_ASAP7_75t_SL g512 ( .A(n_300), .Y(n_512) );
INVx2_ASAP7_75t_L g548 ( .A(n_300), .Y(n_548) );
INVx2_ASAP7_75t_SL g641 ( .A(n_300), .Y(n_641) );
INVx6_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx5_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g342 ( .A(n_305), .Y(n_342) );
BUFx3_ASAP7_75t_L g468 ( .A(n_305), .Y(n_468) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx3_ASAP7_75t_L g471 ( .A(n_307), .Y(n_471) );
INVx2_ASAP7_75t_L g631 ( .A(n_307), .Y(n_631) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx12f_ASAP7_75t_L g343 ( .A(n_308), .Y(n_343) );
BUFx6f_ASAP7_75t_SL g608 ( .A(n_311), .Y(n_608) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx3_ASAP7_75t_L g450 ( .A(n_312), .Y(n_450) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_312), .Y(n_545) );
BUFx4f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx6f_ASAP7_75t_SL g336 ( .A(n_314), .Y(n_336) );
INVx2_ASAP7_75t_L g475 ( .A(n_314), .Y(n_475) );
INVx1_ASAP7_75t_L g610 ( .A(n_314), .Y(n_610) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
XOR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_344), .Y(n_320) );
NAND4xp75_ASAP7_75t_L g321 ( .A(n_322), .B(n_327), .C(n_334), .D(n_340), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx3_ASAP7_75t_L g421 ( .A(n_330), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g479 ( .A1(n_330), .A2(n_480), .B1(n_481), .B2(n_484), .Y(n_479) );
INVx2_ASAP7_75t_L g592 ( .A(n_330), .Y(n_592) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_333), .Y(n_598) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx3_ASAP7_75t_L g424 ( .A(n_343), .Y(n_424) );
INVx2_ASAP7_75t_L g605 ( .A(n_343), .Y(n_605) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
XOR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_377), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_348), .B(n_362), .Y(n_347) );
NOR2x1_ASAP7_75t_L g348 ( .A(n_349), .B(n_355), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx2_ASAP7_75t_SL g538 ( .A(n_351), .Y(n_538) );
INVx1_ASAP7_75t_SL g542 ( .A(n_353), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_359), .Y(n_355) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_363), .B(n_370), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_374), .Y(n_370) );
INVx1_ASAP7_75t_L g429 ( .A(n_378), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_400), .B1(n_426), .B2(n_427), .Y(n_378) );
INVx1_ASAP7_75t_L g426 ( .A(n_379), .Y(n_426) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_383), .B(n_390), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx2_ASAP7_75t_L g427 ( .A(n_400), .Y(n_427) );
BUFx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g425 ( .A(n_403), .Y(n_425) );
NAND4xp75_ASAP7_75t_L g403 ( .A(n_404), .B(n_409), .C(n_413), .D(n_422), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_419), .Y(n_444) );
INVx1_ASAP7_75t_L g483 ( .A(n_419), .Y(n_483) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g591 ( .A(n_420), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B1(n_456), .B2(n_525), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_447), .Y(n_436) );
NAND4xp25_ASAP7_75t_SL g437 ( .A(n_438), .B(n_440), .C(n_442), .D(n_445), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .C(n_452), .D(n_453), .Y(n_447) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx4_ASAP7_75t_L g568 ( .A(n_450), .Y(n_568) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g526 ( .A(n_457), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_501), .B1(n_523), .B2(n_524), .Y(n_457) );
INVx2_ASAP7_75t_L g523 ( .A(n_458), .Y(n_523) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND3x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_478), .C(n_492), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_472), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B1(n_466), .B2(n_469), .C(n_470), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
OAI222xp33_ASAP7_75t_L g600 ( .A1(n_466), .A2(n_601), .B1(n_602), .B2(n_603), .C1(n_604), .C2(n_605), .Y(n_600) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_476), .Y(n_472) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g612 ( .A(n_477), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_485), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g516 ( .A(n_483), .Y(n_516) );
OAI22xp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B1(n_489), .B2(n_490), .Y(n_485) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_488), .Y(n_522) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g524 ( .A(n_501), .Y(n_524) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_513), .Y(n_503) );
NOR2xp67_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
OAI21xp5_ASAP7_75t_SL g505 ( .A1(n_506), .A2(n_507), .B(n_508), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
NOR2x1_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g614 ( .A(n_527), .Y(n_614) );
AOI22xp5_ASAP7_75t_SL g527 ( .A1(n_528), .A2(n_529), .B1(n_579), .B2(n_580), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B1(n_559), .B2(n_560), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
XNOR2x1_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
NAND2x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_549), .Y(n_535) );
NOR2xp67_ASAP7_75t_L g536 ( .A(n_537), .B(n_543), .Y(n_536) );
OAI21xp5_ASAP7_75t_SL g537 ( .A1(n_538), .A2(n_539), .B(n_540), .Y(n_537) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
XOR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_578), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_562), .B(n_571), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_584), .B(n_599), .Y(n_583) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_593), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_600), .B(n_606), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_611), .Y(n_606) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_618), .B(n_621), .Y(n_671) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
OAI222xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_649), .B1(n_651), .B2(n_668), .C1(n_669), .C2(n_672), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_627), .Y(n_648) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR4xp25_ASAP7_75t_L g628 ( .A(n_629), .B(n_633), .C(n_639), .D(n_643), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
XOR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_668), .Y(n_654) );
NAND2x1_ASAP7_75t_L g655 ( .A(n_656), .B(n_661), .Y(n_655) );
NOR2x1_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_670), .Y(n_669) );
CKINVDCx6p67_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_673), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_674), .Y(n_673) );
endmodule