module fake_jpeg_2294_n_607 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_607);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_607;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_7),
.B(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_58),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_60),
.B(n_97),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g145 ( 
.A(n_61),
.Y(n_145)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_64),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_74),
.Y(n_168)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_75),
.Y(n_194)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

CKINVDCx9p33_ASAP7_75t_R g78 ( 
.A(n_18),
.Y(n_78)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_9),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_29),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_85),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_86),
.B(n_96),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_90),
.Y(n_192)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_91),
.Y(n_185)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

BUFx16f_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_95),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_33),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_8),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_102),
.Y(n_182)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_10),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_107),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_55),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_106),
.B(n_110),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_22),
.B(n_29),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_39),
.B(n_10),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_23),
.Y(n_144)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_119),
.B(n_138),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_74),
.A2(n_35),
.B1(n_26),
.B2(n_47),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g238 ( 
.A1(n_128),
.A2(n_188),
.B1(n_126),
.B2(n_179),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_55),
.B1(n_53),
.B2(n_49),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_135),
.A2(n_158),
.B1(n_170),
.B2(n_23),
.Y(n_207)
);

HAxp5_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_57),
.CON(n_136),
.SN(n_136)
);

NOR3xp33_ASAP7_75t_L g232 ( 
.A(n_136),
.B(n_144),
.C(n_38),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_63),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_73),
.A2(n_118),
.B1(n_87),
.B2(n_79),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_141),
.A2(n_92),
.B1(n_72),
.B2(n_34),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_142),
.B(n_30),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_101),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_148),
.B(n_160),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_94),
.A2(n_53),
.B1(n_44),
.B2(n_49),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_91),
.B(n_22),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_93),
.B(n_24),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_172),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_112),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_116),
.B(n_52),
.Y(n_172)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_71),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_90),
.Y(n_202)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g222 ( 
.A(n_186),
.Y(n_222)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_89),
.Y(n_189)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_59),
.Y(n_193)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_196),
.A2(n_225),
.B1(n_220),
.B2(n_184),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_45),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_198),
.B(n_240),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_199),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_201),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_202),
.Y(n_316)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_204),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_139),
.A2(n_35),
.B1(n_43),
.B2(n_45),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_206),
.B(n_224),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_207),
.A2(n_124),
.B1(n_157),
.B2(n_166),
.Y(n_278)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_209),
.Y(n_293)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_210),
.Y(n_295)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_211),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_134),
.B(n_24),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_212),
.B(n_218),
.Y(n_300)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_214),
.Y(n_299)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_215),
.Y(n_291)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_216),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_136),
.A2(n_117),
.B(n_32),
.C(n_82),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g285 ( 
.A1(n_217),
.A2(n_125),
.B1(n_192),
.B2(n_132),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_134),
.B(n_30),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_139),
.A2(n_35),
.B1(n_51),
.B2(n_48),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_219),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_133),
.B(n_103),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_220),
.Y(n_311)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_223),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_143),
.B(n_42),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_141),
.A2(n_34),
.B1(n_42),
.B2(n_52),
.Y(n_225)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_226),
.Y(n_323)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_227),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_143),
.B(n_66),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_228),
.B(n_229),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_123),
.B(n_51),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_160),
.A2(n_38),
.B1(n_43),
.B2(n_48),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_231),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_258),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_159),
.B(n_177),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_163),
.C(n_173),
.Y(n_268)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_234),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_131),
.B(n_82),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_235),
.B(n_236),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_164),
.B(n_26),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_152),
.B(n_67),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_237),
.B(n_239),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_238),
.A2(n_249),
.B1(n_251),
.B2(n_263),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_67),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_156),
.B(n_26),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_241),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_153),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_247),
.Y(n_297)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_162),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_244),
.Y(n_320)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_122),
.Y(n_246)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_127),
.B(n_61),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_174),
.A2(n_61),
.B1(n_47),
.B2(n_49),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_147),
.B(n_47),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_191),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_140),
.A2(n_53),
.B1(n_44),
.B2(n_32),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_137),
.B(n_11),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_254),
.Y(n_303)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_150),
.Y(n_253)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_253),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_140),
.B(n_11),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_151),
.Y(n_255)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_255),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_149),
.Y(n_256)
);

NAND2xp33_ASAP7_75t_SL g286 ( 
.A(n_256),
.B(n_260),
.Y(n_286)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_130),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_257),
.Y(n_270)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_165),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_167),
.B(n_121),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_262),
.Y(n_312)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_146),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_128),
.A2(n_25),
.B(n_32),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_261),
.B(n_25),
.Y(n_315)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_167),
.A2(n_25),
.B1(n_11),
.B2(n_12),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_185),
.A2(n_25),
.B1(n_7),
.B2(n_12),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_264),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_324)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_176),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_265),
.B(n_226),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_266),
.A2(n_222),
.B1(n_211),
.B2(n_209),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_213),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_275),
.B(n_294),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_196),
.A2(n_184),
.B1(n_176),
.B2(n_120),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_276),
.A2(n_278),
.B1(n_287),
.B2(n_313),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_197),
.C(n_198),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_277),
.B(n_282),
.C(n_306),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_171),
.C(n_190),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_120),
.B1(n_166),
.B2(n_157),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_283),
.A2(n_265),
.B1(n_223),
.B2(n_203),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_285),
.B(n_315),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_217),
.A2(n_129),
.B1(n_124),
.B2(n_130),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_145),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_208),
.B(n_145),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_298),
.B(n_307),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_221),
.B(n_149),
.C(n_155),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_200),
.B(n_0),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_261),
.A2(n_25),
.B1(n_16),
.B2(n_15),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_200),
.B(n_15),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_318),
.B(n_216),
.C(n_215),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_321),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_325),
.B(n_348),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_234),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_327),
.Y(n_392)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_280),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_329),
.Y(n_388)
);

INVx13_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_330),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_227),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_331),
.B(n_332),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_293),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_300),
.B(n_213),
.Y(n_333)
);

NAND3xp33_ASAP7_75t_L g412 ( 
.A(n_333),
.B(n_350),
.C(n_262),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_201),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_334),
.B(n_339),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_335),
.A2(n_349),
.B1(n_361),
.B2(n_362),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_195),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_338),
.B(n_369),
.C(n_306),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_293),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_322),
.Y(n_343)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_343),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_309),
.B(n_195),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_356),
.Y(n_383)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_305),
.Y(n_346)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_347),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_278),
.A2(n_238),
.B1(n_241),
.B2(n_230),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_320),
.Y(n_350)
);

INVx13_ASAP7_75t_L g351 ( 
.A(n_273),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_351),
.A2(n_357),
.B1(n_291),
.B2(n_319),
.Y(n_380)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_322),
.Y(n_352)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_352),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_353),
.A2(n_291),
.B1(n_319),
.B2(n_302),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_294),
.B(n_246),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_355),
.B(n_358),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_275),
.B(n_258),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_317),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_303),
.B(n_281),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_296),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_359),
.B(n_299),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_284),
.B(n_297),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_360),
.B(n_364),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_311),
.A2(n_238),
.B1(n_199),
.B2(n_210),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_290),
.A2(n_238),
.B1(n_204),
.B2(n_260),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_312),
.B(n_222),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_285),
.B(n_214),
.Y(n_365)
);

AND2x2_ASAP7_75t_SL g385 ( 
.A(n_365),
.B(n_371),
.Y(n_385)
);

AND2x6_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_256),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_366),
.B(n_368),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_367),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_282),
.B(n_244),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_268),
.B(n_243),
.C(n_245),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_307),
.B(n_318),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_301),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_285),
.B(n_272),
.Y(n_371)
);

OAI32xp33_ASAP7_75t_L g373 ( 
.A1(n_354),
.A2(n_290),
.A3(n_272),
.B1(n_289),
.B2(n_267),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_373),
.B(n_404),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_374),
.B(n_369),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_354),
.A2(n_272),
.B(n_289),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_376),
.A2(n_377),
.B(n_378),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_354),
.A2(n_310),
.B(n_267),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_371),
.A2(n_285),
.B(n_270),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_371),
.A2(n_270),
.B(n_296),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_379),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_380),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_384),
.A2(n_339),
.B1(n_332),
.B2(n_335),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_363),
.A2(n_283),
.B1(n_276),
.B2(n_277),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_386),
.A2(n_401),
.B1(n_402),
.B2(n_411),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_344),
.A2(n_365),
.B(n_366),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_390),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_279),
.Y(n_390)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_361),
.A2(n_308),
.B(n_301),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_398),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_340),
.A2(n_274),
.B(n_292),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_363),
.A2(n_323),
.B1(n_317),
.B2(n_288),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_349),
.A2(n_337),
.B1(n_362),
.B2(n_368),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_346),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_405),
.B(n_327),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_340),
.A2(n_292),
.B(n_274),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_350),
.Y(n_434)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_410),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_337),
.A2(n_323),
.B1(n_269),
.B2(n_302),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_328),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_410),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_422),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_325),
.C(n_336),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_423),
.C(n_433),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_416),
.A2(n_420),
.B1(n_440),
.B2(n_443),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_407),
.B(n_342),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_417),
.B(n_419),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_336),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_449),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_328),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_410),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_392),
.Y(n_424)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_424),
.Y(n_465)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_392),
.Y(n_426)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_400),
.Y(n_428)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_428),
.Y(n_480)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_400),
.Y(n_429)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_342),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_442),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_407),
.B(n_345),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_435),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_374),
.B(n_338),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_434),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_372),
.B(n_391),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_372),
.B(n_320),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_437),
.B(n_441),
.Y(n_482)
);

AO21x2_ASAP7_75t_L g439 ( 
.A1(n_378),
.A2(n_356),
.B(n_359),
.Y(n_439)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_439),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_402),
.A2(n_370),
.B1(n_348),
.B2(n_352),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_388),
.B(n_343),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_403),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_391),
.B(n_341),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_446),
.Y(n_454)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_403),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_393),
.B(n_357),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_448),
.Y(n_456)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_409),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_299),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_447),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_450),
.B(n_468),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_421),
.A2(n_399),
.B1(n_395),
.B2(n_387),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_453),
.A2(n_439),
.B1(n_386),
.B2(n_396),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_383),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_455),
.B(n_458),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_383),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_393),
.Y(n_462)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_462),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_445),
.Y(n_464)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_464),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_415),
.B(n_394),
.Y(n_466)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_466),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_423),
.B(n_376),
.C(n_379),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_471),
.C(n_477),
.Y(n_488)
);

A2O1A1O1Ixp25_ASAP7_75t_L g468 ( 
.A1(n_414),
.A2(n_436),
.B(n_431),
.C(n_440),
.D(n_425),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_424),
.B(n_394),
.Y(n_470)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_470),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_385),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_434),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_473),
.B(n_476),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_424),
.B(n_427),
.Y(n_474)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_474),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_421),
.A2(n_395),
.B1(n_401),
.B2(n_412),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_475),
.A2(n_438),
.B1(n_439),
.B2(n_396),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_427),
.B(n_390),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_431),
.B(n_385),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_425),
.B(n_438),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_398),
.C(n_377),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_463),
.B(n_458),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_486),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_425),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_487),
.A2(n_497),
.B1(n_501),
.B2(n_504),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_466),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_489),
.B(n_495),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_473),
.A2(n_427),
.B1(n_439),
.B2(n_385),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_490),
.A2(n_491),
.B1(n_464),
.B2(n_454),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_451),
.A2(n_439),
.B1(n_385),
.B2(n_430),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_460),
.B(n_409),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_455),
.B(n_373),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_499),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_469),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_498),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_461),
.B(n_482),
.Y(n_500)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_500),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_461),
.A2(n_396),
.B1(n_398),
.B2(n_448),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_457),
.B(n_467),
.C(n_471),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_462),
.C(n_456),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_469),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_457),
.B(n_381),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_505),
.B(n_506),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_477),
.B(n_411),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_479),
.A2(n_408),
.B(n_444),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_507),
.A2(n_510),
.B1(n_375),
.B2(n_397),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_472),
.A2(n_390),
.B1(n_381),
.B2(n_429),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_497),
.A2(n_451),
.B1(n_450),
.B2(n_478),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_512),
.A2(n_516),
.B1(n_397),
.B2(n_347),
.Y(n_551)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_502),
.Y(n_514)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_514),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_494),
.A2(n_478),
.B1(n_452),
.B2(n_474),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_492),
.A2(n_453),
.B1(n_476),
.B2(n_468),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_517),
.A2(n_520),
.B1(n_522),
.B2(n_533),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_518),
.A2(n_485),
.B1(n_510),
.B2(n_483),
.Y(n_542)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_509),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_519),
.B(n_524),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_494),
.A2(n_454),
.B1(n_456),
.B2(n_470),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_521),
.B(n_506),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_491),
.A2(n_465),
.B1(n_481),
.B2(n_480),
.Y(n_522)
);

FAx1_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_465),
.CI(n_480),
.CON(n_523),
.SN(n_523)
);

A2O1A1O1Ixp25_ASAP7_75t_L g541 ( 
.A1(n_523),
.A2(n_508),
.B(n_499),
.C(n_490),
.D(n_485),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_404),
.C(n_481),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_493),
.B(n_459),
.C(n_446),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_525),
.B(n_526),
.Y(n_536)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_509),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_493),
.B(n_459),
.C(n_442),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_529),
.B(n_530),
.C(n_505),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_503),
.B(n_428),
.C(n_426),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_531),
.B(n_507),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_508),
.A2(n_397),
.B1(n_389),
.B2(n_375),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_535),
.B(n_546),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_538),
.B(n_539),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_521),
.B(n_486),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_540),
.B(n_545),
.Y(n_560)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_541),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_542),
.A2(n_543),
.B1(n_553),
.B2(n_518),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_511),
.A2(n_483),
.B1(n_488),
.B2(n_496),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_524),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_534),
.B(n_513),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_513),
.B(n_488),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_549),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_525),
.B(n_389),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_SL g550 ( 
.A(n_527),
.B(n_410),
.C(n_375),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_550),
.B(n_351),
.Y(n_567)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_551),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_512),
.A2(n_269),
.B1(n_295),
.B2(n_279),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_552),
.A2(n_533),
.B1(n_523),
.B2(n_516),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_517),
.A2(n_532),
.B1(n_520),
.B2(n_522),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_554),
.B(n_555),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_545),
.B(n_529),
.C(n_528),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_556),
.B(n_557),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_548),
.A2(n_523),
.B1(n_515),
.B2(n_527),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_551),
.A2(n_515),
.B1(n_295),
.B2(n_271),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_561),
.B(n_568),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_535),
.B(n_271),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_L g581 ( 
.A(n_562),
.B(n_564),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_544),
.B(n_536),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_SL g566 ( 
.A(n_538),
.B(n_330),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_566),
.B(n_567),
.Y(n_574)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_537),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_560),
.B(n_540),
.C(n_549),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_572),
.B(n_576),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_559),
.B(n_539),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_575),
.B(n_582),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_556),
.B(n_547),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_560),
.B(n_552),
.C(n_541),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_577),
.B(n_578),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_558),
.B(n_569),
.Y(n_578)
);

AOI21xp33_ASAP7_75t_L g579 ( 
.A1(n_557),
.A2(n_351),
.B(n_257),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_579),
.A2(n_574),
.B(n_581),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_559),
.A2(n_13),
.B(n_14),
.Y(n_580)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_580),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_563),
.B(n_1),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_575),
.B(n_563),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_585),
.B(n_587),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_573),
.B(n_565),
.Y(n_587)
);

NOR3xp33_ASAP7_75t_L g589 ( 
.A(n_570),
.B(n_566),
.C(n_567),
.Y(n_589)
);

AOI322xp5_ASAP7_75t_L g595 ( 
.A1(n_589),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_574),
.C1(n_582),
.C2(n_586),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_590),
.B(n_577),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_572),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_571),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_592),
.B(n_593),
.Y(n_599)
);

A2O1A1Ixp33_ASAP7_75t_SL g600 ( 
.A1(n_595),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_584),
.B(n_583),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_596),
.A2(n_597),
.B(n_589),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_588),
.Y(n_597)
);

AO21x1_ASAP7_75t_L g601 ( 
.A1(n_598),
.A2(n_599),
.B(n_594),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_600),
.B(n_593),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_601),
.B(n_602),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_603),
.A2(n_4),
.B(n_5),
.Y(n_604)
);

BUFx24_ASAP7_75t_SL g605 ( 
.A(n_604),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_605),
.B(n_4),
.Y(n_606)
);

A2O1A1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_606),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_607)
);


endmodule