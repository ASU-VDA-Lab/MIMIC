module fake_jpeg_6756_n_276 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_0),
.C(n_1),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_24),
.C(n_35),
.Y(n_59)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_43),
.Y(n_60)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_33),
.B1(n_24),
.B2(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_47),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_0),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_16),
.B(n_9),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_18),
.Y(n_96)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_58),
.B(n_67),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_59),
.B(n_73),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_62),
.B(n_74),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_63),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_33),
.B1(n_26),
.B2(n_19),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_64),
.A2(n_78),
.B1(n_82),
.B2(n_36),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_33),
.B1(n_34),
.B2(n_17),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_68),
.A2(n_79),
.B1(n_98),
.B2(n_36),
.Y(n_108)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_39),
.B(n_17),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_29),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_77),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_16),
.B1(n_21),
.B2(n_32),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_34),
.B1(n_27),
.B2(n_32),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_43),
.B(n_22),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_89),
.B(n_99),
.C(n_84),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_41),
.A2(n_26),
.B1(n_27),
.B2(n_21),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_84),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_30),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_40),
.B(n_31),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_36),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_31),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_95),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_29),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_57),
.B(n_11),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_36),
.B1(n_23),
.B2(n_18),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_102),
.A2(n_93),
.B1(n_90),
.B2(n_63),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_105),
.B(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_124),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_23),
.B1(n_36),
.B2(n_0),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_107),
.A2(n_85),
.B1(n_9),
.B2(n_11),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_112),
.B(n_101),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_36),
.B1(n_10),
.B2(n_3),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_10),
.B1(n_15),
.B2(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_0),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_79),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_23),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_130),
.B(n_60),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_59),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_127),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_11),
.B(n_4),
.C(n_6),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_2),
.Y(n_127)
);

NAND2x1_ASAP7_75t_L g130 ( 
.A(n_58),
.B(n_6),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_15),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_7),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_61),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_138),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_128),
.B(n_132),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_137),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_69),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_69),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_162),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_97),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_97),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_70),
.Y(n_146)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_102),
.A2(n_58),
.B1(n_76),
.B2(n_86),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_147),
.A2(n_156),
.B1(n_160),
.B2(n_102),
.Y(n_194)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_152),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_85),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_154),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g152 ( 
.A(n_114),
.B(n_77),
.C(n_98),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_86),
.B1(n_76),
.B2(n_83),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_107),
.Y(n_171)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_75),
.C(n_72),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_159),
.C(n_130),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_113),
.B(n_7),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_163),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_72),
.C(n_77),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_101),
.Y(n_161)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_63),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_12),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_118),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_167),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_133),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_169),
.A2(n_176),
.B(n_103),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_174),
.Y(n_206)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_130),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_177),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_125),
.B(n_102),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_136),
.B(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_143),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_151),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_133),
.Y(n_182)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_186),
.B(n_189),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_137),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_155),
.C(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_192),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_156),
.B1(n_142),
.B2(n_119),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_R g195 ( 
.A1(n_147),
.A2(n_105),
.B1(n_118),
.B2(n_106),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_152),
.C(n_147),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_191),
.C(n_167),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_139),
.B1(n_143),
.B2(n_163),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_205),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_202),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_151),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_207),
.B(n_213),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_187),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_204),
.B(n_210),
.Y(n_222)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_157),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_135),
.B(n_141),
.C(n_149),
.D(n_109),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_160),
.B1(n_153),
.B2(n_142),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_212),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_174),
.A2(n_129),
.B1(n_140),
.B2(n_103),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_129),
.B1(n_158),
.B2(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_179),
.B(n_176),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_126),
.B1(n_148),
.B2(n_117),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_170),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_221),
.C(n_227),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_169),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_206),
.C(n_183),
.Y(n_227)
);

OAI321xp33_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_207),
.A3(n_202),
.B1(n_180),
.B2(n_215),
.C(n_198),
.Y(n_228)
);

OAI321xp33_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_210),
.A3(n_213),
.B1(n_208),
.B2(n_175),
.C(n_214),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_170),
.B(n_208),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_182),
.C(n_192),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_231),
.C(n_237),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_168),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_168),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_233),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_177),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_197),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_181),
.C(n_188),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_235),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_249),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_221),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_220),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_251),
.B(n_222),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_246),
.B(n_185),
.Y(n_262)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_226),
.A2(n_229),
.B1(n_224),
.B2(n_225),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_212),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_224),
.C(n_231),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_253),
.A2(n_260),
.B(n_258),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_234),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_218),
.C(n_211),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_201),
.B1(n_193),
.B2(n_185),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_259),
.A2(n_172),
.B1(n_184),
.B2(n_173),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_247),
.B(n_166),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_248),
.B(n_172),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_244),
.B(n_250),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_263),
.A2(n_266),
.B(n_254),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_173),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_265),
.B(n_184),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_262),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_265),
.A2(n_256),
.B(n_255),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_272),
.B(n_117),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_13),
.Y(n_276)
);


endmodule