module real_jpeg_5846_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_313;
wire n_42;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_0),
.A2(n_273),
.B1(n_276),
.B2(n_277),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_0),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_0),
.A2(n_276),
.B1(n_371),
.B2(n_373),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_0),
.A2(n_72),
.B1(n_276),
.B2(n_405),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_L g466 ( 
.A1(n_0),
.A2(n_276),
.B1(n_341),
.B2(n_467),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_85),
.B1(n_89),
.B2(n_92),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_1),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_1),
.A2(n_92),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_1),
.A2(n_92),
.B1(n_182),
.B2(n_383),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_1),
.A2(n_92),
.B1(n_419),
.B2(n_421),
.Y(n_418)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_2),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_2),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_2),
.Y(n_234)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_2),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_2),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_2),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_2),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_95),
.B1(n_98),
.B2(n_102),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_3),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_3),
.A2(n_102),
.B1(n_131),
.B2(n_134),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_3),
.A2(n_102),
.B1(n_142),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_3),
.A2(n_102),
.B1(n_312),
.B2(n_351),
.Y(n_389)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_4),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_4),
.Y(n_149)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_4),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_4),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_4),
.Y(n_440)
);

INVx6_ASAP7_75t_L g469 ( 
.A(n_4),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_5),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_5),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_127),
.C(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_5),
.B(n_73),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_5),
.B(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_5),
.B(n_129),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_5),
.B(n_97),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_6),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_6),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_6),
.A2(n_183),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_6),
.A2(n_183),
.B1(n_302),
.B2(n_367),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_6),
.A2(n_183),
.B1(n_341),
.B2(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_7),
.Y(n_333)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_8),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_9),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_9),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_9),
.A2(n_170),
.B1(n_200),
.B2(n_203),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_9),
.A2(n_170),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_9),
.A2(n_149),
.B1(n_170),
.B2(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_12),
.Y(n_122)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_12),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_12),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_13),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_13),
.A2(n_57),
.B1(n_311),
.B2(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_13),
.A2(n_57),
.B1(n_396),
.B2(n_398),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_13),
.A2(n_57),
.B1(n_452),
.B2(n_454),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_14),
.Y(n_547)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_16),
.A2(n_32),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_16),
.A2(n_50),
.B1(n_311),
.B2(n_313),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_16),
.A2(n_50),
.B1(n_208),
.B2(n_392),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_16),
.A2(n_50),
.B1(n_267),
.B2(n_410),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_17),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_17),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_17),
.A2(n_209),
.B1(n_227),
.B2(n_230),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_17),
.A2(n_209),
.B1(n_299),
.B2(n_302),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_17),
.A2(n_48),
.B1(n_209),
.B2(n_439),
.Y(n_438)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_543),
.B(n_545),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_152),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_150),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_147),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_23),
.B(n_147),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_138),
.C(n_144),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_24),
.A2(n_25),
.B1(n_539),
.B2(n_540),
.Y(n_538)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_58),
.C(n_103),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_26),
.B(n_531),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_47),
.B1(n_51),
.B2(n_53),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_27),
.A2(n_51),
.B1(n_53),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_27),
.A2(n_51),
.B1(n_139),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_27),
.A2(n_360),
.B(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_27),
.A2(n_51),
.B1(n_413),
.B2(n_438),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_27),
.A2(n_47),
.B1(n_51),
.B2(n_516),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_28),
.A2(n_358),
.B(n_359),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_28),
.B(n_361),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_34),
.Y(n_140)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_39),
.B1(n_42),
.B2(n_45),
.Y(n_38)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_36),
.Y(n_335)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_44),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_44),
.Y(n_268)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_SL g358 ( 
.A1(n_48),
.A2(n_165),
.B(n_338),
.Y(n_358)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_51),
.B(n_165),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_51),
.A2(n_438),
.B(n_470),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_52),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_52),
.B(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_58),
.A2(n_103),
.B1(n_104),
.B2(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_58),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_84),
.B1(n_93),
.B2(n_94),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_59),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_59),
.A2(n_93),
.B1(n_298),
.B2(n_366),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_59),
.A2(n_93),
.B1(n_404),
.B2(n_409),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_59),
.A2(n_84),
.B1(n_93),
.B2(n_520),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_73),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_65),
.B1(n_69),
.B2(n_71),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_68),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_68),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_68),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_69),
.B(n_133),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_73),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_73),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

AOI22x1_ASAP7_75t_L g441 ( 
.A1(n_73),
.A2(n_145),
.B1(n_306),
.B2(n_442),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_73),
.A2(n_145),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_81),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g210 ( 
.A(n_75),
.Y(n_210)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_77),
.Y(n_397)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_79),
.Y(n_372)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_83),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_88),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_88),
.Y(n_411)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_93),
.B(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_93),
.A2(n_298),
.B(n_305),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_101),
.Y(n_262)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_101),
.Y(n_327)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_101),
.Y(n_337)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_101),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_103),
.A2(n_104),
.B1(n_518),
.B2(n_519),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_103),
.B(n_515),
.C(n_518),
.Y(n_526)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_128),
.B(n_130),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_105),
.A2(n_162),
.B(n_166),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_105),
.A2(n_128),
.B1(n_207),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_105),
.A2(n_166),
.B(n_255),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_105),
.A2(n_128),
.B1(n_370),
.B2(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_106),
.B(n_167),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_106),
.A2(n_129),
.B1(n_391),
.B2(n_395),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_106),
.A2(n_129),
.B1(n_395),
.B2(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_106),
.A2(n_129),
.B1(n_418),
.B2(n_457),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_114),
.B2(n_116),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_110),
.Y(n_394)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_SL g208 ( 
.A(n_116),
.Y(n_208)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_117),
.A2(n_207),
.B(n_211),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_123),
.B2(n_126),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_124),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_128),
.A2(n_211),
.B(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_130),
.Y(n_457)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_133),
.Y(n_420)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_136),
.Y(n_283)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_137),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_138),
.B(n_144),
.Y(n_540)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_145),
.A2(n_261),
.B(n_265),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_145),
.B(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_145),
.A2(n_265),
.B(n_483),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_149),
.Y(n_363)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_149),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_537),
.B(n_542),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_509),
.B(n_534),
.Y(n_153)
);

OAI311xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_376),
.A3(n_485),
.B1(n_503),
.C1(n_508),
.Y(n_154)
);

AOI21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_318),
.B(n_375),
.Y(n_155)
);

AO21x1_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_289),
.B(n_317),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_249),
.B(n_288),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_214),
.B(n_248),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_179),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_160),
.B(n_179),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_172),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_161),
.A2(n_172),
.B1(n_173),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_161),
.Y(n_246)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_165),
.A2(n_189),
.B(n_196),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_SL g261 ( 
.A1(n_165),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_165),
.B(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_169),
.Y(n_257)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_171),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx5_ASAP7_75t_L g422 ( 
.A(n_175),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_177),
.Y(n_313)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_204),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_180),
.B(n_205),
.C(n_213),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_189),
.B(n_196),
.Y(n_180)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_186),
.Y(n_277)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_188),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_188),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_189),
.A2(n_344),
.B1(n_345),
.B2(n_348),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_189),
.A2(n_382),
.B1(n_386),
.B2(n_389),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_189),
.A2(n_389),
.B(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_199),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_190),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_190),
.A2(n_272),
.B1(n_310),
.B2(n_314),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_190),
.A2(n_349),
.B1(n_433),
.B2(n_434),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_202),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_212),
.B2(n_213),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_208),
.Y(n_258)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_238),
.B(n_247),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_224),
.B(n_237),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_223),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx8_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_236),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_236),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_232),
.B(n_235),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_234),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_271),
.B(n_278),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_245),
.Y(n_247)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_244),
.Y(n_347)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_244),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_251),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_269),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_259),
.B2(n_260),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_259),
.C(n_269),
.Y(n_290)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI32xp33_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_280),
.A3(n_281),
.B1(n_284),
.B2(n_287),
.Y(n_279)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_268),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_279),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_279),
.Y(n_295)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_275),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_290),
.B(n_291),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_296),
.B2(n_316),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_295),
.C(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_307),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_297),
.B(n_308),
.C(n_309),
.Y(n_352)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx12f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_301),
.Y(n_453)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_310),
.Y(n_344)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_319),
.B(n_320),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_355),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_321)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_324),
.B1(n_342),
.B2(n_343),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_324),
.B(n_342),
.Y(n_481)
);

OAI32xp33_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_328),
.A3(n_331),
.B1(n_334),
.B2(n_338),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_352),
.B(n_353),
.C(n_355),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_364),
.B2(n_374),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_356),
.B(n_365),
.C(n_369),
.Y(n_494)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_364),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_369),
.Y(n_364)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_366),
.Y(n_483)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp33_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_471),
.Y(n_376)
);

A2O1A1Ixp33_ASAP7_75t_SL g503 ( 
.A1(n_377),
.A2(n_471),
.B(n_504),
.C(n_507),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_443),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_378),
.B(n_443),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_415),
.C(n_428),
.Y(n_378)
);

FAx1_ASAP7_75t_SL g484 ( 
.A(n_379),
.B(n_415),
.CI(n_428),
.CON(n_484),
.SN(n_484)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_402),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_380),
.B(n_403),
.C(n_412),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_390),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_381),
.B(n_390),
.Y(n_477)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_391),
.Y(n_431)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx8_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_412),
.Y(n_402)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_409),
.Y(n_450)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_416),
.A2(n_417),
.B1(n_423),
.B2(n_427),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_417),
.B(n_423),
.Y(n_461)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_423),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_423),
.A2(n_427),
.B1(n_463),
.B2(n_464),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_423),
.A2(n_461),
.B(n_464),
.Y(n_512)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_436),
.C(n_441),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_429),
.B(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_430),
.B(n_432),
.Y(n_493)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_436),
.A2(n_437),
.B1(n_441),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_441),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_444),
.B(n_447),
.C(n_459),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_447),
.B1(n_459),
.B2(n_460),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_455),
.B(n_458),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_456),
.Y(n_458)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_451),
.Y(n_520)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

FAx1_ASAP7_75t_SL g511 ( 
.A(n_458),
.B(n_512),
.CI(n_513),
.CON(n_511),
.SN(n_511)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_458),
.B(n_512),
.C(n_513),
.Y(n_533)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_470),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_466),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_468),
.Y(n_467)
);

INVx8_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_484),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_484),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_477),
.C(n_478),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_473),
.A2(n_474),
.B1(n_477),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_496),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.C(n_482),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_479),
.A2(n_480),
.B1(n_482),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g548 ( 
.A(n_484),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_486),
.B(n_498),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_487),
.A2(n_505),
.B(n_506),
.Y(n_504)
);

NOR2x1_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_495),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_495),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_492),
.C(n_494),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_501),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_492),
.A2(n_493),
.B1(n_494),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_494),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_500),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_523),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_511),
.B(n_522),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_511),
.B(n_522),
.Y(n_535)
);

BUFx24_ASAP7_75t_SL g550 ( 
.A(n_511),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_514),
.A2(n_515),
.B1(n_517),
.B2(n_521),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_514),
.A2(n_515),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_514),
.B(n_525),
.C(n_529),
.Y(n_541)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_517),
.Y(n_521)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_523),
.A2(n_535),
.B(n_536),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_524),
.B(n_533),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_533),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_525),
.A2(n_526),
.B1(n_527),
.B2(n_528),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_541),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_541),
.Y(n_542)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx13_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx8_ASAP7_75t_L g546 ( 
.A(n_544),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_547),
.Y(n_545)
);


endmodule