module fake_jpeg_31020_n_93 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_47),
.Y(n_60)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_1),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_50),
.C(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_27),
.B(n_1),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_28),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_35),
.Y(n_61)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_2),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_36),
.B1(n_35),
.B2(n_26),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_34),
.B(n_4),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_58),
.C(n_61),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_43),
.B1(n_51),
.B2(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_61),
.B1(n_34),
.B2(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_60),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_79),
.B(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_80),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_78),
.B1(n_74),
.B2(n_72),
.Y(n_85)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_74),
.C(n_81),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_85),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_38),
.A3(n_37),
.B1(n_31),
.B2(n_10),
.C1(n_13),
.C2(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_7),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_87),
.Y(n_88)
);

OA21x2_ASAP7_75t_SL g90 ( 
.A1(n_88),
.A2(n_19),
.B(n_22),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_89),
.A2(n_24),
.B(n_3),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_91),
.Y(n_93)
);


endmodule