module fake_jpeg_7959_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_14),
.Y(n_67)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_0),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_25),
.B1(n_18),
.B2(n_22),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_59),
.B1(n_60),
.B2(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_18),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_49),
.C(n_55),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_25),
.B1(n_18),
.B2(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_51),
.B1(n_38),
.B2(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_32),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_25),
.B1(n_19),
.B2(n_26),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_54),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_0),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_20),
.C(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_21),
.B1(n_31),
.B2(n_26),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_17),
.B1(n_29),
.B2(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_30),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_17),
.B(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_13),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_28),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_41),
.C(n_40),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_15),
.Y(n_78)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_70),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_71),
.B(n_78),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_72),
.A2(n_75),
.B1(n_90),
.B2(n_93),
.Y(n_120)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_73),
.A2(n_47),
.B1(n_57),
.B2(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_74),
.B(n_86),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_77),
.Y(n_124)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_33),
.B(n_38),
.C(n_34),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_47),
.B(n_57),
.C(n_63),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_15),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_97),
.B(n_99),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_39),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_65),
.C(n_63),
.Y(n_110)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_39),
.B1(n_36),
.B2(n_41),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_41),
.B1(n_40),
.B2(n_28),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_12),
.Y(n_94)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_54),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_102),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_53),
.A2(n_34),
.B1(n_22),
.B2(n_28),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_53),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_34),
.A3(n_28),
.B1(n_22),
.B2(n_35),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_61),
.A3(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_108),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_107),
.A2(n_85),
.B1(n_79),
.B2(n_76),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_49),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_123),
.B(n_128),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_77),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_119),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_53),
.B1(n_54),
.B2(n_59),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_80),
.B1(n_102),
.B2(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_59),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_126),
.B1(n_90),
.B2(n_75),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_40),
.A3(n_41),
.B1(n_32),
.B2(n_7),
.Y(n_126)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_131),
.B(n_134),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_132),
.B(n_141),
.Y(n_184)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_98),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_100),
.B1(n_72),
.B2(n_74),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_139),
.B1(n_120),
.B2(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_92),
.B1(n_101),
.B2(n_93),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_121),
.B1(n_130),
.B2(n_126),
.Y(n_140)
);

AO22x1_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_116),
.B1(n_115),
.B2(n_112),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_103),
.B(n_86),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_142),
.B(n_143),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_103),
.B(n_86),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_87),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_85),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_113),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_158),
.C(n_159),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_154),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_157),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_115),
.A2(n_73),
.B(n_91),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_109),
.B(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_119),
.B(n_11),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_129),
.B(n_10),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_1),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_164),
.A2(n_170),
.B1(n_187),
.B2(n_5),
.Y(n_215)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_153),
.B(n_110),
.CI(n_109),
.CON(n_165),
.SN(n_165)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_165),
.B(n_168),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_120),
.B1(n_112),
.B2(n_127),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_109),
.B(n_110),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_158),
.B(n_159),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_179),
.B(n_181),
.Y(n_193)
);

NOR2x1_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_106),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_174),
.B(n_177),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_152),
.A2(n_114),
.B1(n_89),
.B2(n_111),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_182),
.B(n_6),
.Y(n_207)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_11),
.C(n_16),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_111),
.B1(n_89),
.B2(n_69),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_132),
.B1(n_131),
.B2(n_134),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

AOI32xp33_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_68),
.A3(n_8),
.B1(n_10),
.B2(n_15),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_133),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_189),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_146),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_173),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_192),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_157),
.B1(n_141),
.B2(n_148),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_209),
.B1(n_211),
.B2(n_214),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_151),
.C(n_153),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_201),
.C(n_203),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_207),
.B1(n_210),
.B2(n_176),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_145),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_199),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_154),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_168),
.A2(n_136),
.B(n_140),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_206),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_150),
.C(n_159),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_190),
.B(n_169),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_138),
.C(n_149),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_213),
.C(n_185),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_181),
.A2(n_143),
.B(n_161),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_162),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_174),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_166),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_189),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_6),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_4),
.B1(n_5),
.B2(n_12),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_176),
.B1(n_185),
.B2(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_228),
.B1(n_235),
.B2(n_208),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_213),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_227),
.Y(n_242)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_165),
.C(n_162),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_205),
.C(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_233),
.B1(n_188),
.B2(n_178),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_201),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_237),
.C(n_240),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_203),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_243),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_226),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_200),
.C(n_190),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_245),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_194),
.Y(n_245)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_247),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_170),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_228),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_257),
.B(n_260),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_216),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_256),
.B(n_259),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_231),
.B(n_230),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_249),
.A2(n_232),
.B(n_224),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_239),
.B(n_221),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_183),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_167),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_225),
.B(n_227),
.Y(n_272)
);

OAI221xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_223),
.B1(n_211),
.B2(n_207),
.C(n_244),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_270),
.B(n_198),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_198),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_269),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_240),
.C(n_243),
.Y(n_269)
);

OAI221xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_206),
.B1(n_233),
.B2(n_164),
.C(n_187),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_241),
.C(n_248),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_271),
.B(n_275),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_180),
.B(n_222),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_254),
.C(n_258),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_264),
.C(n_261),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_281),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_267),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_280),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_279),
.A2(n_265),
.B(n_180),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_210),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_222),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_175),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_282),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_290),
.B(n_285),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_286),
.A2(n_277),
.B(n_284),
.C(n_276),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_285),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_SL g294 ( 
.A1(n_292),
.A2(n_293),
.B(n_163),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_163),
.Y(n_295)
);


endmodule