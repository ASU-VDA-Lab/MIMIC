module fake_jpeg_10328_n_199 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_32),
.Y(n_56)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_31),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_24),
.B1(n_23),
.B2(n_28),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_26),
.Y(n_74)
);

CKINVDCx12_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_25),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_71),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_35),
.C(n_39),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_77),
.C(n_31),
.Y(n_98)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_23),
.B1(n_28),
.B2(n_33),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_52),
.B1(n_68),
.B2(n_56),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_34),
.B1(n_39),
.B2(n_46),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_76),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_32),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_51),
.B(n_60),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_98),
.C(n_27),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_46),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_89),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_97),
.B1(n_72),
.B2(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_64),
.B1(n_71),
.B2(n_74),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_80),
.B1(n_56),
.B2(n_44),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_93),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_75),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_15),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_58),
.B(n_52),
.C(n_40),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_27),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_104),
.Y(n_126)
);

AO21x2_ASAP7_75t_SL g102 ( 
.A1(n_99),
.A2(n_69),
.B(n_44),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_102),
.A2(n_108),
.B(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_119),
.C(n_30),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_110),
.Y(n_123)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_25),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_30),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_0),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_21),
.B(n_19),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_91),
.B1(n_84),
.B2(n_94),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_94),
.B1(n_100),
.B2(n_82),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_90),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_21),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_15),
.C(n_19),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_96),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_119),
.C(n_116),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_138),
.C(n_148),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_116),
.C(n_102),
.Y(n_138)
);

OAI321xp33_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_112),
.A3(n_109),
.B1(n_105),
.B2(n_108),
.C(n_26),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_128),
.A3(n_121),
.B1(n_126),
.B2(n_134),
.C1(n_129),
.C2(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_120),
.B(n_112),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_150),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_20),
.B(n_12),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_155),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_131),
.B1(n_136),
.B2(n_132),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_162),
.B1(n_147),
.B2(n_1),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_133),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_160),
.C(n_137),
.Y(n_165)
);

NAND4xp25_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_82),
.C(n_95),
.D(n_21),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_163),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_29),
.C(n_22),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_22),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_9),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_29),
.B1(n_20),
.B2(n_7),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_166),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_148),
.C(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_171),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_147),
.B(n_11),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_168),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_169),
.Y(n_182)
);

AO22x1_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_173),
.A2(n_162),
.B1(n_160),
.B2(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_8),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_178),
.B(n_180),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_155),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_181),
.B(n_2),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_172),
.A3(n_173),
.B1(n_165),
.B2(n_158),
.C1(n_5),
.C2(n_1),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_185),
.B(n_175),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_187),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_2),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_176),
.B(n_178),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_183),
.B1(n_188),
.B2(n_179),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_192),
.Y(n_193)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_3),
.B(n_4),
.Y(n_196)
);

OAI211xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_193),
.B(n_3),
.C(n_6),
.Y(n_198)
);

AOI21x1_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_6),
.B(n_197),
.Y(n_199)
);


endmodule