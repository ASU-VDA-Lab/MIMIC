module fake_jpeg_1062_n_225 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_225);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_1),
.Y(n_94)
);

BUFx4f_ASAP7_75t_SL g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx6p67_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_56),
.B1(n_72),
.B2(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_56),
.B1(n_72),
.B2(n_71),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_79),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_71),
.B1(n_73),
.B2(n_69),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_73),
.B1(n_67),
.B2(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_104),
.Y(n_122)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_54),
.B(n_58),
.C(n_63),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_112),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_95),
.B1(n_80),
.B2(n_87),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_62),
.B1(n_60),
.B2(n_76),
.Y(n_137)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_75),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_70),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_61),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_84),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_25),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_118),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_60),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_121),
.C(n_99),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_55),
.C(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_66),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_102),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_53),
.B(n_74),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_129),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_84),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_53),
.B1(n_84),
.B2(n_55),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_133),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_110),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_62),
.B1(n_60),
.B2(n_76),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_1),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_140),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_136),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_141),
.B(n_146),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_107),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_147),
.Y(n_167)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_99),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_156),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_76),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_169)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_159),
.Y(n_165)
);

INVx5_ASAP7_75t_SL g158 ( 
.A(n_129),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_168)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_48),
.C(n_46),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_30),
.C(n_29),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_3),
.B(n_4),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_7),
.B(n_8),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_124),
.B(n_117),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_175),
.B1(n_28),
.B2(n_27),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_172),
.B1(n_173),
.B2(n_178),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_6),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_170),
.B(n_14),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_156),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_22),
.B1(n_36),
.B2(n_31),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_151),
.B(n_148),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_182),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_192),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_160),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_153),
.B1(n_152),
.B2(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_194),
.B1(n_195),
.B2(n_174),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_142),
.B(n_39),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_191),
.Y(n_201)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_193),
.A2(n_168),
.B1(n_171),
.B2(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_16),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_166),
.C(n_162),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_202),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_205),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_203),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_181),
.C(n_167),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_189),
.A2(n_181),
.B1(n_18),
.B2(n_19),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_191),
.B(n_185),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_212),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_193),
.A3(n_192),
.B1(n_188),
.B2(n_182),
.C1(n_21),
.C2(n_17),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_210),
.B(n_17),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_193),
.B(n_26),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_209),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_216),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_196),
.B1(n_214),
.B2(n_208),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_219),
.A2(n_217),
.B(n_214),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_211),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

OAI311xp33_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_197),
.A3(n_198),
.B1(n_20),
.C1(n_18),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_19),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_20),
.Y(n_225)
);


endmodule