module real_jpeg_6724_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_1),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_1),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_1),
.A2(n_117),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_1),
.A2(n_117),
.B1(n_294),
.B2(n_296),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_1),
.A2(n_117),
.B1(n_364),
.B2(n_369),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_3),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_3),
.A2(n_127),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_3),
.A2(n_90),
.B1(n_127),
.B2(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_3),
.A2(n_127),
.B1(n_173),
.B2(n_398),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_4),
.A2(n_106),
.B1(n_110),
.B2(n_111),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_4),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_4),
.A2(n_110),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_4),
.A2(n_42),
.B1(n_110),
.B2(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_4),
.A2(n_110),
.B1(n_344),
.B2(n_380),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_5),
.B(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_5),
.B(n_168),
.C(n_267),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g270 ( 
.A1(n_5),
.A2(n_271),
.B1(n_272),
.B2(n_274),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_5),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_5),
.B(n_153),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_5),
.A2(n_24),
.B1(n_315),
.B2(n_318),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_5),
.B(n_202),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_5),
.A2(n_235),
.B(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_6),
.A2(n_224),
.B1(n_248),
.B2(n_251),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_6),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_6),
.A2(n_251),
.B1(n_278),
.B2(n_281),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_6),
.A2(n_251),
.B1(n_299),
.B2(n_316),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_6),
.A2(n_251),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_7),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_8),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_8),
.Y(n_189)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_8),
.Y(n_320)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_8),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_9),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_9),
.A2(n_46),
.B1(n_73),
.B2(n_76),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_9),
.A2(n_46),
.B1(n_155),
.B2(n_158),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_10),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_10),
.Y(n_230)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_12),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_12),
.Y(n_120)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_12),
.Y(n_226)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_12),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_13),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_13),
.A2(n_35),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_15),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_15),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_15),
.A2(n_81),
.B1(n_155),
.B2(n_156),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_15),
.A2(n_43),
.B1(n_81),
.B2(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_256),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_254),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_206),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_19),
.B(n_206),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_159),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.C(n_122),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_22),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_23),
.B(n_50),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_38),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_24),
.A2(n_163),
.B(n_165),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_24),
.B(n_41),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_24),
.A2(n_30),
.B1(n_240),
.B2(n_245),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_24),
.A2(n_185),
.B(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_24),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_24),
.A2(n_304),
.B1(n_315),
.B2(n_318),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_24),
.A2(n_38),
.B(n_165),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_27),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_29),
.Y(n_309)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_37),
.Y(n_295)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_37),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_44),
.Y(n_317)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_45),
.Y(n_244)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_48),
.B(n_324),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_71),
.B1(n_78),
.B2(n_85),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_51),
.A2(n_170),
.B(n_177),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_51),
.A2(n_394),
.B(n_395),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_51),
.A2(n_177),
.B(n_397),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_52),
.A2(n_171),
.B1(n_178),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_52),
.A2(n_178),
.B1(n_270),
.B2(n_277),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_52),
.A2(n_178),
.B1(n_277),
.B2(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_52),
.A2(n_178),
.B1(n_288),
.B2(n_363),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_64),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_53)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_54),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_55),
.Y(n_273)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_55),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_61),
.Y(n_282)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_62),
.Y(n_280)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_62),
.Y(n_341)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_63),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_64)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_66),
.Y(n_168)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_70),
.Y(n_268)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_72),
.B(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_75),
.Y(n_289)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_85),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_85),
.B(n_271),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_85),
.B(n_397),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_86),
.A2(n_87),
.B1(n_122),
.B2(n_123),
.Y(n_208)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_105),
.B1(n_114),
.B2(n_121),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_88),
.A2(n_114),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_88),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_88),
.A2(n_121),
.B1(n_414),
.B2(n_417),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_98),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_95),
.Y(n_89)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_90),
.Y(n_201)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_97),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_98),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_100),
.Y(n_223)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_101),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_101),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_105),
.Y(n_253)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_132),
.B(n_152),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_124),
.B(n_134),
.Y(n_218)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_125),
.Y(n_338)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_131),
.Y(n_346)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_131),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_132),
.A2(n_134),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_132),
.A2(n_134),
.B1(n_379),
.B2(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_133),
.B(n_154),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_133),
.A2(n_213),
.B(n_218),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_133),
.A2(n_153),
.B1(n_353),
.B2(n_358),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_143),
.Y(n_133)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_134),
.A2(n_195),
.B(n_196),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_134)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_137),
.Y(n_342)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_139),
.Y(n_349)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_140),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_149),
.B2(n_151),
.Y(n_143)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_180),
.B1(n_204),
.B2(n_205),
.Y(n_159)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_169),
.B2(n_179),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_193),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_190),
.B1(n_191),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_184),
.A2(n_241),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_197),
.B1(n_198),
.B2(n_203),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_202),
.A2(n_247),
.B1(n_252),
.B2(n_253),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_207),
.B(n_209),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_211),
.B(n_422),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.C(n_246),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_212),
.B(n_246),
.Y(n_425)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_213),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx6_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_219),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_239),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_220),
.B(n_239),
.Y(n_407)
);

OAI32xp33_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_224),
.A3(n_227),
.B1(n_231),
.B2(n_234),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g361 ( 
.A(n_223),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_226),
.Y(n_416)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_244),
.Y(n_305)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_247),
.Y(n_417)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_419),
.B(n_432),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_403),
.B(n_418),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_372),
.B(n_402),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_332),
.B(n_371),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_300),
.B(n_331),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_283),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_263),
.B(n_283),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_269),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_264),
.B(n_269),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_271),
.B(n_344),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_SL g353 ( 
.A1(n_271),
.A2(n_343),
.B(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_273),
.Y(n_370)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_292),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_291),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_291),
.C(n_292),
.Y(n_333)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_287),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_290),
.B(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_311),
.B(n_330),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_310),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_310),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_321),
.B(n_329),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_313),
.B(n_314),
.Y(n_329)
);

INVx4_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_325),
.Y(n_387)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_334),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_351),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_335),
.B(n_352),
.C(n_362),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_350),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_336),
.B(n_350),
.Y(n_392)
);

OAI32xp33_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_339),
.A3(n_342),
.B1(n_343),
.B2(n_347),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_362),
.Y(n_351)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_356),
.Y(n_359)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_373),
.B(n_374),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_390),
.B2(n_391),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_393),
.C(n_400),
.Y(n_404)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_384),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_385),
.C(n_389),
.Y(n_408)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_386),
.B1(n_388),
.B2(n_389),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_388),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_392),
.A2(n_393),
.B1(n_400),
.B2(n_401),
.Y(n_391)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_392),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_393),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_405),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_408),
.C(n_409),
.Y(n_429)
);

BUFx24_ASAP7_75t_SL g435 ( 
.A(n_409),
.Y(n_435)
);

FAx1_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_412),
.CI(n_413),
.CON(n_409),
.SN(n_409)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_412),
.C(n_413),
.Y(n_426)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_428),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_420),
.A2(n_433),
.B(n_434),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_423),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_423),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_426),
.C(n_427),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_426),
.B(n_427),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_429),
.B(n_430),
.Y(n_433)
);


endmodule