module fake_ariane_1656_n_3294 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_830, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_850, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_806, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_864, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_520, n_870, n_87, n_714, n_279, n_702, n_207, n_790, n_857, n_363, n_720, n_354, n_41, n_813, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_829, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_855, n_158, n_69, n_259, n_835, n_95, n_808, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_858, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_840, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_3, n_271, n_465, n_486, n_507, n_759, n_247, n_569, n_567, n_825, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_831, n_256, n_868, n_326, n_681, n_778, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_823, n_620, n_228, n_325, n_276, n_93, n_688, n_859, n_636, n_427, n_108, n_587, n_497, n_693, n_863, n_303, n_671, n_442, n_777, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_843, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_775, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_869, n_141, n_846, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_844, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_861, n_175, n_711, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_847, n_371, n_845, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_865, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_860, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_851, n_255, n_560, n_450, n_257, n_842, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_853, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_848, n_804, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_834, n_83, n_389, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_213, n_862, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_785, n_827, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_793, n_852, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_866, n_26, n_246, n_517, n_530, n_0, n_792, n_824, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_773, n_165, n_144, n_317, n_867, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_856, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_618, n_411, n_484, n_712, n_849, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_797, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_828, n_595, n_322, n_251, n_506, n_602, n_799, n_558, n_592, n_116, n_397, n_841, n_854, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_783, n_675, n_3294);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_850;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_864;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_870;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_790;
input n_857;
input n_363;
input n_720;
input n_354;
input n_41;
input n_813;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_829;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_855;
input n_158;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_858;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_840;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_831;
input n_256;
input n_868;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_823;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_859;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_863;
input n_303;
input n_671;
input n_442;
input n_777;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_843;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_869;
input n_141;
input n_846;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_844;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_861;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_847;
input n_371;
input n_845;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_865;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_860;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_851;
input n_255;
input n_560;
input n_450;
input n_257;
input n_842;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_853;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_848;
input n_804;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_83;
input n_389;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_862;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_785;
input n_827;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_793;
input n_852;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_866;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_792;
input n_824;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_773;
input n_165;
input n_144;
input n_317;
input n_867;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_856;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_618;
input n_411;
input n_484;
input n_712;
input n_849;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_841;
input n_854;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_783;
input n_675;

output n_3294;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_3152;
wire n_2346;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_3181;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_924;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_2006;
wire n_952;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_2976;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_3145;
wire n_2248;
wire n_3063;
wire n_3281;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_1062;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_3252;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_3144;
wire n_2359;
wire n_2201;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_1404;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_1900;
wire n_1074;
wire n_3230;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_2650;
wire n_1254;
wire n_929;
wire n_3207;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_3073;
wire n_2060;
wire n_1295;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3013;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1840;
wire n_1230;
wire n_2739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_3271;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_1216;
wire n_3126;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3119;
wire n_1108;
wire n_1590;
wire n_1351;
wire n_3234;
wire n_3280;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_3284;
wire n_2926;
wire n_1442;
wire n_2703;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1468;
wire n_1253;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_3212;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3159;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3250;
wire n_3029;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1972;
wire n_1178;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_1491;
wire n_931;
wire n_2628;
wire n_3219;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_3116;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_990;
wire n_1623;
wire n_1903;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_976;
wire n_909;
wire n_1392;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_3127;
wire n_1731;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_3052;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3179;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_3262;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_3171;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3246;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_2327;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2975;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_3118;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_3286;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_2075;
wire n_1726;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1377;
wire n_1614;
wire n_1162;
wire n_2031;
wire n_3260;
wire n_2118;
wire n_1740;
wire n_3222;
wire n_1602;
wire n_3139;
wire n_2853;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3035;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_2379;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_1708;
wire n_3085;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_1711;
wire n_1219;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2508;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_3151;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_3024;
wire n_2772;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_2893;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_1867;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_2958;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3097;
wire n_876;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_3173;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_1526;
wire n_2991;
wire n_1305;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_2905;
wire n_2884;
wire n_3167;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_3110;
wire n_1321;
wire n_3050;
wire n_3157;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3129;
wire n_1556;
wire n_1561;
wire n_2720;
wire n_2412;
wire n_3107;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_2936;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_2170;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_3236;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_3291;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_3184;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2796;
wire n_2173;
wire n_2715;
wire n_3206;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_914;
wire n_1116;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_1197;
wire n_3011;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_2647;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_2401;
wire n_2935;
wire n_889;
wire n_3255;
wire n_1549;
wire n_1066;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_911;
wire n_2658;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_3243;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_3117;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_3101;
wire n_918;
wire n_1968;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1803;
wire n_1444;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3241;
wire n_1157;
wire n_1584;
wire n_1664;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_2938;
wire n_1612;
wire n_2498;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_2600;
wire n_3092;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_2951;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3259;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_3292;
wire n_2872;
wire n_2126;
wire n_3109;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_3269;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3248;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_3091;
wire n_1024;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_2817;
wire n_2773;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_898;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3111;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_2569;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_2897;
wire n_1322;
wire n_3273;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_3155;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1865;
wire n_1710;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_1094;
wire n_2973;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_1754;
wire n_3146;
wire n_3038;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3188;
wire n_3001;
wire n_3232;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_2088;
wire n_3265;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3285;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_3203;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_2917;
wire n_3137;
wire n_2544;
wire n_3143;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_2430;
wire n_2504;
wire n_910;
wire n_1410;
wire n_939;
wire n_2297;
wire n_3094;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_2957;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_1638;
wire n_3071;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_1946;
wire n_2148;
wire n_933;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_3196;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_3293;
wire n_1683;
wire n_1229;
wire n_2582;
wire n_3228;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_3149;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3202;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_2573;
wire n_2940;
wire n_2336;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_1582;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx1_ASAP7_75t_L g871 ( 
.A(n_436),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_842),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_518),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_302),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_652),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_785),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_361),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_259),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_799),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_484),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_181),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_331),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_771),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_729),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_128),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_741),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_716),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_735),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_265),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_411),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_222),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_776),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_686),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_736),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_768),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_210),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_566),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_712),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_211),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_77),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_755),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_206),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_225),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_806),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_839),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_163),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_589),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_247),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_43),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_788),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_200),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_696),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_781),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_493),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_73),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_127),
.Y(n_916)
);

BUFx10_ASAP7_75t_L g917 ( 
.A(n_852),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_773),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_277),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_574),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_733),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_831),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_861),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_547),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_730),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_866),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_858),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_837),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_300),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_378),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_684),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_144),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_568),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_163),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_751),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_663),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_216),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_460),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_763),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_526),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_845),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_779),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_219),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_85),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_195),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_176),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_680),
.Y(n_947)
);

BUFx5_ASAP7_75t_L g948 ( 
.A(n_105),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_691),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_109),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_505),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_424),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_347),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_580),
.Y(n_954)
);

CKINVDCx16_ASAP7_75t_R g955 ( 
.A(n_550),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_29),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_479),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_122),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_333),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_843),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_570),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_406),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_556),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_827),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_724),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_850),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_644),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_816),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_796),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_824),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_300),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_490),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_371),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_129),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_297),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_48),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_789),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_75),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_77),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_708),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_737),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_75),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_523),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_835),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_502),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_107),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_298),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_812),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_140),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_86),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_471),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_772),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_761),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_766),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_726),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_819),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_519),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_769),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_725),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_164),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_195),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_753),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_145),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_511),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_868),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_473),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_175),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_156),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_299),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_807),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_397),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_854),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_157),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_863),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_36),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_79),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_767),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_834),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_321),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_53),
.Y(n_1020)
);

CKINVDCx16_ASAP7_75t_R g1021 ( 
.A(n_855),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_190),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_110),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_853),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_156),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_88),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_606),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_365),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_744),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_247),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_790),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_141),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_22),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_818),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_172),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_758),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_804),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_780),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_711),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_829),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_358),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_815),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_236),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_793),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_412),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_759),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_169),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_821),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_699),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_616),
.Y(n_1050)
);

BUFx8_ASAP7_75t_SL g1051 ( 
.A(n_100),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_244),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_739),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_584),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_206),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_430),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_817),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_727),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_814),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_757),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_693),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_404),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_721),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_577),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_222),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_538),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_337),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_336),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_634),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_597),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_392),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_862),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_69),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_354),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_340),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_116),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_591),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_22),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_588),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_101),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_347),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_667),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_742),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_743),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_469),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_389),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_402),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_366),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_784),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_344),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_185),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_10),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_851),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_625),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_381),
.Y(n_1095)
);

INVxp67_ASAP7_75t_SL g1096 ( 
.A(n_709),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_98),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_676),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_315),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_326),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_8),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_148),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_162),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_801),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_694),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_552),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_202),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_857),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_803),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_865),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_168),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_823),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_534),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_745),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_841),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_645),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_169),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_856),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_740),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_797),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_825),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_221),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_452),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_96),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_472),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_846),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_764),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_555),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_718),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_467),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_353),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_349),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_277),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_400),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_601),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_160),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_93),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_549),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_661),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_706),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_701),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_371),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_543),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_791),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_777),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_323),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_783),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_125),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_475),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_609),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_707),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_867),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_860),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_808),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_153),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_507),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_762),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_828),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_655),
.Y(n_1159)
);

CKINVDCx16_ASAP7_75t_R g1160 ( 
.A(n_198),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_388),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_836),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_416),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_438),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_732),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_646),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_160),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_295),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_139),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_159),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_765),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_723),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_623),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_127),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_398),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_420),
.Y(n_1176)
);

BUFx5_ASAP7_75t_L g1177 ( 
.A(n_654),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_722),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_702),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_328),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_391),
.Y(n_1181)
);

CKINVDCx16_ASAP7_75t_R g1182 ( 
.A(n_794),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_715),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_802),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_315),
.Y(n_1185)
);

CKINVDCx16_ASAP7_75t_R g1186 ( 
.A(n_838),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_176),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_44),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_343),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_592),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_223),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_713),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_175),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_787),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_809),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_10),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_542),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_197),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_232),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_464),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_669),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_704),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_775),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_599),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_847),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_756),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_458),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_426),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_774),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_626),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_240),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_752),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_291),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_849),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_810),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_323),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_778),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_782),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_714),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_826),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_562),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_335),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_805),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_754),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_848),
.Y(n_1225)
);

CKINVDCx16_ASAP7_75t_R g1226 ( 
.A(n_747),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_524),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_338),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_710),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_728),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_445),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_486),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_428),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_832),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_859),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_172),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_413),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_492),
.Y(n_1238)
);

CKINVDCx14_ASAP7_75t_R g1239 ( 
.A(n_62),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_582),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_404),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_426),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_734),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_864),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_750),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_705),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_330),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_191),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_365),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_811),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_792),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_700),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_113),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_820),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_446),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_703),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_638),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_717),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_760),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_738),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_659),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_406),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_731),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_313),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_605),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_572),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_258),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_456),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_800),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_786),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_795),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_813),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_263),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_749),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_504),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_770),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_840),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_688),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_254),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_719),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_67),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_361),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_116),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_396),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_202),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_383),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_40),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_191),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_746),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_187),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_844),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_379),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_830),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_405),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_720),
.Y(n_1295)
);

BUFx10_ASAP7_75t_L g1296 ( 
.A(n_262),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_273),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_341),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_869),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_748),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_42),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_675),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_132),
.Y(n_1303)
);

CKINVDCx16_ASAP7_75t_R g1304 ( 
.A(n_668),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_161),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_273),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_822),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_798),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_197),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_474),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_833),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_328),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_612),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_915),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_915),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_948),
.Y(n_1316)
);

INVxp67_ASAP7_75t_L g1317 ( 
.A(n_874),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_948),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_948),
.Y(n_1319)
);

INVxp33_ASAP7_75t_L g1320 ( 
.A(n_1292),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_948),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_948),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1239),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_948),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1051),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_891),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_909),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1160),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_886),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_877),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_907),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_878),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_900),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_937),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_946),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_955),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_909),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_953),
.Y(n_1338)
);

INVxp67_ASAP7_75t_SL g1339 ( 
.A(n_909),
.Y(n_1339)
);

CKINVDCx16_ASAP7_75t_R g1340 ( 
.A(n_1021),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_918),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_925),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_1015),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_956),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_962),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1015),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_936),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_1015),
.Y(n_1348)
);

CKINVDCx16_ASAP7_75t_R g1349 ( 
.A(n_1182),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_938),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_975),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_987),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_967),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1001),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1003),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_885),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1097),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1011),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_977),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_984),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_996),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1013),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1016),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_997),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1025),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1026),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1129),
.Y(n_1367)
);

CKINVDCx14_ASAP7_75t_R g1368 ( 
.A(n_917),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1103),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1028),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1032),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1033),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1041),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1166),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1047),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1055),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1062),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1266),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1065),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1074),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1081),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1100),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_881),
.Y(n_1383)
);

INVxp33_ASAP7_75t_SL g1384 ( 
.A(n_882),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1132),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1317),
.A2(n_950),
.B1(n_982),
.B2(n_916),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1339),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1356),
.B(n_1309),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1327),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1337),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1318),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1343),
.B(n_1346),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1336),
.A2(n_1122),
.B1(n_1078),
.B2(n_1073),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1326),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1329),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1348),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1384),
.B(n_904),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1316),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1319),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1368),
.B(n_1186),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1320),
.B(n_1226),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1369),
.B(n_949),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1314),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1315),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1321),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1322),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1324),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1330),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1357),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1332),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1369),
.B(n_1269),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1340),
.A2(n_1170),
.B1(n_989),
.B2(n_1304),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1331),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1349),
.B(n_917),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1333),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1328),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1334),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1335),
.B(n_871),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1338),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1344),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1345),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1351),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1352),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1383),
.A2(n_1030),
.B1(n_1117),
.B2(n_1076),
.Y(n_1424)
);

XNOR2xp5_ASAP7_75t_L g1425 ( 
.A(n_1342),
.B(n_889),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1354),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1355),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1358),
.B(n_1296),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1347),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1362),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1363),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1365),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1341),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1366),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1323),
.B(n_979),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1370),
.B(n_873),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1371),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1372),
.B(n_1296),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1373),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1375),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1350),
.B(n_888),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1367),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1376),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1377),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1379),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1374),
.A2(n_1169),
.B1(n_1087),
.B2(n_896),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1394),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1406),
.B(n_1380),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1445),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1428),
.B(n_1381),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1409),
.Y(n_1451)
);

BUFx4f_ASAP7_75t_L g1452 ( 
.A(n_1416),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1391),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1389),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1403),
.Y(n_1455)
);

INVxp67_ASAP7_75t_SL g1456 ( 
.A(n_1392),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1404),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1430),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1397),
.B(n_1378),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1413),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1395),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1432),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1401),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1399),
.A2(n_899),
.B1(n_1071),
.B2(n_959),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1434),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1442),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1408),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1389),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1398),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1438),
.B(n_1382),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1390),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1410),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1426),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1424),
.A2(n_929),
.B1(n_952),
.B2(n_906),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1400),
.B(n_890),
.Y(n_1475)
);

NAND2xp33_ASAP7_75t_L g1476 ( 
.A(n_1398),
.B(n_1405),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1415),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1446),
.B(n_1388),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1417),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1419),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1387),
.B(n_1385),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1426),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1427),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1390),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1429),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1441),
.A2(n_1096),
.B(n_1310),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1420),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1421),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1386),
.A2(n_943),
.B1(n_1133),
.B2(n_932),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1427),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1407),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1431),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1437),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1439),
.A2(n_1080),
.B1(n_1142),
.B2(n_1137),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1439),
.B(n_902),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1396),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1422),
.B(n_1148),
.Y(n_1497)
);

INVx4_ASAP7_75t_L g1498 ( 
.A(n_1440),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1440),
.B(n_903),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1423),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1443),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1444),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1435),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1418),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1436),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1402),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1411),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1433),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1414),
.B(n_1029),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1412),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1425),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1393),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1403),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1409),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1403),
.Y(n_1515)
);

BUFx8_ASAP7_75t_SL g1516 ( 
.A(n_1395),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1409),
.Y(n_1517)
);

OAI21xp33_ASAP7_75t_SL g1518 ( 
.A1(n_1397),
.A2(n_1196),
.B(n_1161),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1409),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1409),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1466),
.B(n_1353),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1460),
.B(n_1359),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1456),
.B(n_910),
.Y(n_1523)
);

OAI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1506),
.A2(n_911),
.B1(n_919),
.B2(n_908),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1504),
.A2(n_1180),
.B1(n_1236),
.B2(n_1211),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1447),
.B(n_1463),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1507),
.B(n_1360),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1452),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1516),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1461),
.B(n_1361),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1508),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1508),
.B(n_1364),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1503),
.B(n_1325),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1485),
.B(n_1189),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1511),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1496),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1451),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1459),
.B(n_930),
.Y(n_1538)
);

AO22x2_ASAP7_75t_L g1539 ( 
.A1(n_1512),
.A2(n_1216),
.B1(n_1233),
.B2(n_1213),
.Y(n_1539)
);

A2O1A1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1505),
.A2(n_1264),
.B(n_1279),
.C(n_1237),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1449),
.B(n_1154),
.Y(n_1541)
);

AND2x6_ASAP7_75t_L g1542 ( 
.A(n_1510),
.B(n_1282),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1518),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1467),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1514),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1450),
.B(n_1283),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1473),
.B(n_1482),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1509),
.B(n_1305),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1472),
.Y(n_1549)
);

NAND2x1p5_ASAP7_75t_L g1550 ( 
.A(n_1498),
.B(n_1204),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1477),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1483),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1483),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1470),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1490),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1489),
.A2(n_944),
.B1(n_1043),
.B2(n_971),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1490),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1469),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1469),
.B(n_934),
.Y(n_1559)
);

AO22x2_ASAP7_75t_L g1560 ( 
.A1(n_1478),
.A2(n_1290),
.B1(n_1297),
.B2(n_1286),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1517),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1501),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1479),
.Y(n_1563)
);

OAI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1474),
.A2(n_958),
.B1(n_973),
.B2(n_945),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1500),
.B(n_1312),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1480),
.Y(n_1566)
);

AO22x2_ASAP7_75t_L g1567 ( 
.A1(n_1475),
.A2(n_1281),
.B1(n_1303),
.B2(n_1242),
.Y(n_1567)
);

INVx4_ASAP7_75t_L g1568 ( 
.A(n_1497),
.Y(n_1568)
);

INVx5_ASAP7_75t_L g1569 ( 
.A(n_1497),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1487),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1488),
.B(n_974),
.Y(n_1571)
);

INVx6_ASAP7_75t_L g1572 ( 
.A(n_1494),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1454),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1492),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1481),
.B(n_976),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1493),
.B(n_978),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1455),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1457),
.B(n_986),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1468),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1502),
.B(n_990),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1513),
.B(n_1000),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1515),
.B(n_1458),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1491),
.B(n_1007),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1495),
.B(n_1008),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1462),
.B(n_1009),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1499),
.B(n_960),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1465),
.B(n_1019),
.Y(n_1587)
);

AO22x2_ASAP7_75t_L g1588 ( 
.A1(n_1520),
.A2(n_968),
.B1(n_1002),
.B2(n_895),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1486),
.B(n_1298),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1453),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1448),
.B(n_1020),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1519),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1471),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1484),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1476),
.B(n_1022),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1464),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1466),
.B(n_1023),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1447),
.B(n_1035),
.Y(n_1598)
);

INVx8_ASAP7_75t_L g1599 ( 
.A(n_1516),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1508),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1456),
.B(n_1045),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1516),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1485),
.A2(n_1056),
.B1(n_1067),
.B2(n_1052),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1496),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1451),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1456),
.B(n_1068),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1447),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1466),
.B(n_1075),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1461),
.B(n_1086),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1505),
.A2(n_1090),
.B1(n_1091),
.B2(n_1088),
.Y(n_1610)
);

AO22x2_ASAP7_75t_L g1611 ( 
.A1(n_1512),
.A2(n_970),
.B1(n_1058),
.B2(n_933),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1456),
.B(n_1092),
.Y(n_1612)
);

NAND3xp33_ASAP7_75t_L g1613 ( 
.A(n_1506),
.B(n_1099),
.C(n_1095),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1447),
.B(n_1306),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1456),
.B(n_1101),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1518),
.A2(n_1111),
.B1(n_1124),
.B2(n_1107),
.C(n_1102),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1508),
.B(n_1287),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1447),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1466),
.B(n_1131),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1466),
.B(n_1134),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1447),
.B(n_1136),
.Y(n_1621)
);

NOR2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1460),
.B(n_1191),
.Y(n_1622)
);

AOI22x1_ASAP7_75t_L g1623 ( 
.A1(n_1505),
.A2(n_1155),
.B1(n_1163),
.B2(n_1146),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1516),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1516),
.Y(n_1625)
);

INVx8_ASAP7_75t_L g1626 ( 
.A(n_1516),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1516),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1447),
.Y(n_1628)
);

INVx6_ASAP7_75t_L g1629 ( 
.A(n_1466),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1516),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1496),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1516),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1516),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1447),
.B(n_1301),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1447),
.B(n_1167),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1466),
.B(n_1168),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1447),
.B(n_1174),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1496),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1456),
.B(n_1175),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1456),
.B(n_1176),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1461),
.B(n_1181),
.Y(n_1641)
);

NAND2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1452),
.B(n_894),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1451),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1456),
.B(n_1185),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1447),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1451),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1466),
.B(n_1187),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1456),
.B(n_1188),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1496),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1452),
.B(n_926),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1466),
.B(n_1193),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1516),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_R g1653 ( 
.A(n_1485),
.B(n_872),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1496),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1505),
.A2(n_1199),
.B1(n_1208),
.B2(n_1198),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1496),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1496),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1451),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1516),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1456),
.B(n_1222),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1569),
.B(n_875),
.Y(n_1661)
);

INVxp67_ASAP7_75t_SL g1662 ( 
.A(n_1531),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1537),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1628),
.B(n_1228),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1569),
.B(n_1554),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1536),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1629),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1530),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1601),
.A2(n_880),
.B(n_879),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1604),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1548),
.A2(n_1247),
.B1(n_1248),
.B2(n_1241),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1552),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1631),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1599),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1545),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1607),
.B(n_1249),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1638),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1527),
.A2(n_884),
.B1(n_893),
.B2(n_876),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1543),
.A2(n_905),
.B1(n_912),
.B2(n_898),
.Y(n_1679)
);

BUFx8_ASAP7_75t_L g1680 ( 
.A(n_1602),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1521),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1538),
.A2(n_957),
.B1(n_965),
.B2(n_940),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1560),
.A2(n_1262),
.B1(n_1267),
.B2(n_1253),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1532),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1624),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1561),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1553),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1649),
.Y(n_1688)
);

INVx5_ASAP7_75t_L g1689 ( 
.A(n_1625),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1654),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1618),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1542),
.A2(n_1284),
.B1(n_1285),
.B2(n_1273),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1656),
.Y(n_1693)
);

AND2x2_ASAP7_75t_SL g1694 ( 
.A(n_1522),
.B(n_897),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1657),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1523),
.B(n_1288),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1660),
.A2(n_983),
.B(n_980),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1645),
.B(n_1568),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1575),
.B(n_1294),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1526),
.B(n_1024),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_1627),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1598),
.B(n_0),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1544),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1614),
.A2(n_1039),
.B1(n_1046),
.B2(n_1027),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1606),
.B(n_1048),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1534),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1556),
.A2(n_1082),
.B1(n_1093),
.B2(n_1059),
.Y(n_1707)
);

NOR2xp67_ASAP7_75t_L g1708 ( 
.A(n_1528),
.B(n_1110),
.Y(n_1708)
);

INVx4_ASAP7_75t_L g1709 ( 
.A(n_1626),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1600),
.B(n_1157),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1605),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1549),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1643),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1612),
.B(n_1615),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1551),
.Y(n_1715)
);

O2A1O1Ixp33_ASAP7_75t_L g1716 ( 
.A1(n_1564),
.A2(n_1143),
.B(n_1158),
.C(n_1127),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1563),
.A2(n_1162),
.B(n_1165),
.C(n_1159),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1566),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1555),
.B(n_1171),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1558),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1639),
.B(n_883),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1640),
.B(n_1179),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1570),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1574),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1621),
.B(n_0),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1644),
.B(n_1183),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1653),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1648),
.B(n_1192),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1557),
.B(n_1205),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1533),
.B(n_1206),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1577),
.B(n_1210),
.Y(n_1731)
);

AND2x6_ASAP7_75t_L g1732 ( 
.A(n_1596),
.B(n_1214),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1609),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1550),
.Y(n_1734)
);

BUFx12f_ASAP7_75t_SL g1735 ( 
.A(n_1630),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1547),
.B(n_1221),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1634),
.A2(n_1256),
.B1(n_1260),
.B2(n_1246),
.Y(n_1737)
);

NOR3xp33_ASAP7_75t_L g1738 ( 
.A(n_1616),
.B(n_1280),
.C(n_1263),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1582),
.B(n_1291),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1641),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1529),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1576),
.B(n_887),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1637),
.A2(n_901),
.B1(n_913),
.B2(n_892),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1591),
.A2(n_1571),
.B1(n_1581),
.B2(n_1578),
.Y(n_1744)
);

BUFx3_ASAP7_75t_L g1745 ( 
.A(n_1632),
.Y(n_1745)
);

NOR2x1p5_ASAP7_75t_L g1746 ( 
.A(n_1633),
.B(n_1108),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1635),
.B(n_1),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1603),
.B(n_1),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1646),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1572),
.B(n_914),
.Y(n_1750)
);

INVx4_ASAP7_75t_L g1751 ( 
.A(n_1652),
.Y(n_1751)
);

AND3x1_ASAP7_75t_L g1752 ( 
.A(n_1540),
.B(n_942),
.C(n_939),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1658),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1659),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1585),
.B(n_920),
.Y(n_1755)
);

BUFx3_ASAP7_75t_L g1756 ( 
.A(n_1573),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1541),
.Y(n_1757)
);

OAI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1613),
.A2(n_1070),
.B(n_1060),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1587),
.B(n_921),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1562),
.B(n_922),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1597),
.B(n_923),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1579),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1546),
.B(n_924),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1535),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1542),
.A2(n_1258),
.B1(n_1308),
.B2(n_1251),
.Y(n_1765)
);

INVx5_ASAP7_75t_L g1766 ( 
.A(n_1586),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1608),
.Y(n_1767)
);

INVx5_ASAP7_75t_L g1768 ( 
.A(n_1619),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1622),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1611),
.A2(n_1218),
.B1(n_1254),
.B2(n_1089),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_R g1771 ( 
.A(n_1620),
.B(n_927),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1590),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1642),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1592),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1583),
.B(n_928),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1593),
.Y(n_1776)
);

BUFx6f_ASAP7_75t_SL g1777 ( 
.A(n_1636),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1594),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1584),
.A2(n_935),
.B1(n_941),
.B2(n_931),
.Y(n_1779)
);

INVx3_ASAP7_75t_L g1780 ( 
.A(n_1650),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1588),
.Y(n_1781)
);

BUFx3_ASAP7_75t_L g1782 ( 
.A(n_1647),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1524),
.B(n_947),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1651),
.B(n_951),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1565),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1589),
.B(n_961),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1539),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1595),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1525),
.B(n_963),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1567),
.A2(n_964),
.B1(n_1018),
.B2(n_954),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1559),
.Y(n_1791)
);

INVx2_ASAP7_75t_SL g1792 ( 
.A(n_1580),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1623),
.Y(n_1793)
);

INVx5_ASAP7_75t_L g1794 ( 
.A(n_1617),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1610),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1655),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1569),
.B(n_966),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1537),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1569),
.B(n_2),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1560),
.A2(n_964),
.B1(n_1018),
.B2(n_954),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1554),
.B(n_969),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1529),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1536),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1569),
.B(n_2),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_L g1805 ( 
.A(n_1531),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1569),
.B(n_972),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1554),
.B(n_981),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_1530),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1569),
.B(n_985),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1537),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1569),
.B(n_988),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1554),
.B(n_991),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1554),
.B(n_992),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1536),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1527),
.B(n_3),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1537),
.Y(n_1816)
);

OR2x2_ASAP7_75t_SL g1817 ( 
.A(n_1629),
.B(n_954),
.Y(n_1817)
);

INVx2_ASAP7_75t_SL g1818 ( 
.A(n_1629),
.Y(n_1818)
);

NAND2x1p5_ASAP7_75t_L g1819 ( 
.A(n_1600),
.B(n_964),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1569),
.B(n_993),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1531),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1537),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1537),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1569),
.B(n_994),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1629),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1537),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_SL g1827 ( 
.A1(n_1616),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.C(n_6),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1554),
.B(n_995),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1629),
.Y(n_1829)
);

AND2x6_ASAP7_75t_L g1830 ( 
.A(n_1528),
.B(n_1018),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1569),
.B(n_998),
.Y(n_1831)
);

AOI21xp33_ASAP7_75t_L g1832 ( 
.A1(n_1548),
.A2(n_1004),
.B(n_999),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1554),
.B(n_1005),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_SL g1834 ( 
.A1(n_1548),
.A2(n_1010),
.B1(n_1012),
.B2(n_1006),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1556),
.A2(n_1017),
.B1(n_1031),
.B2(n_1014),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1536),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1536),
.Y(n_1837)
);

BUFx4f_ASAP7_75t_L g1838 ( 
.A(n_1602),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1536),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1536),
.Y(n_1840)
);

AND2x4_ASAP7_75t_L g1841 ( 
.A(n_1569),
.B(n_4),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1569),
.B(n_1034),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1537),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1628),
.B(n_5),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1560),
.A2(n_1255),
.B1(n_1302),
.B2(n_1115),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_SL g1846 ( 
.A(n_1529),
.B(n_1037),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1548),
.B(n_1036),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1629),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1554),
.B(n_1038),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1560),
.A2(n_1255),
.B1(n_1302),
.B2(n_1115),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1628),
.Y(n_1851)
);

O2A1O1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1548),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_1852)
);

INVx2_ASAP7_75t_SL g1853 ( 
.A(n_1629),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1536),
.Y(n_1854)
);

BUFx3_ASAP7_75t_L g1855 ( 
.A(n_1629),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1700),
.B(n_7),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1666),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1847),
.B(n_9),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_SL g1859 ( 
.A(n_1735),
.B(n_1299),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1829),
.B(n_9),
.Y(n_1860)
);

BUFx3_ASAP7_75t_L g1861 ( 
.A(n_1855),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1667),
.B(n_11),
.Y(n_1862)
);

OR2x6_ASAP7_75t_L g1863 ( 
.A(n_1818),
.B(n_1115),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1795),
.B(n_11),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1694),
.B(n_1733),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1707),
.A2(n_1042),
.B1(n_1044),
.B2(n_1040),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1741),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1732),
.A2(n_1302),
.B1(n_1255),
.B2(n_1177),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1772),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1714),
.A2(n_1274),
.B(n_1272),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1750),
.B(n_12),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1851),
.B(n_12),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1796),
.B(n_13),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1854),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1670),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_1825),
.Y(n_1876)
);

CKINVDCx20_ASAP7_75t_R g1877 ( 
.A(n_1680),
.Y(n_1877)
);

BUFx2_ASAP7_75t_L g1878 ( 
.A(n_1672),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1673),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1848),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1698),
.B(n_1276),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1691),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1677),
.B(n_13),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1688),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1853),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1690),
.B(n_1693),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1740),
.B(n_14),
.Y(n_1887)
);

INVx1_ASAP7_75t_SL g1888 ( 
.A(n_1764),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1774),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1695),
.Y(n_1890)
);

INVx4_ASAP7_75t_L g1891 ( 
.A(n_1689),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1703),
.B(n_14),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1732),
.A2(n_1177),
.B1(n_1050),
.B2(n_1053),
.Y(n_1893)
);

A2O1A1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1697),
.A2(n_1054),
.B(n_1105),
.C(n_1077),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1712),
.Y(n_1895)
);

INVxp67_ASAP7_75t_SL g1896 ( 
.A(n_1805),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1663),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1715),
.B(n_15),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1706),
.B(n_1049),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1808),
.B(n_1664),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1732),
.A2(n_1177),
.B1(n_1061),
.B2(n_1063),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1718),
.B(n_15),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1681),
.B(n_16),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1723),
.B(n_16),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1815),
.B(n_17),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1702),
.B(n_17),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1744),
.B(n_1057),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1724),
.B(n_18),
.Y(n_1908)
);

NAND3xp33_ASAP7_75t_L g1909 ( 
.A(n_1783),
.B(n_1066),
.C(n_1064),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1768),
.B(n_18),
.Y(n_1910)
);

NOR2xp67_ASAP7_75t_L g1911 ( 
.A(n_1768),
.B(n_1069),
.Y(n_1911)
);

AO22x1_ASAP7_75t_L g1912 ( 
.A1(n_1748),
.A2(n_1079),
.B1(n_1083),
.B2(n_1072),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1803),
.B(n_19),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1675),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1802),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1814),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1686),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1727),
.B(n_1300),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1683),
.A2(n_1177),
.B1(n_1085),
.B2(n_1094),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1711),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1836),
.A2(n_1313),
.B1(n_1123),
.B2(n_1140),
.Y(n_1921)
);

NOR3xp33_ASAP7_75t_L g1922 ( 
.A(n_1671),
.B(n_1125),
.C(n_1112),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1837),
.B(n_19),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1839),
.B(n_20),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1840),
.B(n_20),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1713),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1763),
.B(n_21),
.Y(n_1927)
);

BUFx3_ASAP7_75t_L g1928 ( 
.A(n_1674),
.Y(n_1928)
);

OAI221xp5_ASAP7_75t_L g1929 ( 
.A1(n_1678),
.A2(n_1104),
.B1(n_1106),
.B2(n_1098),
.C(n_1084),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1749),
.Y(n_1930)
);

BUFx2_ASAP7_75t_L g1931 ( 
.A(n_1782),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1725),
.B(n_1747),
.Y(n_1932)
);

AO22x1_ASAP7_75t_L g1933 ( 
.A1(n_1766),
.A2(n_1113),
.B1(n_1114),
.B2(n_1109),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1696),
.B(n_21),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1753),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1798),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1739),
.B(n_23),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1668),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1810),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1767),
.B(n_23),
.Y(n_1940)
);

NOR2xp67_ASAP7_75t_L g1941 ( 
.A(n_1709),
.B(n_1116),
.Y(n_1941)
);

BUFx3_ASAP7_75t_L g1942 ( 
.A(n_1745),
.Y(n_1942)
);

INVx3_ASAP7_75t_L g1943 ( 
.A(n_1751),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1730),
.B(n_24),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1816),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1822),
.Y(n_1946)
);

INVxp67_ASAP7_75t_L g1947 ( 
.A(n_1844),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1805),
.B(n_1118),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1823),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1821),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1781),
.B(n_24),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1788),
.B(n_1801),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1826),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1682),
.A2(n_1120),
.B1(n_1121),
.B2(n_1119),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1843),
.Y(n_1955)
);

INVxp67_ASAP7_75t_SL g1956 ( 
.A(n_1821),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1776),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1778),
.Y(n_1958)
);

OAI31xp33_ASAP7_75t_SL g1959 ( 
.A1(n_1834),
.A2(n_1832),
.A3(n_1793),
.B(n_1721),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1835),
.A2(n_1128),
.B1(n_1130),
.B2(n_1126),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1787),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1731),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1799),
.B(n_25),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1785),
.Y(n_1964)
);

AND3x1_ASAP7_75t_SL g1965 ( 
.A(n_1746),
.B(n_25),
.C(n_26),
.Y(n_1965)
);

BUFx4f_ASAP7_75t_L g1966 ( 
.A(n_1685),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1807),
.B(n_26),
.Y(n_1967)
);

INVx4_ASAP7_75t_L g1968 ( 
.A(n_1689),
.Y(n_1968)
);

OR2x6_ASAP7_75t_L g1969 ( 
.A(n_1685),
.B(n_27),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1791),
.Y(n_1970)
);

BUFx3_ASAP7_75t_L g1971 ( 
.A(n_1838),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1819),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1756),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1687),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1812),
.B(n_27),
.Y(n_1975)
);

INVx2_ASAP7_75t_SL g1976 ( 
.A(n_1701),
.Y(n_1976)
);

INVx5_ASAP7_75t_L g1977 ( 
.A(n_1701),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1679),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1804),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1841),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1720),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1813),
.B(n_28),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1792),
.B(n_28),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1771),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1828),
.B(n_29),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1684),
.B(n_30),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1833),
.B(n_30),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1754),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1754),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1849),
.B(n_31),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1762),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1766),
.B(n_1135),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1705),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1722),
.Y(n_1994)
);

BUFx4f_ASAP7_75t_L g1995 ( 
.A(n_1830),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1726),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1728),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1699),
.B(n_31),
.Y(n_1998)
);

INVxp67_ASAP7_75t_L g1999 ( 
.A(n_1882),
.Y(n_1999)
);

INVx5_ASAP7_75t_L g2000 ( 
.A(n_1891),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1997),
.B(n_1784),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1900),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1878),
.B(n_1817),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1861),
.B(n_1662),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1877),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1932),
.B(n_1736),
.Y(n_2006)
);

BUFx8_ASAP7_75t_L g2007 ( 
.A(n_1984),
.Y(n_2007)
);

CKINVDCx6p67_ASAP7_75t_R g2008 ( 
.A(n_1971),
.Y(n_2008)
);

O2A1O1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1856),
.A2(n_1716),
.B(n_1852),
.C(n_1738),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1928),
.B(n_1773),
.Y(n_2010)
);

NOR2xp67_ASAP7_75t_SL g2011 ( 
.A(n_1867),
.B(n_1769),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1857),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1942),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1950),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1974),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1907),
.A2(n_1737),
.B1(n_1704),
.B2(n_1779),
.Y(n_2016)
);

OAI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1858),
.A2(n_1775),
.B1(n_1742),
.B2(n_1743),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1874),
.Y(n_2018)
);

OAI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_1959),
.A2(n_1692),
.B1(n_1846),
.B2(n_1759),
.C(n_1755),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_1950),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1875),
.Y(n_2021)
);

BUFx6f_ASAP7_75t_L g2022 ( 
.A(n_1966),
.Y(n_2022)
);

AND2x4_ASAP7_75t_L g2023 ( 
.A(n_1876),
.B(n_1780),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1977),
.Y(n_2024)
);

INVx3_ASAP7_75t_L g2025 ( 
.A(n_1968),
.Y(n_2025)
);

NAND2xp33_ASAP7_75t_L g2026 ( 
.A(n_1922),
.B(n_1830),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_SL g2027 ( 
.A1(n_1978),
.A2(n_1786),
.B1(n_1777),
.B2(n_1661),
.Y(n_2027)
);

NAND2x1p5_ASAP7_75t_L g2028 ( 
.A(n_1977),
.B(n_1757),
.Y(n_2028)
);

BUFx8_ASAP7_75t_L g2029 ( 
.A(n_1988),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1952),
.B(n_1708),
.Y(n_2030)
);

BUFx2_ASAP7_75t_L g2031 ( 
.A(n_1931),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1988),
.Y(n_2032)
);

OR2x6_ASAP7_75t_L g2033 ( 
.A(n_1976),
.B(n_1734),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1915),
.Y(n_2034)
);

OR2x6_ASAP7_75t_L g2035 ( 
.A(n_1969),
.B(n_1665),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1872),
.B(n_1719),
.Y(n_2036)
);

INVx4_ASAP7_75t_L g2037 ( 
.A(n_1943),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1937),
.A2(n_1886),
.B(n_1967),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1879),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1884),
.Y(n_2040)
);

BUFx3_ASAP7_75t_L g2041 ( 
.A(n_1880),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1890),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1885),
.B(n_1794),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1869),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1895),
.Y(n_2045)
);

BUFx2_ASAP7_75t_L g2046 ( 
.A(n_1981),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1944),
.B(n_1865),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_SL g2048 ( 
.A(n_1995),
.B(n_1794),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1866),
.A2(n_1752),
.B1(n_1710),
.B2(n_1676),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1993),
.B(n_1770),
.Y(n_2050)
);

AND2x4_ASAP7_75t_L g2051 ( 
.A(n_1896),
.B(n_1729),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1975),
.A2(n_1760),
.B(n_1669),
.Y(n_2052)
);

OAI221xp5_ASAP7_75t_L g2053 ( 
.A1(n_1871),
.A2(n_1827),
.B1(n_1717),
.B2(n_1761),
.C(n_1765),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1889),
.Y(n_2054)
);

INVx4_ASAP7_75t_L g2055 ( 
.A(n_1989),
.Y(n_2055)
);

OR2x6_ASAP7_75t_L g2056 ( 
.A(n_1969),
.B(n_1910),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1956),
.B(n_1797),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1940),
.B(n_1758),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1916),
.Y(n_2059)
);

BUFx2_ASAP7_75t_L g2060 ( 
.A(n_1888),
.Y(n_2060)
);

INVx2_ASAP7_75t_SL g2061 ( 
.A(n_1973),
.Y(n_2061)
);

INVx3_ASAP7_75t_L g2062 ( 
.A(n_1991),
.Y(n_2062)
);

INVx1_ASAP7_75t_SL g2063 ( 
.A(n_1938),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1994),
.B(n_1800),
.Y(n_2064)
);

OAI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_1927),
.A2(n_1850),
.B1(n_1845),
.B2(n_1790),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1958),
.Y(n_2066)
);

BUFx12f_ASAP7_75t_L g2067 ( 
.A(n_1860),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1897),
.Y(n_2068)
);

CKINVDCx20_ASAP7_75t_R g2069 ( 
.A(n_1965),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1930),
.Y(n_2070)
);

INVx3_ASAP7_75t_L g2071 ( 
.A(n_1964),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1936),
.Y(n_2072)
);

AOI22xp33_ASAP7_75t_L g2073 ( 
.A1(n_1962),
.A2(n_1789),
.B1(n_1830),
.B2(n_1809),
.Y(n_2073)
);

INVx2_ASAP7_75t_SL g2074 ( 
.A(n_1979),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1914),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1996),
.B(n_1806),
.Y(n_2076)
);

CKINVDCx20_ASAP7_75t_R g2077 ( 
.A(n_1899),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1917),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1947),
.B(n_1811),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1980),
.B(n_1820),
.Y(n_2080)
);

AOI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1960),
.A2(n_1831),
.B1(n_1842),
.B2(n_1824),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1920),
.Y(n_2082)
);

AOI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_1912),
.A2(n_1139),
.B1(n_1141),
.B2(n_1138),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1939),
.Y(n_2084)
);

INVx1_ASAP7_75t_SL g2085 ( 
.A(n_1887),
.Y(n_2085)
);

BUFx2_ASAP7_75t_L g2086 ( 
.A(n_1863),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1945),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_1905),
.A2(n_1177),
.B1(n_1145),
.B2(n_1147),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_1863),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1963),
.B(n_32),
.Y(n_2090)
);

INVx4_ASAP7_75t_L g2091 ( 
.A(n_1862),
.Y(n_2091)
);

BUFx6f_ASAP7_75t_L g2092 ( 
.A(n_1926),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1970),
.B(n_32),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_1919),
.A2(n_1906),
.B1(n_1929),
.B2(n_1935),
.Y(n_2094)
);

CKINVDCx11_ASAP7_75t_R g2095 ( 
.A(n_1903),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1946),
.Y(n_2096)
);

INVx1_ASAP7_75t_SL g2097 ( 
.A(n_1983),
.Y(n_2097)
);

BUFx8_ASAP7_75t_SL g2098 ( 
.A(n_1986),
.Y(n_2098)
);

OAI221xp5_ASAP7_75t_L g2099 ( 
.A1(n_1998),
.A2(n_1150),
.B1(n_1231),
.B2(n_1219),
.C(n_1201),
.Y(n_2099)
);

NOR2x1_ASAP7_75t_SL g2100 ( 
.A(n_1864),
.B(n_1873),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1911),
.B(n_435),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1953),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1957),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_1881),
.B(n_1144),
.Y(n_2104)
);

HB1xp67_ASAP7_75t_L g2105 ( 
.A(n_1961),
.Y(n_2105)
);

O2A1O1Ixp5_ASAP7_75t_L g2106 ( 
.A1(n_1982),
.A2(n_1177),
.B(n_35),
.C(n_33),
.Y(n_2106)
);

OAI21x1_ASAP7_75t_L g2107 ( 
.A1(n_1985),
.A2(n_439),
.B(n_437),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1992),
.B(n_33),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1949),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1955),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1859),
.B(n_1149),
.Y(n_2111)
);

BUFx6f_ASAP7_75t_L g2112 ( 
.A(n_1972),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_1941),
.B(n_440),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_1883),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1951),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_1918),
.Y(n_2116)
);

OR2x6_ASAP7_75t_SL g2117 ( 
.A(n_1909),
.B(n_1151),
.Y(n_2117)
);

INVx1_ASAP7_75t_SL g2118 ( 
.A(n_1933),
.Y(n_2118)
);

BUFx6f_ASAP7_75t_L g2119 ( 
.A(n_1892),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1934),
.B(n_34),
.Y(n_2120)
);

CKINVDCx5p33_ASAP7_75t_R g2121 ( 
.A(n_1948),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1898),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1902),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1904),
.Y(n_2124)
);

NOR2xp67_ASAP7_75t_L g2125 ( 
.A(n_1987),
.B(n_441),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1908),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1913),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1923),
.Y(n_2128)
);

INVx2_ASAP7_75t_SL g2129 ( 
.A(n_1924),
.Y(n_2129)
);

NOR2x1_ASAP7_75t_SL g2130 ( 
.A(n_1925),
.B(n_34),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_1990),
.Y(n_2131)
);

BUFx3_ASAP7_75t_L g2132 ( 
.A(n_1954),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1921),
.Y(n_2133)
);

A2O1A1Ixp33_ASAP7_75t_L g2134 ( 
.A1(n_1894),
.A2(n_1153),
.B(n_1156),
.C(n_1152),
.Y(n_2134)
);

O2A1O1Ixp33_ASAP7_75t_L g2135 ( 
.A1(n_1870),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1868),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1893),
.Y(n_2137)
);

AOI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1901),
.A2(n_1172),
.B1(n_1173),
.B2(n_1164),
.Y(n_2138)
);

BUFx2_ASAP7_75t_L g2139 ( 
.A(n_1861),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1997),
.B(n_37),
.Y(n_2140)
);

A2O1A1Ixp33_ASAP7_75t_L g2141 ( 
.A1(n_1907),
.A2(n_1184),
.B(n_1190),
.C(n_1178),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1857),
.Y(n_2142)
);

AOI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_1907),
.A2(n_1195),
.B1(n_1197),
.B2(n_1194),
.Y(n_2143)
);

OAI21x1_ASAP7_75t_L g2144 ( 
.A1(n_2107),
.A2(n_443),
.B(n_442),
.Y(n_2144)
);

OAI21x1_ASAP7_75t_L g2145 ( 
.A1(n_2052),
.A2(n_447),
.B(n_444),
.Y(n_2145)
);

OAI21x1_ASAP7_75t_L g2146 ( 
.A1(n_2038),
.A2(n_449),
.B(n_448),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2002),
.B(n_38),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2105),
.B(n_2085),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2012),
.Y(n_2149)
);

BUFx2_ASAP7_75t_L g2150 ( 
.A(n_2031),
.Y(n_2150)
);

AOI22xp5_ASAP7_75t_L g2151 ( 
.A1(n_2016),
.A2(n_1202),
.B1(n_1203),
.B2(n_1200),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_2022),
.Y(n_2152)
);

CKINVDCx20_ASAP7_75t_R g2153 ( 
.A(n_2005),
.Y(n_2153)
);

OA21x2_ASAP7_75t_L g2154 ( 
.A1(n_2106),
.A2(n_1209),
.B(n_1207),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2044),
.Y(n_2155)
);

OAI21x1_ASAP7_75t_L g2156 ( 
.A1(n_2018),
.A2(n_451),
.B(n_450),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2021),
.B(n_38),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_2034),
.Y(n_2158)
);

INVx2_ASAP7_75t_SL g2159 ( 
.A(n_2029),
.Y(n_2159)
);

OAI21x1_ASAP7_75t_L g2160 ( 
.A1(n_2039),
.A2(n_454),
.B(n_453),
.Y(n_2160)
);

INVxp67_ASAP7_75t_SL g2161 ( 
.A(n_1999),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2040),
.Y(n_2162)
);

OAI21x1_ASAP7_75t_L g2163 ( 
.A1(n_2042),
.A2(n_457),
.B(n_455),
.Y(n_2163)
);

OA21x2_ASAP7_75t_L g2164 ( 
.A1(n_2115),
.A2(n_1215),
.B(n_1212),
.Y(n_2164)
);

AO21x2_ASAP7_75t_L g2165 ( 
.A1(n_2100),
.A2(n_1220),
.B(n_1217),
.Y(n_2165)
);

OA21x2_ASAP7_75t_L g2166 ( 
.A1(n_2120),
.A2(n_1224),
.B(n_1223),
.Y(n_2166)
);

OA21x2_ASAP7_75t_L g2167 ( 
.A1(n_2122),
.A2(n_1227),
.B(n_1225),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2054),
.Y(n_2168)
);

NAND2x1p5_ASAP7_75t_L g2169 ( 
.A(n_2024),
.B(n_459),
.Y(n_2169)
);

NOR2xp67_ASAP7_75t_L g2170 ( 
.A(n_2000),
.B(n_461),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2045),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2059),
.Y(n_2172)
);

OR2x2_ASAP7_75t_L g2173 ( 
.A(n_2142),
.B(n_39),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2068),
.Y(n_2174)
);

OAI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_2017),
.A2(n_2009),
.B(n_2019),
.Y(n_2175)
);

OAI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2132),
.A2(n_1230),
.B1(n_1232),
.B2(n_1229),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2066),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2001),
.B(n_39),
.Y(n_2178)
);

CKINVDCx11_ASAP7_75t_R g2179 ( 
.A(n_2022),
.Y(n_2179)
);

OAI22xp33_ASAP7_75t_SL g2180 ( 
.A1(n_2030),
.A2(n_1235),
.B1(n_1238),
.B2(n_1234),
.Y(n_2180)
);

OAI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2143),
.A2(n_1243),
.B1(n_1244),
.B2(n_1240),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2139),
.Y(n_2182)
);

BUFx10_ASAP7_75t_L g2183 ( 
.A(n_2014),
.Y(n_2183)
);

BUFx2_ASAP7_75t_SL g2184 ( 
.A(n_2000),
.Y(n_2184)
);

INVx2_ASAP7_75t_SL g2185 ( 
.A(n_2013),
.Y(n_2185)
);

OAI21x1_ASAP7_75t_L g2186 ( 
.A1(n_2125),
.A2(n_463),
.B(n_462),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_2014),
.Y(n_2187)
);

INVx1_ASAP7_75t_SL g2188 ( 
.A(n_2060),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2070),
.Y(n_2189)
);

OAI21x1_ASAP7_75t_L g2190 ( 
.A1(n_2072),
.A2(n_466),
.B(n_465),
.Y(n_2190)
);

OAI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2133),
.A2(n_1250),
.B1(n_1257),
.B2(n_1252),
.Y(n_2191)
);

OAI21x1_ASAP7_75t_L g2192 ( 
.A1(n_2084),
.A2(n_470),
.B(n_468),
.Y(n_2192)
);

BUFx2_ASAP7_75t_L g2193 ( 
.A(n_2046),
.Y(n_2193)
);

AO32x2_ASAP7_75t_L g2194 ( 
.A1(n_2129),
.A2(n_42),
.A3(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_2015),
.Y(n_2195)
);

OAI21x1_ASAP7_75t_L g2196 ( 
.A1(n_2087),
.A2(n_477),
.B(n_476),
.Y(n_2196)
);

CKINVDCx20_ASAP7_75t_R g2197 ( 
.A(n_2007),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2075),
.Y(n_2198)
);

CKINVDCx12_ASAP7_75t_R g2199 ( 
.A(n_2056),
.Y(n_2199)
);

OAI21x1_ASAP7_75t_L g2200 ( 
.A1(n_2096),
.A2(n_480),
.B(n_478),
.Y(n_2200)
);

CKINVDCx16_ASAP7_75t_R g2201 ( 
.A(n_2067),
.Y(n_2201)
);

OAI21x1_ASAP7_75t_L g2202 ( 
.A1(n_2110),
.A2(n_482),
.B(n_481),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2078),
.Y(n_2203)
);

OAI222xp33_ASAP7_75t_L g2204 ( 
.A1(n_2065),
.A2(n_1265),
.B1(n_1259),
.B2(n_1268),
.C1(n_1261),
.C2(n_1245),
.Y(n_2204)
);

INVx1_ASAP7_75t_SL g2205 ( 
.A(n_2077),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_2008),
.Y(n_2206)
);

AO31x2_ASAP7_75t_L g2207 ( 
.A1(n_2123),
.A2(n_485),
.A3(n_487),
.B(n_483),
.Y(n_2207)
);

NOR2xp33_ASAP7_75t_R g2208 ( 
.A(n_2048),
.B(n_1270),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2082),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2102),
.Y(n_2210)
);

OA21x2_ASAP7_75t_L g2211 ( 
.A1(n_2124),
.A2(n_1275),
.B(n_1271),
.Y(n_2211)
);

OAI21x1_ASAP7_75t_SL g2212 ( 
.A1(n_2130),
.A2(n_41),
.B(n_44),
.Y(n_2212)
);

OAI21x1_ASAP7_75t_L g2213 ( 
.A1(n_2126),
.A2(n_489),
.B(n_488),
.Y(n_2213)
);

OA21x2_ASAP7_75t_L g2214 ( 
.A1(n_2127),
.A2(n_1278),
.B(n_1277),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_L g2215 ( 
.A(n_2091),
.B(n_45),
.Y(n_2215)
);

OAI22xp5_ASAP7_75t_SL g2216 ( 
.A1(n_2069),
.A2(n_1293),
.B1(n_1295),
.B2(n_1289),
.Y(n_2216)
);

OAI21x1_ASAP7_75t_L g2217 ( 
.A1(n_2128),
.A2(n_494),
.B(n_491),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2103),
.Y(n_2218)
);

INVx3_ASAP7_75t_SL g2219 ( 
.A(n_2023),
.Y(n_2219)
);

AOI22xp33_ASAP7_75t_L g2220 ( 
.A1(n_2053),
.A2(n_1311),
.B1(n_1307),
.B2(n_47),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_2013),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2092),
.Y(n_2222)
);

OAI22xp33_ASAP7_75t_L g2223 ( 
.A1(n_2056),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2047),
.B(n_46),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2063),
.B(n_48),
.Y(n_2225)
);

NAND2x1p5_ASAP7_75t_L g2226 ( 
.A(n_2011),
.B(n_495),
.Y(n_2226)
);

OAI21x1_ASAP7_75t_L g2227 ( 
.A1(n_2135),
.A2(n_497),
.B(n_496),
.Y(n_2227)
);

OAI21x1_ASAP7_75t_L g2228 ( 
.A1(n_2071),
.A2(n_499),
.B(n_498),
.Y(n_2228)
);

OAI221xp5_ASAP7_75t_L g2229 ( 
.A1(n_2049),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.C(n_52),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_2041),
.Y(n_2230)
);

INVx2_ASAP7_75t_SL g2231 ( 
.A(n_2032),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2109),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2006),
.B(n_49),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_2073),
.A2(n_501),
.B(n_500),
.Y(n_2234)
);

AO21x2_ASAP7_75t_L g2235 ( 
.A1(n_2064),
.A2(n_506),
.B(n_503),
.Y(n_2235)
);

NAND2x1p5_ASAP7_75t_L g2236 ( 
.A(n_2032),
.B(n_508),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2109),
.Y(n_2237)
);

OAI21x1_ASAP7_75t_L g2238 ( 
.A1(n_2093),
.A2(n_510),
.B(n_509),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2114),
.B(n_50),
.Y(n_2239)
);

NOR2xp67_ASAP7_75t_L g2240 ( 
.A(n_2037),
.B(n_512),
.Y(n_2240)
);

BUFx2_ASAP7_75t_L g2241 ( 
.A(n_2150),
.Y(n_2241)
);

AOI22xp33_ASAP7_75t_L g2242 ( 
.A1(n_2175),
.A2(n_2229),
.B1(n_2036),
.B2(n_2137),
.Y(n_2242)
);

OAI221xp5_ASAP7_75t_L g2243 ( 
.A1(n_2151),
.A2(n_2027),
.B1(n_2081),
.B2(n_2131),
.C(n_2108),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_2220),
.A2(n_2094),
.B1(n_2088),
.B2(n_2117),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2155),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2223),
.A2(n_2141),
.B1(n_2099),
.B2(n_2118),
.Y(n_2246)
);

AOI22xp33_ASAP7_75t_SL g2247 ( 
.A1(n_2212),
.A2(n_2058),
.B1(n_2119),
.B2(n_2050),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2149),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2161),
.B(n_2119),
.Y(n_2249)
);

HB1xp67_ASAP7_75t_L g2250 ( 
.A(n_2195),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2162),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2168),
.Y(n_2252)
);

AOI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_2164),
.A2(n_2092),
.B1(n_2097),
.B2(n_2051),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2174),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2148),
.B(n_2140),
.Y(n_2255)
);

BUFx2_ASAP7_75t_L g2256 ( 
.A(n_2193),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2198),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2188),
.B(n_2090),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2171),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_2172),
.B(n_2003),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_2232),
.Y(n_2261)
);

OAI211xp5_ASAP7_75t_L g2262 ( 
.A1(n_2178),
.A2(n_2104),
.B(n_2083),
.C(n_2134),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2209),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2215),
.A2(n_2035),
.B1(n_2026),
.B2(n_2121),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_2158),
.Y(n_2265)
);

INVx2_ASAP7_75t_SL g2266 ( 
.A(n_2183),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2182),
.B(n_2074),
.Y(n_2267)
);

AOI221xp5_ASAP7_75t_L g2268 ( 
.A1(n_2204),
.A2(n_2076),
.B1(n_2079),
.B2(n_2111),
.C(n_2080),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_SL g2269 ( 
.A1(n_2166),
.A2(n_2086),
.B1(n_2136),
.B2(n_2089),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2189),
.Y(n_2270)
);

INVx1_ASAP7_75t_SL g2271 ( 
.A(n_2205),
.Y(n_2271)
);

A2O1A1Ixp33_ASAP7_75t_L g2272 ( 
.A1(n_2227),
.A2(n_2116),
.B(n_2113),
.C(n_2101),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_2226),
.B(n_2180),
.Y(n_2273)
);

HB1xp67_ASAP7_75t_L g2274 ( 
.A(n_2177),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2224),
.B(n_2020),
.Y(n_2275)
);

BUFx2_ASAP7_75t_L g2276 ( 
.A(n_2237),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2203),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2210),
.Y(n_2278)
);

INVx1_ASAP7_75t_SL g2279 ( 
.A(n_2219),
.Y(n_2279)
);

AOI21xp33_ASAP7_75t_L g2280 ( 
.A1(n_2167),
.A2(n_2061),
.B(n_2035),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2233),
.B(n_2062),
.Y(n_2281)
);

AOI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_2176),
.A2(n_2095),
.B1(n_2057),
.B2(n_2043),
.Y(n_2282)
);

INVx1_ASAP7_75t_SL g2283 ( 
.A(n_2230),
.Y(n_2283)
);

OAI221xp5_ASAP7_75t_L g2284 ( 
.A1(n_2216),
.A2(n_2239),
.B1(n_2225),
.B2(n_2147),
.C(n_2173),
.Y(n_2284)
);

AOI22xp33_ASAP7_75t_L g2285 ( 
.A1(n_2211),
.A2(n_2112),
.B1(n_2098),
.B2(n_2004),
.Y(n_2285)
);

AOI22xp33_ASAP7_75t_L g2286 ( 
.A1(n_2214),
.A2(n_2112),
.B1(n_2033),
.B2(n_2138),
.Y(n_2286)
);

INVx4_ASAP7_75t_L g2287 ( 
.A(n_2187),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_2179),
.Y(n_2288)
);

OAI21xp5_ASAP7_75t_L g2289 ( 
.A1(n_2191),
.A2(n_2025),
.B(n_2028),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2157),
.B(n_2055),
.Y(n_2290)
);

AOI22xp33_ASAP7_75t_L g2291 ( 
.A1(n_2218),
.A2(n_2033),
.B1(n_2010),
.B2(n_53),
.Y(n_2291)
);

A2O1A1Ixp33_ASAP7_75t_L g2292 ( 
.A1(n_2186),
.A2(n_54),
.B(n_51),
.C(n_52),
.Y(n_2292)
);

INVxp67_ASAP7_75t_L g2293 ( 
.A(n_2231),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_2241),
.B(n_2159),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2250),
.B(n_2185),
.Y(n_2295)
);

NOR2x1p5_ASAP7_75t_L g2296 ( 
.A(n_2288),
.B(n_2221),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2274),
.B(n_2255),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2244),
.A2(n_2222),
.B1(n_2165),
.B2(n_2235),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2243),
.A2(n_2154),
.B1(n_2152),
.B2(n_2234),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_2256),
.B(n_2201),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2275),
.B(n_2184),
.Y(n_2301)
);

OR2x2_ASAP7_75t_L g2302 ( 
.A(n_2248),
.B(n_2207),
.Y(n_2302)
);

OR2x6_ASAP7_75t_L g2303 ( 
.A(n_2249),
.B(n_2169),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2276),
.B(n_2194),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2251),
.B(n_54),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_R g2306 ( 
.A(n_2265),
.B(n_2153),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2259),
.B(n_55),
.Y(n_2307)
);

NAND3xp33_ASAP7_75t_SL g2308 ( 
.A(n_2284),
.B(n_2208),
.C(n_2197),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_R g2309 ( 
.A(n_2279),
.B(n_2206),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2277),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2270),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_R g2312 ( 
.A(n_2283),
.B(n_2199),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_2271),
.Y(n_2313)
);

AOI22xp33_ASAP7_75t_L g2314 ( 
.A1(n_2246),
.A2(n_2238),
.B1(n_2181),
.B2(n_2217),
.Y(n_2314)
);

OAI221xp5_ASAP7_75t_SL g2315 ( 
.A1(n_2242),
.A2(n_2262),
.B1(n_2291),
.B2(n_2292),
.C(n_2264),
.Y(n_2315)
);

OAI222xp33_ASAP7_75t_L g2316 ( 
.A1(n_2269),
.A2(n_2194),
.B1(n_2236),
.B2(n_2207),
.C1(n_2146),
.C2(n_2213),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2281),
.B(n_2240),
.Y(n_2317)
);

OAI22xp33_ASAP7_75t_L g2318 ( 
.A1(n_2273),
.A2(n_2170),
.B1(n_2160),
.B2(n_2163),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2261),
.B(n_2228),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_2266),
.Y(n_2320)
);

INVx4_ASAP7_75t_L g2321 ( 
.A(n_2287),
.Y(n_2321)
);

NAND2xp33_ASAP7_75t_SL g2322 ( 
.A(n_2287),
.B(n_55),
.Y(n_2322)
);

NAND4xp25_ASAP7_75t_L g2323 ( 
.A(n_2247),
.B(n_58),
.C(n_56),
.D(n_57),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2272),
.B(n_2156),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2261),
.B(n_56),
.Y(n_2325)
);

HB1xp67_ASAP7_75t_L g2326 ( 
.A(n_2267),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_R g2327 ( 
.A(n_2290),
.B(n_57),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_2293),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2258),
.B(n_2190),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2278),
.Y(n_2330)
);

AND2x2_ASAP7_75t_SL g2331 ( 
.A(n_2285),
.B(n_2192),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2260),
.B(n_58),
.Y(n_2332)
);

OAI21xp5_ASAP7_75t_SL g2333 ( 
.A1(n_2282),
.A2(n_2268),
.B(n_2289),
.Y(n_2333)
);

CKINVDCx5p33_ASAP7_75t_R g2334 ( 
.A(n_2245),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2252),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2254),
.B(n_59),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2257),
.B(n_59),
.Y(n_2337)
);

A2O1A1Ixp33_ASAP7_75t_L g2338 ( 
.A1(n_2280),
.A2(n_2200),
.B(n_2202),
.C(n_2196),
.Y(n_2338)
);

CKINVDCx16_ASAP7_75t_R g2339 ( 
.A(n_2263),
.Y(n_2339)
);

NAND2xp33_ASAP7_75t_R g2340 ( 
.A(n_2253),
.B(n_61),
.Y(n_2340)
);

A2O1A1Ixp33_ASAP7_75t_L g2341 ( 
.A1(n_2286),
.A2(n_2145),
.B(n_2144),
.C(n_62),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2256),
.B(n_60),
.Y(n_2342)
);

OAI22xp5_ASAP7_75t_L g2343 ( 
.A1(n_2242),
.A2(n_63),
.B1(n_60),
.B2(n_61),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2256),
.B(n_63),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_2265),
.Y(n_2345)
);

CKINVDCx16_ASAP7_75t_R g2346 ( 
.A(n_2275),
.Y(n_2346)
);

BUFx2_ASAP7_75t_L g2347 ( 
.A(n_2250),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2277),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_R g2349 ( 
.A(n_2288),
.B(n_64),
.Y(n_2349)
);

NAND3xp33_ASAP7_75t_SL g2350 ( 
.A(n_2284),
.B(n_64),
.C(n_65),
.Y(n_2350)
);

BUFx2_ASAP7_75t_L g2351 ( 
.A(n_2347),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2310),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2330),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2346),
.B(n_65),
.Y(n_2354)
);

BUFx2_ASAP7_75t_L g2355 ( 
.A(n_2300),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_2313),
.Y(n_2356)
);

INVx2_ASAP7_75t_SL g2357 ( 
.A(n_2320),
.Y(n_2357)
);

INVx2_ASAP7_75t_SL g2358 ( 
.A(n_2320),
.Y(n_2358)
);

BUFx2_ASAP7_75t_L g2359 ( 
.A(n_2312),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2297),
.B(n_66),
.Y(n_2360)
);

BUFx2_ASAP7_75t_L g2361 ( 
.A(n_2295),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2311),
.Y(n_2362)
);

INVx2_ASAP7_75t_SL g2363 ( 
.A(n_2301),
.Y(n_2363)
);

OR2x2_ASAP7_75t_L g2364 ( 
.A(n_2326),
.B(n_66),
.Y(n_2364)
);

INVx3_ASAP7_75t_L g2365 ( 
.A(n_2321),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2348),
.Y(n_2366)
);

AND2x4_ASAP7_75t_L g2367 ( 
.A(n_2294),
.B(n_67),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2302),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2339),
.B(n_68),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2304),
.B(n_68),
.Y(n_2370)
);

NOR2x1_ASAP7_75t_L g2371 ( 
.A(n_2325),
.B(n_69),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2335),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2305),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2328),
.B(n_70),
.Y(n_2374)
);

HB1xp67_ASAP7_75t_L g2375 ( 
.A(n_2329),
.Y(n_2375)
);

INVx5_ASAP7_75t_L g2376 ( 
.A(n_2303),
.Y(n_2376)
);

HB1xp67_ASAP7_75t_L g2377 ( 
.A(n_2307),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2317),
.B(n_70),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2334),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2319),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2336),
.Y(n_2381)
);

INVx3_ASAP7_75t_L g2382 ( 
.A(n_2303),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2332),
.B(n_71),
.Y(n_2383)
);

OAI22xp5_ASAP7_75t_L g2384 ( 
.A1(n_2315),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_2384)
);

INVxp67_ASAP7_75t_L g2385 ( 
.A(n_2342),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2344),
.B(n_2309),
.Y(n_2386)
);

NOR2x1_ASAP7_75t_L g2387 ( 
.A(n_2296),
.B(n_2324),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2337),
.Y(n_2388)
);

AOI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2318),
.A2(n_72),
.B(n_74),
.Y(n_2389)
);

AOI22xp33_ASAP7_75t_L g2390 ( 
.A1(n_2350),
.A2(n_78),
.B1(n_74),
.B2(n_76),
.Y(n_2390)
);

HB1xp67_ASAP7_75t_L g2391 ( 
.A(n_2331),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2343),
.Y(n_2392)
);

INVx3_ASAP7_75t_L g2393 ( 
.A(n_2345),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2316),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2338),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2333),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2327),
.B(n_76),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2340),
.Y(n_2398)
);

INVxp67_ASAP7_75t_L g2399 ( 
.A(n_2308),
.Y(n_2399)
);

BUFx3_ASAP7_75t_L g2400 ( 
.A(n_2306),
.Y(n_2400)
);

INVxp67_ASAP7_75t_SL g2401 ( 
.A(n_2298),
.Y(n_2401)
);

INVx3_ASAP7_75t_L g2402 ( 
.A(n_2322),
.Y(n_2402)
);

AOI21xp5_ASAP7_75t_SL g2403 ( 
.A1(n_2341),
.A2(n_80),
.B(n_79),
.Y(n_2403)
);

HB1xp67_ASAP7_75t_L g2404 ( 
.A(n_2323),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2314),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2349),
.B(n_78),
.Y(n_2406)
);

NAND3xp33_ASAP7_75t_L g2407 ( 
.A(n_2299),
.B(n_80),
.C(n_81),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2297),
.B(n_81),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2311),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2310),
.Y(n_2410)
);

AOI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2324),
.A2(n_82),
.B(n_83),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2311),
.Y(n_2412)
);

BUFx3_ASAP7_75t_L g2413 ( 
.A(n_2313),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2310),
.Y(n_2414)
);

BUFx2_ASAP7_75t_L g2415 ( 
.A(n_2347),
.Y(n_2415)
);

INVx5_ASAP7_75t_SL g2416 ( 
.A(n_2303),
.Y(n_2416)
);

INVxp67_ASAP7_75t_SL g2417 ( 
.A(n_2297),
.Y(n_2417)
);

HB1xp67_ASAP7_75t_L g2418 ( 
.A(n_2347),
.Y(n_2418)
);

AOI22xp33_ASAP7_75t_L g2419 ( 
.A1(n_2350),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2347),
.B(n_84),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2311),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2347),
.B(n_85),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2310),
.Y(n_2423)
);

BUFx2_ASAP7_75t_L g2424 ( 
.A(n_2347),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2310),
.Y(n_2425)
);

INVxp67_ASAP7_75t_L g2426 ( 
.A(n_2347),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2310),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2311),
.Y(n_2428)
);

NOR2x1_ASAP7_75t_L g2429 ( 
.A(n_2300),
.B(n_86),
.Y(n_2429)
);

BUFx6f_ASAP7_75t_L g2430 ( 
.A(n_2320),
.Y(n_2430)
);

AOI21xp5_ASAP7_75t_SL g2431 ( 
.A1(n_2395),
.A2(n_95),
.B(n_87),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2355),
.B(n_87),
.Y(n_2432)
);

AOI22xp33_ASAP7_75t_L g2433 ( 
.A1(n_2394),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2351),
.B(n_89),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2400),
.B(n_90),
.Y(n_2435)
);

OA21x2_ASAP7_75t_L g2436 ( 
.A1(n_2401),
.A2(n_91),
.B(n_92),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2417),
.B(n_91),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_SL g2438 ( 
.A(n_2387),
.B(n_2376),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2377),
.B(n_2373),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2405),
.B(n_92),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2381),
.B(n_2351),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2415),
.B(n_93),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2424),
.B(n_94),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2418),
.B(n_94),
.Y(n_2444)
);

OAI21xp33_ASAP7_75t_L g2445 ( 
.A1(n_2384),
.A2(n_95),
.B(n_96),
.Y(n_2445)
);

AND2x2_ASAP7_75t_SL g2446 ( 
.A(n_2359),
.B(n_97),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2361),
.B(n_2375),
.Y(n_2447)
);

OAI22xp5_ASAP7_75t_L g2448 ( 
.A1(n_2404),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_2448)
);

INVxp67_ASAP7_75t_SL g2449 ( 
.A(n_2391),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2363),
.B(n_99),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2426),
.B(n_100),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2385),
.B(n_101),
.Y(n_2452)
);

AOI22xp33_ASAP7_75t_L g2453 ( 
.A1(n_2396),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_2453)
);

OAI22xp5_ASAP7_75t_L g2454 ( 
.A1(n_2392),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2380),
.B(n_105),
.Y(n_2455)
);

AOI22xp33_ASAP7_75t_SL g2456 ( 
.A1(n_2398),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2362),
.B(n_106),
.Y(n_2457)
);

NAND3xp33_ASAP7_75t_L g2458 ( 
.A(n_2389),
.B(n_108),
.C(n_109),
.Y(n_2458)
);

OAI221xp5_ASAP7_75t_SL g2459 ( 
.A1(n_2390),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.C(n_113),
.Y(n_2459)
);

NAND4xp25_ASAP7_75t_L g2460 ( 
.A(n_2419),
.B(n_114),
.C(n_111),
.D(n_112),
.Y(n_2460)
);

OAI221xp5_ASAP7_75t_SL g2461 ( 
.A1(n_2403),
.A2(n_117),
.B1(n_114),
.B2(n_115),
.C(n_118),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2409),
.B(n_115),
.Y(n_2462)
);

OAI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2429),
.A2(n_117),
.B(n_118),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2386),
.B(n_119),
.Y(n_2464)
);

OAI22xp5_ASAP7_75t_L g2465 ( 
.A1(n_2402),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_2465)
);

OAI22xp5_ASAP7_75t_L g2466 ( 
.A1(n_2407),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2376),
.B(n_123),
.Y(n_2467)
);

OAI22xp33_ASAP7_75t_L g2468 ( 
.A1(n_2376),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_2468)
);

OAI22xp5_ASAP7_75t_L g2469 ( 
.A1(n_2399),
.A2(n_128),
.B1(n_124),
.B2(n_126),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2354),
.B(n_126),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2357),
.B(n_129),
.Y(n_2471)
);

OAI221xp5_ASAP7_75t_L g2472 ( 
.A1(n_2411),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.C(n_133),
.Y(n_2472)
);

NAND3xp33_ASAP7_75t_L g2473 ( 
.A(n_2371),
.B(n_130),
.C(n_131),
.Y(n_2473)
);

AOI211xp5_ASAP7_75t_L g2474 ( 
.A1(n_2397),
.A2(n_141),
.B(n_149),
.C(n_133),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2358),
.B(n_134),
.Y(n_2475)
);

NOR2xp33_ASAP7_75t_SL g2476 ( 
.A(n_2356),
.B(n_134),
.Y(n_2476)
);

NAND4xp25_ASAP7_75t_SL g2477 ( 
.A(n_2374),
.B(n_137),
.C(n_135),
.D(n_136),
.Y(n_2477)
);

OAI221xp5_ASAP7_75t_L g2478 ( 
.A1(n_2388),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.C(n_138),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2412),
.B(n_138),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2421),
.B(n_2428),
.Y(n_2480)
);

AOI22xp33_ASAP7_75t_L g2481 ( 
.A1(n_2370),
.A2(n_142),
.B1(n_139),
.B2(n_140),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2430),
.B(n_142),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2368),
.B(n_143),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2408),
.B(n_143),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2430),
.B(n_144),
.Y(n_2485)
);

NAND3xp33_ASAP7_75t_L g2486 ( 
.A(n_2364),
.B(n_145),
.C(n_146),
.Y(n_2486)
);

NAND2x1_ASAP7_75t_L g2487 ( 
.A(n_2365),
.B(n_2382),
.Y(n_2487)
);

NAND3xp33_ASAP7_75t_L g2488 ( 
.A(n_2383),
.B(n_146),
.C(n_147),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2360),
.B(n_2420),
.Y(n_2489)
);

AOI221xp5_ASAP7_75t_L g2490 ( 
.A1(n_2369),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.C(n_150),
.Y(n_2490)
);

OAI21xp5_ASAP7_75t_SL g2491 ( 
.A1(n_2406),
.A2(n_2422),
.B(n_2367),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2378),
.B(n_150),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2413),
.B(n_151),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2372),
.B(n_151),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2366),
.B(n_152),
.Y(n_2495)
);

AOI22xp5_ASAP7_75t_L g2496 ( 
.A1(n_2379),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2416),
.B(n_154),
.Y(n_2497)
);

OAI21xp5_ASAP7_75t_SL g2498 ( 
.A1(n_2393),
.A2(n_155),
.B(n_157),
.Y(n_2498)
);

AOI22xp33_ASAP7_75t_SL g2499 ( 
.A1(n_2416),
.A2(n_159),
.B1(n_155),
.B2(n_158),
.Y(n_2499)
);

NAND3xp33_ASAP7_75t_L g2500 ( 
.A(n_2352),
.B(n_158),
.C(n_161),
.Y(n_2500)
);

OAI22xp5_ASAP7_75t_L g2501 ( 
.A1(n_2353),
.A2(n_165),
.B1(n_162),
.B2(n_164),
.Y(n_2501)
);

OAI21xp5_ASAP7_75t_L g2502 ( 
.A1(n_2410),
.A2(n_165),
.B(n_166),
.Y(n_2502)
);

NAND4xp25_ASAP7_75t_L g2503 ( 
.A(n_2414),
.B(n_168),
.C(n_166),
.D(n_167),
.Y(n_2503)
);

NAND3xp33_ASAP7_75t_L g2504 ( 
.A(n_2423),
.B(n_167),
.C(n_170),
.Y(n_2504)
);

NOR3xp33_ASAP7_75t_SL g2505 ( 
.A(n_2425),
.B(n_170),
.C(n_171),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_SL g2506 ( 
.A(n_2427),
.B(n_171),
.Y(n_2506)
);

NAND3xp33_ASAP7_75t_L g2507 ( 
.A(n_2395),
.B(n_173),
.C(n_174),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2355),
.B(n_173),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2355),
.B(n_174),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2417),
.B(n_177),
.Y(n_2510)
);

OR2x2_ASAP7_75t_L g2511 ( 
.A(n_2417),
.B(n_177),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2417),
.B(n_178),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2417),
.B(n_178),
.Y(n_2513)
);

NOR2xp33_ASAP7_75t_L g2514 ( 
.A(n_2400),
.B(n_179),
.Y(n_2514)
);

NAND3xp33_ASAP7_75t_L g2515 ( 
.A(n_2395),
.B(n_179),
.C(n_180),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2417),
.B(n_180),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2355),
.B(n_181),
.Y(n_2517)
);

AND2x2_ASAP7_75t_SL g2518 ( 
.A(n_2359),
.B(n_182),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2355),
.B(n_182),
.Y(n_2519)
);

NAND3xp33_ASAP7_75t_L g2520 ( 
.A(n_2395),
.B(n_183),
.C(n_184),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2417),
.B(n_183),
.Y(n_2521)
);

OAI221xp5_ASAP7_75t_SL g2522 ( 
.A1(n_2396),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.C(n_187),
.Y(n_2522)
);

OAI21xp33_ASAP7_75t_L g2523 ( 
.A1(n_2395),
.A2(n_186),
.B(n_188),
.Y(n_2523)
);

NOR3xp33_ASAP7_75t_L g2524 ( 
.A(n_2384),
.B(n_188),
.C(n_189),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2417),
.B(n_189),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2417),
.B(n_190),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2355),
.B(n_192),
.Y(n_2527)
);

NAND4xp25_ASAP7_75t_L g2528 ( 
.A(n_2384),
.B(n_194),
.C(n_192),
.D(n_193),
.Y(n_2528)
);

AND2x2_ASAP7_75t_SL g2529 ( 
.A(n_2359),
.B(n_193),
.Y(n_2529)
);

OA21x2_ASAP7_75t_L g2530 ( 
.A1(n_2394),
.A2(n_194),
.B(n_196),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2368),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2355),
.B(n_196),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2417),
.B(n_198),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2355),
.B(n_199),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2417),
.B(n_199),
.Y(n_2535)
);

OAI21xp5_ASAP7_75t_SL g2536 ( 
.A1(n_2384),
.A2(n_200),
.B(n_201),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2417),
.B(n_201),
.Y(n_2537)
);

AOI21xp33_ASAP7_75t_SL g2538 ( 
.A1(n_2386),
.A2(n_203),
.B(n_204),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_2355),
.B(n_203),
.Y(n_2539)
);

OAI21xp5_ASAP7_75t_L g2540 ( 
.A1(n_2396),
.A2(n_204),
.B(n_205),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2417),
.B(n_205),
.Y(n_2541)
);

OAI221xp5_ASAP7_75t_SL g2542 ( 
.A1(n_2396),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.C(n_210),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2355),
.B(n_207),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_SL g2544 ( 
.A(n_2387),
.B(n_208),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2355),
.B(n_209),
.Y(n_2545)
);

INVxp67_ASAP7_75t_L g2546 ( 
.A(n_2441),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2480),
.Y(n_2547)
);

NAND2x1p5_ASAP7_75t_L g2548 ( 
.A(n_2438),
.B(n_211),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2447),
.B(n_212),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2531),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2530),
.Y(n_2551)
);

OR2x2_ASAP7_75t_L g2552 ( 
.A(n_2439),
.B(n_212),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2530),
.Y(n_2553)
);

INVxp67_ASAP7_75t_L g2554 ( 
.A(n_2440),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2449),
.B(n_213),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2437),
.B(n_213),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2495),
.Y(n_2557)
);

INVxp67_ASAP7_75t_L g2558 ( 
.A(n_2544),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2494),
.Y(n_2559)
);

HB1xp67_ASAP7_75t_L g2560 ( 
.A(n_2434),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2510),
.B(n_214),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2457),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2462),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2487),
.B(n_214),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2489),
.B(n_215),
.Y(n_2565)
);

AND2x4_ASAP7_75t_L g2566 ( 
.A(n_2455),
.B(n_2450),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2512),
.B(n_215),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2436),
.Y(n_2568)
);

HB1xp67_ASAP7_75t_L g2569 ( 
.A(n_2513),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2483),
.Y(n_2570)
);

HB1xp67_ASAP7_75t_L g2571 ( 
.A(n_2516),
.Y(n_2571)
);

OR2x2_ASAP7_75t_L g2572 ( 
.A(n_2511),
.B(n_216),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2521),
.Y(n_2573)
);

BUFx2_ASAP7_75t_L g2574 ( 
.A(n_2432),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2525),
.B(n_2526),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2508),
.B(n_217),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2509),
.B(n_217),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2533),
.B(n_218),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2517),
.B(n_218),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2519),
.B(n_219),
.Y(n_2580)
);

OR2x2_ASAP7_75t_L g2581 ( 
.A(n_2535),
.B(n_220),
.Y(n_2581)
);

NAND3xp33_ASAP7_75t_L g2582 ( 
.A(n_2474),
.B(n_220),
.C(n_221),
.Y(n_2582)
);

NAND3xp33_ASAP7_75t_L g2583 ( 
.A(n_2524),
.B(n_223),
.C(n_224),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2527),
.B(n_224),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2532),
.B(n_225),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2537),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2541),
.B(n_226),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2444),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2534),
.B(n_226),
.Y(n_2589)
);

INVx1_ASAP7_75t_SL g2590 ( 
.A(n_2446),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2539),
.B(n_227),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2479),
.Y(n_2592)
);

INVx2_ASAP7_75t_SL g2593 ( 
.A(n_2543),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2436),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2545),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2442),
.B(n_2443),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2451),
.B(n_227),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2452),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2506),
.Y(n_2599)
);

BUFx2_ASAP7_75t_L g2600 ( 
.A(n_2464),
.Y(n_2600)
);

NAND3xp33_ASAP7_75t_L g2601 ( 
.A(n_2536),
.B(n_228),
.C(n_229),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2484),
.B(n_228),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2491),
.B(n_229),
.Y(n_2603)
);

CKINVDCx16_ASAP7_75t_R g2604 ( 
.A(n_2476),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2493),
.B(n_230),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2470),
.B(n_230),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2471),
.B(n_2475),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2482),
.Y(n_2608)
);

HB1xp67_ASAP7_75t_L g2609 ( 
.A(n_2492),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2486),
.B(n_231),
.Y(n_2610)
);

AND2x4_ASAP7_75t_L g2611 ( 
.A(n_2485),
.B(n_231),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2488),
.B(n_232),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2518),
.B(n_233),
.Y(n_2613)
);

OR2x2_ASAP7_75t_L g2614 ( 
.A(n_2497),
.B(n_233),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2500),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2504),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2473),
.Y(n_2617)
);

NOR2xp67_ASAP7_75t_L g2618 ( 
.A(n_2538),
.B(n_234),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2529),
.B(n_234),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2498),
.B(n_235),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2507),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2523),
.B(n_235),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2515),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2520),
.B(n_236),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2467),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2435),
.B(n_237),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2431),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2454),
.Y(n_2628)
);

INVx4_ASAP7_75t_L g2629 ( 
.A(n_2514),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2463),
.B(n_237),
.Y(n_2630)
);

OR2x2_ASAP7_75t_L g2631 ( 
.A(n_2503),
.B(n_2477),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2481),
.B(n_238),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2465),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2496),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2502),
.B(n_238),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2505),
.B(n_239),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2540),
.B(n_239),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2490),
.B(n_240),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2501),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2478),
.Y(n_2640)
);

AND2x4_ASAP7_75t_L g2641 ( 
.A(n_2458),
.B(n_241),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2448),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2469),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2468),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2456),
.B(n_241),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2445),
.B(n_242),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2499),
.B(n_242),
.Y(n_2647)
);

OR2x2_ASAP7_75t_L g2648 ( 
.A(n_2528),
.B(n_243),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2472),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2466),
.B(n_243),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2460),
.B(n_244),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2433),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2522),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2542),
.Y(n_2654)
);

AND2x4_ASAP7_75t_L g2655 ( 
.A(n_2453),
.B(n_245),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2461),
.B(n_245),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2459),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2439),
.B(n_246),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2439),
.B(n_246),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2531),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2480),
.Y(n_2661)
);

OR2x2_ASAP7_75t_L g2662 ( 
.A(n_2439),
.B(n_248),
.Y(n_2662)
);

OR2x2_ASAP7_75t_L g2663 ( 
.A(n_2439),
.B(n_248),
.Y(n_2663)
);

OAI21xp33_ASAP7_75t_L g2664 ( 
.A1(n_2536),
.A2(n_249),
.B(n_250),
.Y(n_2664)
);

AND2x2_ASAP7_75t_L g2665 ( 
.A(n_2447),
.B(n_249),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2447),
.B(n_250),
.Y(n_2666)
);

AND2x4_ASAP7_75t_L g2667 ( 
.A(n_2447),
.B(n_251),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2531),
.Y(n_2668)
);

INVxp67_ASAP7_75t_L g2669 ( 
.A(n_2441),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2447),
.B(n_251),
.Y(n_2670)
);

INVx1_ASAP7_75t_SL g2671 ( 
.A(n_2446),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2447),
.B(n_252),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2480),
.Y(n_2673)
);

OR2x2_ASAP7_75t_L g2674 ( 
.A(n_2439),
.B(n_252),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2447),
.B(n_253),
.Y(n_2675)
);

OR2x2_ASAP7_75t_L g2676 ( 
.A(n_2439),
.B(n_253),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2480),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2447),
.B(n_254),
.Y(n_2678)
);

AND2x4_ASAP7_75t_L g2679 ( 
.A(n_2447),
.B(n_255),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2480),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2480),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2480),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2439),
.B(n_255),
.Y(n_2683)
);

BUFx2_ASAP7_75t_L g2684 ( 
.A(n_2574),
.Y(n_2684)
);

HB1xp67_ASAP7_75t_L g2685 ( 
.A(n_2569),
.Y(n_2685)
);

OR2x2_ASAP7_75t_L g2686 ( 
.A(n_2574),
.B(n_256),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2593),
.B(n_256),
.Y(n_2687)
);

INVxp67_ASAP7_75t_L g2688 ( 
.A(n_2627),
.Y(n_2688)
);

BUFx3_ASAP7_75t_L g2689 ( 
.A(n_2611),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2571),
.B(n_257),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2550),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2600),
.B(n_257),
.Y(n_2692)
);

AND2x4_ASAP7_75t_L g2693 ( 
.A(n_2566),
.B(n_258),
.Y(n_2693)
);

INVx2_ASAP7_75t_SL g2694 ( 
.A(n_2607),
.Y(n_2694)
);

OR2x2_ASAP7_75t_L g2695 ( 
.A(n_2547),
.B(n_259),
.Y(n_2695)
);

OR2x2_ASAP7_75t_L g2696 ( 
.A(n_2661),
.B(n_260),
.Y(n_2696)
);

INVxp67_ASAP7_75t_SL g2697 ( 
.A(n_2560),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2551),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2673),
.Y(n_2699)
);

OR2x2_ASAP7_75t_L g2700 ( 
.A(n_2677),
.B(n_260),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2680),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2681),
.B(n_261),
.Y(n_2702)
);

OR2x2_ASAP7_75t_L g2703 ( 
.A(n_2682),
.B(n_261),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2660),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2596),
.B(n_262),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_2546),
.B(n_263),
.Y(n_2706)
);

INVx1_ASAP7_75t_SL g2707 ( 
.A(n_2590),
.Y(n_2707)
);

AND2x4_ASAP7_75t_L g2708 ( 
.A(n_2595),
.B(n_264),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2573),
.B(n_264),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2668),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2594),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2559),
.Y(n_2712)
);

NOR2xp67_ASAP7_75t_L g2713 ( 
.A(n_2629),
.B(n_265),
.Y(n_2713)
);

AND2x4_ASAP7_75t_L g2714 ( 
.A(n_2608),
.B(n_266),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2553),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2586),
.B(n_266),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2568),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2562),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2625),
.Y(n_2719)
);

OR2x2_ASAP7_75t_L g2720 ( 
.A(n_2669),
.B(n_267),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2609),
.B(n_267),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2588),
.B(n_268),
.Y(n_2722)
);

INVx2_ASAP7_75t_SL g2723 ( 
.A(n_2667),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2563),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2549),
.B(n_268),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2554),
.B(n_269),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2557),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2665),
.B(n_269),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2570),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2599),
.Y(n_2730)
);

OR2x2_ASAP7_75t_L g2731 ( 
.A(n_2575),
.B(n_270),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2564),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2666),
.B(n_270),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2644),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2639),
.Y(n_2735)
);

OR2x2_ASAP7_75t_L g2736 ( 
.A(n_2592),
.B(n_2552),
.Y(n_2736)
);

INVxp67_ASAP7_75t_L g2737 ( 
.A(n_2657),
.Y(n_2737)
);

AND2x4_ASAP7_75t_L g2738 ( 
.A(n_2679),
.B(n_271),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2670),
.B(n_271),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2617),
.Y(n_2740)
);

INVxp33_ASAP7_75t_L g2741 ( 
.A(n_2618),
.Y(n_2741)
);

OR2x2_ASAP7_75t_L g2742 ( 
.A(n_2662),
.B(n_2663),
.Y(n_2742)
);

NOR2x1_ASAP7_75t_L g2743 ( 
.A(n_2603),
.B(n_272),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2598),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2548),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2615),
.B(n_272),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2616),
.B(n_274),
.Y(n_2747)
);

OR2x2_ASAP7_75t_L g2748 ( 
.A(n_2674),
.B(n_274),
.Y(n_2748)
);

NAND4xp25_ASAP7_75t_L g2749 ( 
.A(n_2601),
.B(n_278),
.C(n_275),
.D(n_276),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2628),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2658),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2659),
.Y(n_2752)
);

BUFx2_ASAP7_75t_L g2753 ( 
.A(n_2621),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2683),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2555),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2676),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2623),
.Y(n_2757)
);

INVxp67_ASAP7_75t_SL g2758 ( 
.A(n_2558),
.Y(n_2758)
);

AOI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2664),
.A2(n_278),
.B1(n_275),
.B2(n_276),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2643),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2633),
.Y(n_2761)
);

OR2x2_ASAP7_75t_L g2762 ( 
.A(n_2642),
.B(n_2634),
.Y(n_2762)
);

AND2x6_ASAP7_75t_SL g2763 ( 
.A(n_2606),
.B(n_279),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2672),
.B(n_279),
.Y(n_2764)
);

INVx1_ASAP7_75t_SL g2765 ( 
.A(n_2671),
.Y(n_2765)
);

OR2x2_ASAP7_75t_L g2766 ( 
.A(n_2572),
.B(n_280),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2675),
.B(n_2678),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2614),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2565),
.B(n_280),
.Y(n_2769)
);

OR2x2_ASAP7_75t_L g2770 ( 
.A(n_2649),
.B(n_281),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2576),
.B(n_281),
.Y(n_2771)
);

OR2x2_ASAP7_75t_L g2772 ( 
.A(n_2578),
.B(n_282),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2653),
.B(n_2640),
.Y(n_2773)
);

OR2x2_ASAP7_75t_L g2774 ( 
.A(n_2581),
.B(n_282),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2654),
.B(n_283),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2597),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2577),
.B(n_283),
.Y(n_2777)
);

NOR2xp67_ASAP7_75t_L g2778 ( 
.A(n_2619),
.B(n_284),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2579),
.B(n_284),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2652),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2556),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2605),
.Y(n_2782)
);

OR2x2_ASAP7_75t_L g2783 ( 
.A(n_2561),
.B(n_285),
.Y(n_2783)
);

NOR2xp67_ASAP7_75t_R g2784 ( 
.A(n_2604),
.B(n_285),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2567),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2587),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2580),
.B(n_286),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2610),
.Y(n_2788)
);

OR2x2_ASAP7_75t_L g2789 ( 
.A(n_2602),
.B(n_286),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2584),
.B(n_2585),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_2631),
.B(n_287),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2612),
.Y(n_2792)
);

OR2x2_ASAP7_75t_L g2793 ( 
.A(n_2648),
.B(n_287),
.Y(n_2793)
);

NOR2x1_ASAP7_75t_L g2794 ( 
.A(n_2589),
.B(n_288),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2641),
.B(n_288),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2591),
.B(n_289),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2624),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2646),
.Y(n_2798)
);

OR2x2_ASAP7_75t_L g2799 ( 
.A(n_2656),
.B(n_289),
.Y(n_2799)
);

INVx2_ASAP7_75t_SL g2800 ( 
.A(n_2626),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2636),
.B(n_290),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2613),
.B(n_290),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2622),
.Y(n_2803)
);

OR2x2_ASAP7_75t_L g2804 ( 
.A(n_2651),
.B(n_291),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2620),
.B(n_292),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2637),
.B(n_292),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2630),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2635),
.Y(n_2808)
);

OR2x2_ASAP7_75t_L g2809 ( 
.A(n_2650),
.B(n_293),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2647),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2638),
.B(n_2583),
.Y(n_2811)
);

AND2x4_ASAP7_75t_L g2812 ( 
.A(n_2582),
.B(n_293),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2645),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2655),
.B(n_294),
.Y(n_2814)
);

AND2x2_ASAP7_75t_L g2815 ( 
.A(n_2632),
.B(n_294),
.Y(n_2815)
);

NOR2x1p5_ASAP7_75t_L g2816 ( 
.A(n_2631),
.B(n_295),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2550),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2574),
.B(n_296),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2629),
.B(n_296),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2550),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2550),
.Y(n_2821)
);

OR2x2_ASAP7_75t_L g2822 ( 
.A(n_2574),
.B(n_297),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2574),
.B(n_298),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2550),
.Y(n_2824)
);

OR2x2_ASAP7_75t_L g2825 ( 
.A(n_2574),
.B(n_299),
.Y(n_2825)
);

OR2x2_ASAP7_75t_L g2826 ( 
.A(n_2574),
.B(n_301),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2550),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2550),
.Y(n_2828)
);

OR2x2_ASAP7_75t_L g2829 ( 
.A(n_2574),
.B(n_301),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2574),
.B(n_302),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2574),
.B(n_303),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2569),
.B(n_303),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2574),
.B(n_304),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2574),
.B(n_304),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2574),
.B(n_305),
.Y(n_2835)
);

NAND2x1p5_ASAP7_75t_L g2836 ( 
.A(n_2667),
.B(n_305),
.Y(n_2836)
);

OAI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2631),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2574),
.B(n_306),
.Y(n_2838)
);

HB1xp67_ASAP7_75t_L g2839 ( 
.A(n_2569),
.Y(n_2839)
);

AND2x2_ASAP7_75t_L g2840 ( 
.A(n_2574),
.B(n_307),
.Y(n_2840)
);

OR2x2_ASAP7_75t_L g2841 ( 
.A(n_2574),
.B(n_308),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2574),
.B(n_309),
.Y(n_2842)
);

BUFx2_ASAP7_75t_L g2843 ( 
.A(n_2574),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2550),
.Y(n_2844)
);

AND2x4_ASAP7_75t_L g2845 ( 
.A(n_2574),
.B(n_309),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2550),
.Y(n_2846)
);

INVx2_ASAP7_75t_SL g2847 ( 
.A(n_2607),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2569),
.B(n_310),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2574),
.B(n_310),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2574),
.B(n_311),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2574),
.B(n_311),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2550),
.Y(n_2852)
);

NAND2x1p5_ASAP7_75t_L g2853 ( 
.A(n_2667),
.B(n_312),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2574),
.B(n_312),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_L g2855 ( 
.A(n_2629),
.B(n_313),
.Y(n_2855)
);

INVx3_ASAP7_75t_L g2856 ( 
.A(n_2566),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2574),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2574),
.B(n_314),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2574),
.B(n_314),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2550),
.Y(n_2860)
);

OR2x2_ASAP7_75t_L g2861 ( 
.A(n_2574),
.B(n_316),
.Y(n_2861)
);

AND2x2_ASAP7_75t_L g2862 ( 
.A(n_2574),
.B(n_316),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2574),
.B(n_317),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2550),
.Y(n_2864)
);

INVx3_ASAP7_75t_L g2865 ( 
.A(n_2566),
.Y(n_2865)
);

OR2x2_ASAP7_75t_L g2866 ( 
.A(n_2574),
.B(n_317),
.Y(n_2866)
);

AND2x4_ASAP7_75t_L g2867 ( 
.A(n_2574),
.B(n_318),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2550),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_2574),
.B(n_318),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2550),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2574),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2569),
.B(n_319),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2569),
.B(n_319),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2569),
.B(n_320),
.Y(n_2874)
);

BUFx2_ASAP7_75t_L g2875 ( 
.A(n_2574),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2550),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2685),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2839),
.Y(n_2878)
);

HB1xp67_ASAP7_75t_L g2879 ( 
.A(n_2707),
.Y(n_2879)
);

INVxp67_ASAP7_75t_L g2880 ( 
.A(n_2784),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2711),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2684),
.B(n_320),
.Y(n_2882)
);

HB1xp67_ASAP7_75t_L g2883 ( 
.A(n_2765),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2735),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2750),
.Y(n_2885)
);

OAI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2758),
.A2(n_324),
.B1(n_321),
.B2(n_322),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2800),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2691),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2813),
.A2(n_325),
.B1(n_322),
.B2(n_324),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2817),
.Y(n_2890)
);

INVx1_ASAP7_75t_SL g2891 ( 
.A(n_2790),
.Y(n_2891)
);

OAI222xp33_ASAP7_75t_L g2892 ( 
.A1(n_2688),
.A2(n_2803),
.B1(n_2780),
.B2(n_2798),
.C1(n_2743),
.C2(n_2753),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2684),
.B(n_2737),
.Y(n_2893)
);

AOI22xp33_ASAP7_75t_L g2894 ( 
.A1(n_2698),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_2894)
);

AND2x2_ASAP7_75t_L g2895 ( 
.A(n_2856),
.B(n_327),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2820),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2821),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2824),
.Y(n_2898)
);

O2A1O1Ixp5_ASAP7_75t_R g2899 ( 
.A1(n_2811),
.A2(n_331),
.B(n_329),
.C(n_330),
.Y(n_2899)
);

BUFx2_ASAP7_75t_L g2900 ( 
.A(n_2843),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2827),
.Y(n_2901)
);

OAI322xp33_ASAP7_75t_L g2902 ( 
.A1(n_2757),
.A2(n_336),
.A3(n_335),
.B1(n_333),
.B2(n_329),
.C1(n_332),
.C2(n_334),
.Y(n_2902)
);

OAI322xp33_ASAP7_75t_L g2903 ( 
.A1(n_2740),
.A2(n_340),
.A3(n_339),
.B1(n_337),
.B2(n_332),
.C1(n_334),
.C2(n_338),
.Y(n_2903)
);

OR3x2_ASAP7_75t_L g2904 ( 
.A(n_2749),
.B(n_2822),
.C(n_2686),
.Y(n_2904)
);

OR2x2_ASAP7_75t_L g2905 ( 
.A(n_2760),
.B(n_339),
.Y(n_2905)
);

AOI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2812),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.Y(n_2906)
);

OAI22xp33_ASAP7_75t_SL g2907 ( 
.A1(n_2825),
.A2(n_345),
.B1(n_342),
.B2(n_344),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2828),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2844),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2846),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2852),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2860),
.Y(n_2912)
);

INVxp67_ASAP7_75t_SL g2913 ( 
.A(n_2816),
.Y(n_2913)
);

NOR4xp25_ASAP7_75t_L g2914 ( 
.A(n_2797),
.B(n_348),
.C(n_345),
.D(n_346),
.Y(n_2914)
);

AOI32xp33_ASAP7_75t_L g2915 ( 
.A1(n_2741),
.A2(n_349),
.A3(n_351),
.B1(n_348),
.B2(n_350),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2782),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2818),
.B(n_346),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2823),
.B(n_350),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2865),
.Y(n_2919)
);

INVx1_ASAP7_75t_SL g2920 ( 
.A(n_2689),
.Y(n_2920)
);

OA222x2_ASAP7_75t_L g2921 ( 
.A1(n_2826),
.A2(n_353),
.B1(n_355),
.B2(n_351),
.C1(n_352),
.C2(n_354),
.Y(n_2921)
);

OA222x2_ASAP7_75t_L g2922 ( 
.A1(n_2829),
.A2(n_356),
.B1(n_358),
.B2(n_352),
.C1(n_355),
.C2(n_357),
.Y(n_2922)
);

AND3x1_ASAP7_75t_SL g2923 ( 
.A(n_2755),
.B(n_356),
.C(n_357),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2830),
.B(n_359),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2694),
.B(n_359),
.Y(n_2925)
);

BUFx3_ASAP7_75t_L g2926 ( 
.A(n_2738),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2864),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2831),
.B(n_360),
.Y(n_2928)
);

INVx2_ASAP7_75t_SL g2929 ( 
.A(n_2845),
.Y(n_2929)
);

NAND3xp33_ASAP7_75t_L g2930 ( 
.A(n_2759),
.B(n_360),
.C(n_362),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2868),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2870),
.Y(n_2932)
);

NAND4xp75_ASAP7_75t_L g2933 ( 
.A(n_2794),
.B(n_364),
.C(n_362),
.D(n_363),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2876),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2718),
.Y(n_2935)
);

NAND3xp33_ASAP7_75t_L g2936 ( 
.A(n_2875),
.B(n_363),
.C(n_364),
.Y(n_2936)
);

AOI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2778),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2724),
.Y(n_2938)
);

AND2x2_ASAP7_75t_L g2939 ( 
.A(n_2847),
.B(n_2767),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2727),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2729),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2833),
.B(n_367),
.Y(n_2942)
);

AOI322xp5_ASAP7_75t_L g2943 ( 
.A1(n_2810),
.A2(n_374),
.A3(n_373),
.B1(n_370),
.B2(n_368),
.C1(n_369),
.C2(n_372),
.Y(n_2943)
);

OR2x2_ASAP7_75t_L g2944 ( 
.A(n_2744),
.B(n_369),
.Y(n_2944)
);

AOI32xp33_ASAP7_75t_L g2945 ( 
.A1(n_2806),
.A2(n_373),
.A3(n_375),
.B1(n_372),
.B2(n_374),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2834),
.B(n_370),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2776),
.Y(n_2947)
);

HB1xp67_ASAP7_75t_L g2948 ( 
.A(n_2857),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2712),
.Y(n_2949)
);

AOI22xp5_ASAP7_75t_L g2950 ( 
.A1(n_2788),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2732),
.Y(n_2951)
);

AOI22xp5_ASAP7_75t_L g2952 ( 
.A1(n_2792),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_2952)
);

BUFx2_ASAP7_75t_L g2953 ( 
.A(n_2697),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2699),
.Y(n_2954)
);

A2O1A1Ixp33_ASAP7_75t_L g2955 ( 
.A1(n_2791),
.A2(n_381),
.B(n_379),
.C(n_380),
.Y(n_2955)
);

NOR2xp67_ASAP7_75t_L g2956 ( 
.A(n_2871),
.B(n_380),
.Y(n_2956)
);

AOI22xp5_ASAP7_75t_L g2957 ( 
.A1(n_2768),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2742),
.Y(n_2958)
);

INVxp67_ASAP7_75t_SL g2959 ( 
.A(n_2713),
.Y(n_2959)
);

XOR2x2_ASAP7_75t_L g2960 ( 
.A(n_2836),
.B(n_384),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2701),
.Y(n_2961)
);

INVxp67_ASAP7_75t_L g2962 ( 
.A(n_2773),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2734),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2835),
.B(n_382),
.Y(n_2964)
);

OAI22xp5_ASAP7_75t_L g2965 ( 
.A1(n_2807),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_2965)
);

OR2x2_ASAP7_75t_L g2966 ( 
.A(n_2781),
.B(n_385),
.Y(n_2966)
);

BUFx3_ASAP7_75t_L g2967 ( 
.A(n_2693),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2867),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2704),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2710),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2838),
.B(n_386),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2840),
.B(n_387),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2761),
.Y(n_2973)
);

OR2x2_ASAP7_75t_L g2974 ( 
.A(n_2785),
.B(n_388),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2736),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2745),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2841),
.Y(n_2977)
);

AND4x1_ASAP7_75t_L g2978 ( 
.A(n_2819),
.B(n_2855),
.C(n_2842),
.D(n_2850),
.Y(n_2978)
);

A2O1A1Ixp33_ASAP7_75t_L g2979 ( 
.A1(n_2804),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2717),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2762),
.Y(n_2981)
);

AOI22xp5_ASAP7_75t_L g2982 ( 
.A1(n_2837),
.A2(n_393),
.B1(n_390),
.B2(n_392),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2690),
.Y(n_2983)
);

OAI21xp33_ASAP7_75t_L g2984 ( 
.A1(n_2719),
.A2(n_393),
.B(n_394),
.Y(n_2984)
);

AOI22xp33_ASAP7_75t_L g2985 ( 
.A1(n_2715),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_2985)
);

OR2x2_ASAP7_75t_L g2986 ( 
.A(n_2786),
.B(n_395),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2832),
.Y(n_2987)
);

INVx1_ASAP7_75t_SL g2988 ( 
.A(n_2802),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2849),
.B(n_397),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2861),
.Y(n_2990)
);

INVxp67_ASAP7_75t_L g2991 ( 
.A(n_2746),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2848),
.Y(n_2992)
);

AND2x4_ASAP7_75t_L g2993 ( 
.A(n_2723),
.B(n_398),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2872),
.Y(n_2994)
);

OR2x2_ASAP7_75t_L g2995 ( 
.A(n_2751),
.B(n_399),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2873),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2851),
.B(n_399),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2874),
.Y(n_2998)
);

INVxp67_ASAP7_75t_SL g2999 ( 
.A(n_2866),
.Y(n_2999)
);

OR2x6_ASAP7_75t_L g3000 ( 
.A(n_2853),
.B(n_400),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2770),
.Y(n_3001)
);

INVxp67_ASAP7_75t_L g3002 ( 
.A(n_2747),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2730),
.Y(n_3003)
);

AND2x2_ASAP7_75t_L g3004 ( 
.A(n_2854),
.B(n_2858),
.Y(n_3004)
);

OR2x2_ASAP7_75t_L g3005 ( 
.A(n_2752),
.B(n_401),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2721),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2859),
.B(n_401),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2756),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2862),
.B(n_402),
.Y(n_3009)
);

OA222x2_ASAP7_75t_L g3010 ( 
.A1(n_2720),
.A2(n_407),
.B1(n_409),
.B2(n_403),
.C1(n_405),
.C2(n_408),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2863),
.Y(n_3011)
);

AND2x2_ASAP7_75t_L g3012 ( 
.A(n_2869),
.B(n_403),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2731),
.Y(n_3013)
);

INVx1_ASAP7_75t_SL g3014 ( 
.A(n_2705),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2726),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2692),
.B(n_407),
.Y(n_3016)
);

OAI22xp33_ASAP7_75t_SL g3017 ( 
.A1(n_2793),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_3017)
);

NAND2x1_ASAP7_75t_L g3018 ( 
.A(n_2953),
.B(n_2687),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2999),
.B(n_2879),
.Y(n_3019)
);

AND2x4_ASAP7_75t_L g3020 ( 
.A(n_2920),
.B(n_2754),
.Y(n_3020)
);

HB1xp67_ASAP7_75t_L g3021 ( 
.A(n_2883),
.Y(n_3021)
);

OR2x2_ASAP7_75t_L g3022 ( 
.A(n_2891),
.B(n_2702),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2958),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_3004),
.B(n_2801),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2939),
.B(n_2706),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2881),
.Y(n_3026)
);

AOI22xp5_ASAP7_75t_L g3027 ( 
.A1(n_2899),
.A2(n_2808),
.B1(n_2805),
.B2(n_2815),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2963),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2988),
.B(n_2722),
.Y(n_3029)
);

HB1xp67_ASAP7_75t_L g3030 ( 
.A(n_2900),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2926),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_3011),
.B(n_2725),
.Y(n_3032)
);

INVx2_ASAP7_75t_SL g3033 ( 
.A(n_2967),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_3014),
.B(n_2695),
.Y(n_3034)
);

OR2x2_ASAP7_75t_L g3035 ( 
.A(n_2975),
.B(n_2709),
.Y(n_3035)
);

INVx1_ASAP7_75t_SL g3036 ( 
.A(n_2960),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2977),
.B(n_2696),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2973),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2919),
.B(n_2887),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2884),
.Y(n_3040)
);

AOI21xp33_ASAP7_75t_SL g3041 ( 
.A1(n_2880),
.A2(n_2809),
.B(n_2795),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2885),
.Y(n_3042)
);

HB1xp67_ASAP7_75t_L g3043 ( 
.A(n_2948),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2993),
.Y(n_3044)
);

AND2x2_ASAP7_75t_L g3045 ( 
.A(n_2929),
.B(n_2728),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2925),
.B(n_2733),
.Y(n_3046)
);

INVx2_ASAP7_75t_SL g3047 ( 
.A(n_2993),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_3008),
.Y(n_3048)
);

INVx1_ASAP7_75t_SL g3049 ( 
.A(n_2964),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2888),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2890),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2896),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2897),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2968),
.B(n_2739),
.Y(n_3054)
);

AOI22xp5_ASAP7_75t_L g3055 ( 
.A1(n_2959),
.A2(n_2904),
.B1(n_2913),
.B2(n_2923),
.Y(n_3055)
);

OR2x2_ASAP7_75t_L g3056 ( 
.A(n_2990),
.B(n_2716),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2914),
.B(n_2700),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2898),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2893),
.B(n_2764),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2901),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2877),
.B(n_2878),
.Y(n_3061)
);

OR2x2_ASAP7_75t_L g3062 ( 
.A(n_2962),
.B(n_2703),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2908),
.Y(n_3063)
);

OA21x2_ASAP7_75t_L g3064 ( 
.A1(n_2892),
.A2(n_2978),
.B(n_2882),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_3013),
.B(n_2769),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2909),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2991),
.B(n_2771),
.Y(n_3067)
);

AOI22xp33_ASAP7_75t_L g3068 ( 
.A1(n_2976),
.A2(n_2799),
.B1(n_2775),
.B2(n_2814),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_2895),
.B(n_2777),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2910),
.Y(n_3070)
);

INVxp67_ASAP7_75t_L g3071 ( 
.A(n_2956),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_3002),
.B(n_2779),
.Y(n_3072)
);

OR2x2_ASAP7_75t_L g3073 ( 
.A(n_3015),
.B(n_2748),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2911),
.Y(n_3074)
);

OR2x2_ASAP7_75t_L g3075 ( 
.A(n_2983),
.B(n_2766),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2907),
.B(n_2987),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2912),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2992),
.B(n_2787),
.Y(n_3078)
);

OR2x2_ASAP7_75t_L g3079 ( 
.A(n_2994),
.B(n_2772),
.Y(n_3079)
);

NAND2xp33_ASAP7_75t_SL g3080 ( 
.A(n_2971),
.B(n_2796),
.Y(n_3080)
);

AND2x2_ASAP7_75t_L g3081 ( 
.A(n_2996),
.B(n_2783),
.Y(n_3081)
);

OR2x2_ASAP7_75t_L g3082 ( 
.A(n_2998),
.B(n_2774),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_SL g3083 ( 
.A(n_3006),
.B(n_2708),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2927),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_3012),
.B(n_2789),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2966),
.B(n_2763),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2974),
.B(n_2714),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2931),
.Y(n_3088)
);

INVxp67_ASAP7_75t_L g3089 ( 
.A(n_2986),
.Y(n_3089)
);

AOI22xp33_ASAP7_75t_SL g3090 ( 
.A1(n_3017),
.A2(n_2930),
.B1(n_2981),
.B2(n_2980),
.Y(n_3090)
);

OAI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_2906),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_3016),
.B(n_413),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2995),
.B(n_414),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2932),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2934),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_3005),
.B(n_414),
.Y(n_3096)
);

OAI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_2982),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_2905),
.B(n_2944),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_3021),
.Y(n_3099)
);

OAI31xp33_ASAP7_75t_L g3100 ( 
.A1(n_3057),
.A2(n_2979),
.A3(n_2955),
.B(n_2886),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_3043),
.Y(n_3101)
);

AOI22xp33_ASAP7_75t_L g3102 ( 
.A1(n_3064),
.A2(n_3001),
.B1(n_2947),
.B2(n_2951),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_3019),
.Y(n_3103)
);

AOI21xp33_ASAP7_75t_L g3104 ( 
.A1(n_3064),
.A2(n_3003),
.B(n_2970),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_3030),
.Y(n_3105)
);

AOI221xp5_ASAP7_75t_L g3106 ( 
.A1(n_3090),
.A2(n_2945),
.B1(n_2965),
.B2(n_2915),
.C(n_2984),
.Y(n_3106)
);

AOI22xp5_ASAP7_75t_L g3107 ( 
.A1(n_3098),
.A2(n_2937),
.B1(n_2933),
.B2(n_2957),
.Y(n_3107)
);

OA21x2_ASAP7_75t_SL g3108 ( 
.A1(n_3076),
.A2(n_2922),
.B(n_2921),
.Y(n_3108)
);

INVx2_ASAP7_75t_SL g3109 ( 
.A(n_3045),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_3073),
.Y(n_3110)
);

OA21x2_ASAP7_75t_L g3111 ( 
.A1(n_3055),
.A2(n_2942),
.B(n_2918),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_3049),
.B(n_2916),
.Y(n_3112)
);

INVx2_ASAP7_75t_SL g3113 ( 
.A(n_3046),
.Y(n_3113)
);

OAI221xp5_ASAP7_75t_L g3114 ( 
.A1(n_3086),
.A2(n_2952),
.B1(n_2950),
.B2(n_2936),
.C(n_3000),
.Y(n_3114)
);

NAND4xp25_ASAP7_75t_SL g3115 ( 
.A(n_3027),
.B(n_2943),
.C(n_2917),
.D(n_2928),
.Y(n_3115)
);

OAI32xp33_ASAP7_75t_L g3116 ( 
.A1(n_3080),
.A2(n_2924),
.A3(n_2989),
.B1(n_2972),
.B2(n_2946),
.Y(n_3116)
);

AND2x2_ASAP7_75t_L g3117 ( 
.A(n_3024),
.B(n_2935),
.Y(n_3117)
);

OAI221xp5_ASAP7_75t_L g3118 ( 
.A1(n_3036),
.A2(n_3000),
.B1(n_2889),
.B2(n_2985),
.C(n_2894),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_3078),
.B(n_3085),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_3069),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_3079),
.Y(n_3121)
);

AOI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_3071),
.A2(n_2997),
.B1(n_3009),
.B2(n_3007),
.Y(n_3122)
);

AOI21xp33_ASAP7_75t_L g3123 ( 
.A1(n_3022),
.A2(n_2969),
.B(n_2940),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_3082),
.Y(n_3124)
);

NOR2xp33_ASAP7_75t_L g3125 ( 
.A(n_3047),
.B(n_2938),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_3032),
.Y(n_3126)
);

HB1xp67_ASAP7_75t_L g3127 ( 
.A(n_3020),
.Y(n_3127)
);

INVxp67_ASAP7_75t_L g3128 ( 
.A(n_3033),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_3054),
.Y(n_3129)
);

AOI22xp5_ASAP7_75t_L g3130 ( 
.A1(n_3089),
.A2(n_3010),
.B1(n_2949),
.B2(n_2954),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_3075),
.Y(n_3131)
);

INVx3_ASAP7_75t_L g3132 ( 
.A(n_3020),
.Y(n_3132)
);

OAI32xp33_ASAP7_75t_L g3133 ( 
.A1(n_3062),
.A2(n_2941),
.A3(n_2961),
.B1(n_2903),
.B2(n_2902),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_3025),
.B(n_415),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_3081),
.B(n_417),
.Y(n_3135)
);

AOI21xp33_ASAP7_75t_L g3136 ( 
.A1(n_3028),
.A2(n_3056),
.B(n_3023),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_3044),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_3026),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_3040),
.Y(n_3139)
);

INVx1_ASAP7_75t_SL g3140 ( 
.A(n_3092),
.Y(n_3140)
);

AOI21xp33_ASAP7_75t_L g3141 ( 
.A1(n_3048),
.A2(n_418),
.B(n_419),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_3059),
.B(n_418),
.Y(n_3142)
);

INVx1_ASAP7_75t_SL g3143 ( 
.A(n_3029),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_3042),
.Y(n_3144)
);

NOR3xp33_ASAP7_75t_L g3145 ( 
.A(n_3041),
.B(n_419),
.C(n_420),
.Y(n_3145)
);

INVx1_ASAP7_75t_SL g3146 ( 
.A(n_3065),
.Y(n_3146)
);

AOI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_3087),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_3050),
.Y(n_3148)
);

OAI21xp33_ASAP7_75t_L g3149 ( 
.A1(n_3039),
.A2(n_421),
.B(n_422),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_3051),
.Y(n_3150)
);

INVx3_ASAP7_75t_L g3151 ( 
.A(n_3031),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_3067),
.B(n_423),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_3018),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_3072),
.B(n_424),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_3061),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3052),
.Y(n_3156)
);

AOI32xp33_ASAP7_75t_L g3157 ( 
.A1(n_3091),
.A2(n_428),
.A3(n_425),
.B1(n_427),
.B2(n_429),
.Y(n_3157)
);

OAI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_3097),
.A2(n_425),
.B(n_427),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_3127),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3135),
.Y(n_3160)
);

AND2x2_ASAP7_75t_L g3161 ( 
.A(n_3132),
.B(n_3035),
.Y(n_3161)
);

AOI21xp33_ASAP7_75t_L g3162 ( 
.A1(n_3102),
.A2(n_3038),
.B(n_3053),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_3128),
.B(n_3083),
.Y(n_3163)
);

INVxp67_ASAP7_75t_L g3164 ( 
.A(n_3134),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_3140),
.B(n_3034),
.Y(n_3165)
);

INVx1_ASAP7_75t_SL g3166 ( 
.A(n_3119),
.Y(n_3166)
);

AOI22xp5_ASAP7_75t_L g3167 ( 
.A1(n_3130),
.A2(n_3037),
.B1(n_3068),
.B2(n_3093),
.Y(n_3167)
);

NAND2xp33_ASAP7_75t_SL g3168 ( 
.A(n_3113),
.B(n_3058),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3105),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_3099),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_3117),
.B(n_3060),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_3101),
.Y(n_3172)
);

OAI33xp33_ASAP7_75t_L g3173 ( 
.A1(n_3110),
.A2(n_3074),
.A3(n_3066),
.B1(n_3077),
.B2(n_3070),
.B3(n_3063),
.Y(n_3173)
);

AOI22xp5_ASAP7_75t_L g3174 ( 
.A1(n_3106),
.A2(n_3096),
.B1(n_3088),
.B2(n_3094),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3142),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_3152),
.Y(n_3176)
);

AOI221xp5_ASAP7_75t_L g3177 ( 
.A1(n_3104),
.A2(n_3136),
.B1(n_3133),
.B2(n_3116),
.C(n_3123),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3154),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_3145),
.B(n_3084),
.Y(n_3179)
);

AOI22xp33_ASAP7_75t_L g3180 ( 
.A1(n_3115),
.A2(n_3095),
.B1(n_431),
.B2(n_429),
.Y(n_3180)
);

OAI21xp33_ASAP7_75t_L g3181 ( 
.A1(n_3151),
.A2(n_430),
.B(n_431),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3121),
.Y(n_3182)
);

O2A1O1Ixp33_ASAP7_75t_L g3183 ( 
.A1(n_3100),
.A2(n_434),
.B(n_432),
.C(n_433),
.Y(n_3183)
);

INVxp67_ASAP7_75t_SL g3184 ( 
.A(n_3153),
.Y(n_3184)
);

OAI22xp5_ASAP7_75t_L g3185 ( 
.A1(n_3114),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_3124),
.Y(n_3186)
);

NAND2xp33_ASAP7_75t_L g3187 ( 
.A(n_3109),
.B(n_513),
.Y(n_3187)
);

OAI221xp5_ASAP7_75t_SL g3188 ( 
.A1(n_3108),
.A2(n_3146),
.B1(n_3143),
.B2(n_3107),
.C(n_3131),
.Y(n_3188)
);

NOR3xp33_ASAP7_75t_L g3189 ( 
.A(n_3103),
.B(n_514),
.C(n_515),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_3137),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_3112),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_3129),
.B(n_516),
.Y(n_3192)
);

OAI22xp5_ASAP7_75t_L g3193 ( 
.A1(n_3120),
.A2(n_521),
.B1(n_517),
.B2(n_520),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3126),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3155),
.B(n_522),
.Y(n_3195)
);

OAI21xp33_ASAP7_75t_SL g3196 ( 
.A1(n_3125),
.A2(n_525),
.B(n_527),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3159),
.Y(n_3197)
);

AOI22xp33_ASAP7_75t_L g3198 ( 
.A1(n_3177),
.A2(n_3111),
.B1(n_3118),
.B2(n_3122),
.Y(n_3198)
);

INVxp67_ASAP7_75t_L g3199 ( 
.A(n_3161),
.Y(n_3199)
);

A2O1A1Ixp33_ASAP7_75t_L g3200 ( 
.A1(n_3188),
.A2(n_3158),
.B(n_3149),
.C(n_3157),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_3165),
.Y(n_3201)
);

INVx1_ASAP7_75t_SL g3202 ( 
.A(n_3166),
.Y(n_3202)
);

OR2x2_ASAP7_75t_L g3203 ( 
.A(n_3171),
.B(n_3111),
.Y(n_3203)
);

NOR4xp25_ASAP7_75t_L g3204 ( 
.A(n_3183),
.B(n_3139),
.C(n_3144),
.D(n_3138),
.Y(n_3204)
);

AOI21xp33_ASAP7_75t_SL g3205 ( 
.A1(n_3163),
.A2(n_3141),
.B(n_3156),
.Y(n_3205)
);

AOI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3167),
.A2(n_3147),
.B1(n_3150),
.B2(n_3148),
.Y(n_3206)
);

AND2x2_ASAP7_75t_L g3207 ( 
.A(n_3184),
.B(n_528),
.Y(n_3207)
);

NOR2xp33_ASAP7_75t_L g3208 ( 
.A(n_3164),
.B(n_529),
.Y(n_3208)
);

A2O1A1Ixp33_ASAP7_75t_L g3209 ( 
.A1(n_3196),
.A2(n_3162),
.B(n_3180),
.C(n_3174),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_3187),
.A2(n_530),
.B(n_531),
.Y(n_3210)
);

NOR2xp67_ASAP7_75t_L g3211 ( 
.A(n_3194),
.B(n_532),
.Y(n_3211)
);

A2O1A1Ixp33_ASAP7_75t_L g3212 ( 
.A1(n_3179),
.A2(n_536),
.B(n_533),
.C(n_535),
.Y(n_3212)
);

AOI221xp5_ASAP7_75t_L g3213 ( 
.A1(n_3176),
.A2(n_540),
.B1(n_537),
.B2(n_539),
.C(n_541),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_3175),
.B(n_544),
.Y(n_3214)
);

AOI221xp5_ASAP7_75t_L g3215 ( 
.A1(n_3178),
.A2(n_548),
.B1(n_545),
.B2(n_546),
.C(n_551),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_3160),
.B(n_870),
.Y(n_3216)
);

O2A1O1Ixp33_ASAP7_75t_L g3217 ( 
.A1(n_3185),
.A2(n_557),
.B(n_553),
.C(n_554),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_3190),
.Y(n_3218)
);

OAI221xp5_ASAP7_75t_L g3219 ( 
.A1(n_3191),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.C(n_561),
.Y(n_3219)
);

NAND4xp25_ASAP7_75t_L g3220 ( 
.A(n_3168),
.B(n_565),
.C(n_563),
.D(n_564),
.Y(n_3220)
);

OAI21xp5_ASAP7_75t_SL g3221 ( 
.A1(n_3182),
.A2(n_567),
.B(n_569),
.Y(n_3221)
);

AOI32xp33_ASAP7_75t_L g3222 ( 
.A1(n_3186),
.A2(n_575),
.A3(n_571),
.B1(n_573),
.B2(n_576),
.Y(n_3222)
);

NAND4xp25_ASAP7_75t_L g3223 ( 
.A(n_3169),
.B(n_581),
.C(n_578),
.D(n_579),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3170),
.Y(n_3224)
);

AOI21xp5_ASAP7_75t_L g3225 ( 
.A1(n_3173),
.A2(n_583),
.B(n_585),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_SL g3226 ( 
.A(n_3172),
.B(n_586),
.Y(n_3226)
);

AOI22xp33_ASAP7_75t_L g3227 ( 
.A1(n_3189),
.A2(n_593),
.B1(n_587),
.B2(n_590),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_3192),
.Y(n_3228)
);

OA211x2_ASAP7_75t_L g3229 ( 
.A1(n_3181),
.A2(n_596),
.B(n_594),
.C(n_595),
.Y(n_3229)
);

AOI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_3195),
.A2(n_3193),
.B1(n_602),
.B2(n_598),
.Y(n_3230)
);

AOI322xp5_ASAP7_75t_L g3231 ( 
.A1(n_3177),
.A2(n_610),
.A3(n_608),
.B1(n_604),
.B2(n_600),
.C1(n_603),
.C2(n_607),
.Y(n_3231)
);

OAI221xp5_ASAP7_75t_L g3232 ( 
.A1(n_3188),
.A2(n_614),
.B1(n_611),
.B2(n_613),
.C(n_615),
.Y(n_3232)
);

NOR4xp25_ASAP7_75t_L g3233 ( 
.A(n_3188),
.B(n_619),
.C(n_617),
.D(n_618),
.Y(n_3233)
);

AND2x2_ASAP7_75t_L g3234 ( 
.A(n_3202),
.B(n_620),
.Y(n_3234)
);

NAND3xp33_ASAP7_75t_L g3235 ( 
.A(n_3198),
.B(n_621),
.C(n_622),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3199),
.Y(n_3236)
);

INVx2_ASAP7_75t_SL g3237 ( 
.A(n_3203),
.Y(n_3237)
);

NOR3xp33_ASAP7_75t_L g3238 ( 
.A(n_3232),
.B(n_624),
.C(n_627),
.Y(n_3238)
);

AOI211xp5_ASAP7_75t_L g3239 ( 
.A1(n_3233),
.A2(n_630),
.B(n_628),
.C(n_629),
.Y(n_3239)
);

AOI221xp5_ASAP7_75t_L g3240 ( 
.A1(n_3204),
.A2(n_633),
.B1(n_631),
.B2(n_632),
.C(n_635),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3207),
.B(n_636),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_3208),
.B(n_637),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3197),
.Y(n_3243)
);

NOR2x1p5_ASAP7_75t_L g3244 ( 
.A(n_3201),
.B(n_639),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_3200),
.B(n_640),
.Y(n_3245)
);

AOI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_3209),
.A2(n_641),
.B(n_642),
.Y(n_3246)
);

OAI21xp33_ASAP7_75t_L g3247 ( 
.A1(n_3206),
.A2(n_643),
.B(n_647),
.Y(n_3247)
);

NAND2xp33_ASAP7_75t_L g3248 ( 
.A(n_3224),
.B(n_648),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3214),
.Y(n_3249)
);

AND3x4_ASAP7_75t_L g3250 ( 
.A(n_3228),
.B(n_649),
.C(n_650),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3216),
.Y(n_3251)
);

AOI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_3225),
.A2(n_651),
.B(n_653),
.Y(n_3252)
);

NOR2xp33_ASAP7_75t_L g3253 ( 
.A(n_3205),
.B(n_3218),
.Y(n_3253)
);

NOR3x1_ASAP7_75t_L g3254 ( 
.A(n_3220),
.B(n_656),
.C(n_657),
.Y(n_3254)
);

INVxp67_ASAP7_75t_SL g3255 ( 
.A(n_3226),
.Y(n_3255)
);

AOI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_3221),
.A2(n_658),
.B(n_660),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3231),
.B(n_662),
.Y(n_3257)
);

OAI21xp5_ASAP7_75t_L g3258 ( 
.A1(n_3240),
.A2(n_3210),
.B(n_3217),
.Y(n_3258)
);

NOR3xp33_ASAP7_75t_L g3259 ( 
.A(n_3237),
.B(n_3212),
.C(n_3219),
.Y(n_3259)
);

NAND4xp25_ASAP7_75t_L g3260 ( 
.A(n_3253),
.B(n_3229),
.C(n_3223),
.D(n_3230),
.Y(n_3260)
);

OAI21xp33_ASAP7_75t_SL g3261 ( 
.A1(n_3236),
.A2(n_3211),
.B(n_3222),
.Y(n_3261)
);

NOR2x1_ASAP7_75t_L g3262 ( 
.A(n_3243),
.B(n_3213),
.Y(n_3262)
);

NAND4xp25_ASAP7_75t_L g3263 ( 
.A(n_3246),
.B(n_3227),
.C(n_3215),
.D(n_666),
.Y(n_3263)
);

OAI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_3252),
.A2(n_664),
.B(n_665),
.Y(n_3264)
);

NOR2x1p5_ASAP7_75t_L g3265 ( 
.A(n_3255),
.B(n_670),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3234),
.B(n_3249),
.Y(n_3266)
);

NAND3xp33_ASAP7_75t_L g3267 ( 
.A(n_3248),
.B(n_671),
.C(n_672),
.Y(n_3267)
);

AOI211x1_ASAP7_75t_L g3268 ( 
.A1(n_3235),
.A2(n_677),
.B(n_673),
.C(n_674),
.Y(n_3268)
);

NOR3xp33_ASAP7_75t_L g3269 ( 
.A(n_3245),
.B(n_678),
.C(n_679),
.Y(n_3269)
);

NOR3xp33_ASAP7_75t_L g3270 ( 
.A(n_3261),
.B(n_3251),
.C(n_3247),
.Y(n_3270)
);

NOR2xp67_ASAP7_75t_L g3271 ( 
.A(n_3260),
.B(n_3257),
.Y(n_3271)
);

AND2x4_ASAP7_75t_L g3272 ( 
.A(n_3262),
.B(n_3244),
.Y(n_3272)
);

NOR3xp33_ASAP7_75t_L g3273 ( 
.A(n_3266),
.B(n_3241),
.C(n_3242),
.Y(n_3273)
);

OR2x2_ASAP7_75t_L g3274 ( 
.A(n_3259),
.B(n_3256),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3272),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3274),
.Y(n_3276)
);

AOI22xp5_ASAP7_75t_L g3277 ( 
.A1(n_3276),
.A2(n_3271),
.B1(n_3270),
.B2(n_3273),
.Y(n_3277)
);

OAI21xp5_ASAP7_75t_SL g3278 ( 
.A1(n_3275),
.A2(n_3258),
.B(n_3263),
.Y(n_3278)
);

BUFx2_ASAP7_75t_L g3279 ( 
.A(n_3277),
.Y(n_3279)
);

NAND2xp33_ASAP7_75t_R g3280 ( 
.A(n_3278),
.B(n_3264),
.Y(n_3280)
);

AOI31xp33_ASAP7_75t_L g3281 ( 
.A1(n_3277),
.A2(n_3239),
.A3(n_3267),
.B(n_3265),
.Y(n_3281)
);

OR2x2_ASAP7_75t_L g3282 ( 
.A(n_3279),
.B(n_3269),
.Y(n_3282)
);

HB1xp67_ASAP7_75t_SL g3283 ( 
.A(n_3280),
.Y(n_3283)
);

XNOR2x1_ASAP7_75t_L g3284 ( 
.A(n_3281),
.B(n_3250),
.Y(n_3284)
);

INVx2_ASAP7_75t_SL g3285 ( 
.A(n_3284),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3283),
.Y(n_3286)
);

XOR2xp5_ASAP7_75t_L g3287 ( 
.A(n_3286),
.B(n_3282),
.Y(n_3287)
);

OR2x2_ASAP7_75t_L g3288 ( 
.A(n_3287),
.B(n_3285),
.Y(n_3288)
);

XNOR2x1_ASAP7_75t_L g3289 ( 
.A(n_3288),
.B(n_3268),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3289),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3290),
.B(n_3254),
.Y(n_3291)
);

AOI322xp5_ASAP7_75t_L g3292 ( 
.A1(n_3291),
.A2(n_3238),
.A3(n_682),
.B1(n_683),
.B2(n_685),
.C1(n_687),
.C2(n_689),
.Y(n_3292)
);

AOI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_3292),
.A2(n_692),
.B1(n_681),
.B2(n_690),
.Y(n_3293)
);

AOI211xp5_ASAP7_75t_L g3294 ( 
.A1(n_3293),
.A2(n_698),
.B(n_695),
.C(n_697),
.Y(n_3294)
);


endmodule