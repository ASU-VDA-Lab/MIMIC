module fake_netlist_6_344_n_2026 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2026);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2026;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1774;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1475;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_15),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_12),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_204),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_22),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_2),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_40),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_128),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_126),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_200),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_122),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_172),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_143),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_50),
.Y(n_222)
);

BUFx8_ASAP7_75t_SL g223 ( 
.A(n_97),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_82),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_43),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_65),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_35),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_121),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_125),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_170),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_153),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_103),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_198),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_165),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_206),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_105),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_114),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_79),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_8),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_148),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_71),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_76),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_137),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_23),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_140),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_168),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_2),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_149),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_80),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_5),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_156),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_41),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_42),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_34),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_64),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_46),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_151),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_157),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_96),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_93),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_164),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_85),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_67),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_107),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_63),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_117),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_205),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_32),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_70),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_20),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_43),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_77),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_67),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_202),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_72),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_141),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_110),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_57),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_94),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_1),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_174),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_196),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_83),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_127),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_65),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_150),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_138),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_23),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_53),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_120),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_90),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_46),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_33),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_135),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_11),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_5),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_142),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_180),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_136),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_109),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_41),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_186),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_147),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_44),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_19),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_166),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_145),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_194),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_146),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_178),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_102),
.Y(n_314)
);

INVx4_ASAP7_75t_R g315 ( 
.A(n_181),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_188),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_118),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_27),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_8),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_19),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_81),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_74),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_38),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_171),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_163),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_69),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_38),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_57),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_173),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_100),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_3),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_42),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_25),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_189),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_32),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_76),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_51),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_6),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_45),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_30),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_139),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_160),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_144),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_31),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_24),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_91),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_201),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_50),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_20),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_60),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_169),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_175),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_7),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_191),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_119),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_29),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_7),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_87),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_66),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_183),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_26),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_31),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_184),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_89),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_61),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_24),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_40),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_35),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_134),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_36),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_60),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_48),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_129),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_73),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_28),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_84),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_45),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_28),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_179),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_25),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_52),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_155),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_53),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_152),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_158),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_26),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_75),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_190),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_113),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_4),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_47),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_106),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_116),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_1),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_75),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_70),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_185),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_61),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_92),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_71),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_37),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_69),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_98),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_0),
.Y(n_404)
);

INVxp33_ASAP7_75t_SL g405 ( 
.A(n_3),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_62),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_22),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_15),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_132),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_88),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_162),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_233),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_230),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_257),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_238),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_257),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_227),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_257),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_257),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_247),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_240),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_257),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_257),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_230),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_257),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_241),
.B(n_0),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_257),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_257),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g429 ( 
.A(n_222),
.B(n_4),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_226),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_221),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_241),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_243),
.B(n_6),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_263),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_221),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_232),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_400),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_357),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_357),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_314),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_370),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_232),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_236),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_236),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_248),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_370),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_209),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_211),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_224),
.B(n_9),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_213),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_225),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_346),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_244),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_248),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_246),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_384),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_260),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_260),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_261),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_261),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_223),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_284),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_249),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_284),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_256),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_258),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_265),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_207),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_250),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_285),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_299),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_277),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_210),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_285),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_283),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_302),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_212),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_288),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_295),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_296),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_302),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_305),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_305),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_306),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_215),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_306),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_313),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_208),
.B(n_9),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_298),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_282),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g491 ( 
.A(n_208),
.B(n_10),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_304),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_292),
.B(n_10),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_313),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_308),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_216),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_217),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_318),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_320),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_322),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_323),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_321),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_218),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_219),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_326),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_321),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_220),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_228),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_224),
.B(n_11),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_229),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_231),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_328),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_214),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_325),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_331),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_335),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_337),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_234),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_325),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_417),
.B(n_310),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_461),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_SL g522 ( 
.A(n_509),
.B(n_417),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_282),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_513),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_468),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_416),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_431),
.B(n_282),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_418),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_438),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_416),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_412),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_419),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_473),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_477),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_422),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_423),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_425),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_490),
.B(n_214),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_R g540 ( 
.A(n_447),
.B(n_405),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_435),
.B(n_303),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_490),
.B(n_254),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_427),
.B(n_214),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_428),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_485),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_426),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_496),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_497),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_421),
.B(n_469),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_436),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_442),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_443),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_444),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_R g554 ( 
.A(n_503),
.B(n_235),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_445),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_504),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_507),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_R g558 ( 
.A(n_508),
.B(n_237),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_415),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_519),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_454),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_510),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_457),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_458),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_459),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_460),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_462),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_511),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_464),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_518),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_470),
.B(n_214),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_474),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_476),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_481),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_482),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_483),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_447),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_484),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_487),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_448),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_494),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_502),
.B(n_214),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_420),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_413),
.B(n_254),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_506),
.B(n_303),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_514),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_426),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_438),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_SL g590 ( 
.A(n_437),
.B(n_214),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_449),
.B(n_355),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_448),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_433),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_433),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_450),
.B(n_411),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_450),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_488),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_451),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_451),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_437),
.B(n_251),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_424),
.B(n_254),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_453),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_453),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_491),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_432),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_591),
.B(n_262),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_525),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_527),
.Y(n_608)
);

AND2x6_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_262),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_532),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_600),
.B(n_546),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_594),
.B(n_430),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_546),
.B(n_455),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_527),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_531),
.Y(n_615)
);

AO22x2_ASAP7_75t_L g616 ( 
.A1(n_546),
.A2(n_309),
.B1(n_262),
.B2(n_252),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_595),
.A2(n_441),
.B1(n_439),
.B2(n_455),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_531),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_525),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_594),
.B(n_316),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_546),
.A2(n_365),
.B1(n_327),
.B2(n_348),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_529),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_589),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_577),
.B(n_446),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_542),
.B(n_465),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_529),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_530),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_533),
.B(n_463),
.Y(n_628)
);

OAI22xp33_ASAP7_75t_L g629 ( 
.A1(n_594),
.A2(n_340),
.B1(n_471),
.B2(n_441),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_595),
.B(n_463),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_599),
.B(n_466),
.Y(n_631)
);

BUFx4f_ASAP7_75t_L g632 ( 
.A(n_538),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_527),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_554),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_603),
.B(n_466),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_599),
.B(n_467),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_599),
.B(n_467),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_533),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_536),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_L g641 ( 
.A1(n_540),
.A2(n_439),
.B1(n_429),
.B2(n_349),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_R g642 ( 
.A(n_530),
.B(n_472),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_542),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_599),
.B(n_603),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_603),
.B(n_475),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_603),
.B(n_475),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_588),
.B(n_500),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_531),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_537),
.B(n_478),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_544),
.Y(n_650)
);

CKINVDCx14_ASAP7_75t_R g651 ( 
.A(n_558),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_599),
.B(n_309),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_605),
.B(n_478),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_605),
.B(n_528),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_531),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_599),
.B(n_479),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_544),
.B(n_479),
.Y(n_657)
);

BUFx4f_ASAP7_75t_L g658 ( 
.A(n_538),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_549),
.B(n_480),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_523),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_549),
.B(n_489),
.C(n_480),
.Y(n_661)
);

AND3x2_ASAP7_75t_L g662 ( 
.A(n_589),
.B(n_363),
.C(n_309),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_551),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_551),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_552),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_590),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_523),
.B(n_489),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_531),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_523),
.B(n_303),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_524),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_523),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_528),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_585),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_539),
.B(n_492),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_539),
.B(n_492),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_524),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_605),
.B(n_345),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_528),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_581),
.B(n_495),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_531),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_538),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_592),
.B(n_498),
.Y(n_682)
);

AND2x2_ASAP7_75t_SL g683 ( 
.A(n_541),
.B(n_286),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_552),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_541),
.B(n_586),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_541),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_585),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_588),
.B(n_498),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_596),
.B(n_499),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_522),
.A2(n_501),
.B1(n_516),
.B2(n_515),
.Y(n_690)
);

NOR2x1p5_ASAP7_75t_L g691 ( 
.A(n_598),
.B(n_499),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_541),
.B(n_586),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_602),
.B(n_501),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_550),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_593),
.B(n_505),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_550),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_550),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_520),
.B(n_512),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_593),
.A2(n_365),
.B1(n_292),
.B2(n_327),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_553),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_550),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_555),
.B(n_512),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_569),
.Y(n_703)
);

INVx6_ASAP7_75t_L g704 ( 
.A(n_586),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_601),
.A2(n_365),
.B1(n_356),
.B2(n_348),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_555),
.Y(n_706)
);

INVx5_ASAP7_75t_L g707 ( 
.A(n_538),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_601),
.B(n_515),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_597),
.B(n_517),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_526),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_559),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_534),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_563),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_538),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_564),
.B(n_517),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_564),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_597),
.B(n_310),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_560),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_569),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_560),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_560),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_574),
.B(n_264),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_566),
.B(n_345),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_604),
.A2(n_381),
.B1(n_350),
.B2(n_353),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_574),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_566),
.B(n_345),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_560),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_604),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_572),
.B(n_310),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_572),
.A2(n_359),
.B1(n_362),
.B2(n_339),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_573),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_573),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_535),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_576),
.A2(n_371),
.B1(n_386),
.B2(n_408),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_576),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_574),
.B(n_239),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_563),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_563),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_580),
.B(n_374),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_579),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_579),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_582),
.A2(n_365),
.B1(n_356),
.B2(n_383),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_582),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_580),
.B(n_434),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_565),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_580),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_565),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_565),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_545),
.B(n_310),
.Y(n_749)
);

AND2x2_ASAP7_75t_SL g750 ( 
.A(n_571),
.B(n_286),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_652),
.B(n_316),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_643),
.B(n_567),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_611),
.B(n_659),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_SL g754 ( 
.A(n_634),
.B(n_547),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_652),
.B(n_580),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_660),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_672),
.B(n_678),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_606),
.B(n_560),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_606),
.A2(n_609),
.B1(n_687),
.B2(n_683),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_632),
.A2(n_543),
.B(n_571),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_606),
.B(n_609),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_670),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_606),
.A2(n_440),
.B1(n_452),
.B2(n_456),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_632),
.A2(n_543),
.B(n_583),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_L g765 ( 
.A(n_630),
.B(n_556),
.C(n_548),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_660),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_606),
.B(n_561),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_702),
.B(n_367),
.C(n_366),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_643),
.B(n_567),
.Y(n_769)
);

INVx8_ASAP7_75t_L g770 ( 
.A(n_677),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_609),
.B(n_561),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_609),
.B(n_561),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_671),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_671),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_674),
.B(n_561),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_609),
.A2(n_290),
.B1(n_242),
.B2(n_409),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_685),
.Y(n_777)
);

AND2x6_ASAP7_75t_SL g778 ( 
.A(n_698),
.B(n_243),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_670),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_685),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_676),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_675),
.B(n_368),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_612),
.B(n_557),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_687),
.A2(n_287),
.B1(n_403),
.B2(n_245),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_692),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_654),
.B(n_567),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_654),
.B(n_575),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_692),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_612),
.B(n_562),
.Y(n_789)
);

NOR2x1p5_ASAP7_75t_L g790 ( 
.A(n_634),
.B(n_568),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_661),
.B(n_617),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_672),
.B(n_575),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_676),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_619),
.B(n_578),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_713),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_713),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_638),
.B(n_578),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_737),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_638),
.B(n_578),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_639),
.B(n_587),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_678),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_686),
.Y(n_802)
);

O2A1O1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_673),
.A2(n_583),
.B(n_587),
.C(n_383),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_628),
.B(n_372),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_750),
.B(n_316),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_649),
.B(n_375),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_639),
.B(n_587),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_640),
.B(n_607),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_737),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_623),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_686),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_750),
.A2(n_380),
.B1(n_291),
.B2(n_336),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_616),
.A2(n_380),
.B1(n_291),
.B2(n_336),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_704),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_738),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_657),
.B(n_378),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_663),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_664),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_665),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_684),
.Y(n_820)
);

BUFx6f_ASAP7_75t_SL g821 ( 
.A(n_728),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_SL g822 ( 
.A(n_624),
.B(n_570),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_653),
.B(n_390),
.C(n_387),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_635),
.B(n_316),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_738),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_640),
.B(n_329),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_622),
.B(n_329),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_626),
.B(n_650),
.Y(n_828)
);

OAI221xp5_ASAP7_75t_L g829 ( 
.A1(n_705),
.A2(n_493),
.B1(n_275),
.B2(n_272),
.C(n_344),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_745),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_732),
.B(n_376),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_645),
.B(n_316),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_704),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_745),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_688),
.B(n_395),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_632),
.A2(n_358),
.B(n_343),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_700),
.Y(n_837)
);

INVx8_ASAP7_75t_L g838 ( 
.A(n_677),
.Y(n_838)
);

O2A1O1Ixp5_ASAP7_75t_L g839 ( 
.A1(n_644),
.A2(n_343),
.B(n_410),
.C(n_358),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_688),
.B(n_396),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_695),
.B(n_401),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_732),
.B(n_376),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_747),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_L g844 ( 
.A(n_690),
.B(n_521),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_653),
.B(n_299),
.Y(n_845)
);

AOI221xp5_ASAP7_75t_L g846 ( 
.A1(n_629),
.A2(n_338),
.B1(n_332),
.B2(n_407),
.C(n_319),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_625),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_706),
.Y(n_848)
);

INVxp33_ASAP7_75t_L g849 ( 
.A(n_625),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_716),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_708),
.B(n_299),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_731),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_747),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_722),
.B(n_382),
.Y(n_854)
);

NOR3xp33_ASAP7_75t_L g855 ( 
.A(n_641),
.B(n_406),
.C(n_402),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_646),
.B(n_316),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_647),
.B(n_374),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_613),
.B(n_393),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_694),
.B(n_385),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_667),
.B(n_393),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_647),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_694),
.B(n_385),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_708),
.B(n_299),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_735),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_715),
.B(n_584),
.Y(n_865)
);

NOR2x1p5_ASAP7_75t_L g866 ( 
.A(n_715),
.B(n_374),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_748),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_696),
.B(n_385),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_748),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_709),
.B(n_399),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_741),
.B(n_389),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_704),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_608),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_627),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_743),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_696),
.B(n_385),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_623),
.B(n_740),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_746),
.B(n_410),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_631),
.B(n_636),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_637),
.B(n_253),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_651),
.B(n_280),
.Y(n_881)
);

O2A1O1Ixp5_ASAP7_75t_L g882 ( 
.A1(n_736),
.A2(n_404),
.B(n_398),
.C(n_255),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_697),
.B(n_259),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_697),
.B(n_701),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_701),
.B(n_266),
.Y(n_885)
);

AOI221xp5_ASAP7_75t_L g886 ( 
.A1(n_734),
.A2(n_404),
.B1(n_398),
.B2(n_255),
.C(n_394),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_648),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_SL g888 ( 
.A(n_710),
.B(n_268),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_658),
.A2(n_397),
.B(n_269),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_608),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_703),
.B(n_385),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_620),
.A2(n_394),
.B(n_267),
.C(n_391),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_703),
.B(n_274),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_616),
.A2(n_252),
.B1(n_391),
.B2(n_333),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_719),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_610),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_614),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_651),
.B(n_377),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_719),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_614),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_725),
.B(n_276),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_723),
.B(n_377),
.Y(n_902)
);

AND2x4_ASAP7_75t_SL g903 ( 
.A(n_677),
.B(n_267),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_725),
.B(n_278),
.Y(n_904)
);

NOR3xp33_ASAP7_75t_L g905 ( 
.A(n_744),
.B(n_270),
.C(n_271),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_739),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_739),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_610),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_669),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_666),
.B(n_385),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_656),
.B(n_279),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_770),
.B(n_710),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_753),
.B(n_858),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_753),
.B(n_666),
.Y(n_914)
);

AO21x1_ASAP7_75t_L g915 ( 
.A1(n_858),
.A2(n_749),
.B(n_669),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_906),
.B(n_669),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_777),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_758),
.A2(n_658),
.B(n_618),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_849),
.B(n_679),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_792),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_907),
.B(n_677),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_910),
.A2(n_717),
.B(n_729),
.C(n_730),
.Y(n_922)
);

NOR3xp33_ASAP7_75t_L g923 ( 
.A(n_846),
.B(n_689),
.C(n_682),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_849),
.B(n_693),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_755),
.A2(n_680),
.B(n_621),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_767),
.A2(n_615),
.B(n_714),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_792),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_782),
.B(n_680),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_762),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_782),
.B(n_616),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_860),
.B(n_804),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_860),
.B(n_616),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_771),
.A2(n_772),
.B(n_786),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_787),
.A2(n_681),
.B(n_714),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_910),
.A2(n_724),
.B(n_726),
.C(n_723),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_804),
.B(n_668),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_806),
.B(n_668),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_780),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_874),
.B(n_711),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_SL g940 ( 
.A(n_905),
.B(n_733),
.C(n_712),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_877),
.B(n_712),
.Y(n_941)
);

BUFx4f_ASAP7_75t_L g942 ( 
.A(n_770),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_814),
.A2(n_721),
.B(n_720),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_879),
.A2(n_642),
.B1(n_691),
.B2(n_718),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_806),
.B(n_668),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_SL g946 ( 
.A(n_754),
.B(n_733),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_814),
.A2(n_720),
.B(n_721),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_805),
.A2(n_726),
.B(n_699),
.C(n_742),
.Y(n_948)
);

OAI21xp33_ASAP7_75t_L g949 ( 
.A1(n_835),
.A2(n_270),
.B(n_271),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_762),
.Y(n_950)
);

OAI21xp33_ASAP7_75t_L g951 ( 
.A1(n_835),
.A2(n_840),
.B(n_841),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_775),
.A2(n_721),
.B(n_720),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_816),
.B(n_718),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_816),
.B(n_727),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_805),
.A2(n_633),
.B(n_273),
.C(n_272),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_824),
.A2(n_633),
.B(n_648),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_752),
.B(n_727),
.Y(n_957)
);

AO22x1_ASAP7_75t_L g958 ( 
.A1(n_841),
.A2(n_273),
.B1(n_275),
.B2(n_307),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_884),
.A2(n_727),
.B(n_361),
.Y(n_959)
);

NAND3xp33_ASAP7_75t_L g960 ( 
.A(n_840),
.B(n_662),
.C(n_289),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_752),
.B(n_648),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_751),
.A2(n_307),
.B(n_361),
.C(n_344),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_801),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_887),
.A2(n_655),
.B(n_707),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_810),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_783),
.B(n_655),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_769),
.B(n_655),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_845),
.B(n_333),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_861),
.B(n_377),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_870),
.A2(n_342),
.B(n_293),
.C(n_392),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_769),
.B(n_281),
.Y(n_971)
);

BUFx4f_ASAP7_75t_L g972 ( 
.A(n_770),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_757),
.B(n_78),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_812),
.A2(n_365),
.B1(n_388),
.B2(n_294),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_812),
.A2(n_365),
.B1(n_388),
.B2(n_297),
.Y(n_975)
);

BUFx12f_ASAP7_75t_L g976 ( 
.A(n_896),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_759),
.A2(n_388),
.B1(n_300),
.B2(n_347),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_813),
.A2(n_388),
.B1(n_301),
.B2(n_351),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_801),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_SL g980 ( 
.A(n_822),
.B(n_311),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_785),
.B(n_312),
.Y(n_981)
);

INVx11_ASAP7_75t_L g982 ( 
.A(n_908),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_813),
.A2(n_388),
.B1(n_379),
.B2(n_373),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_872),
.A2(n_369),
.B(n_364),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_801),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_872),
.A2(n_360),
.B(n_354),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_788),
.B(n_317),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_801),
.Y(n_988)
);

AO21x1_ASAP7_75t_L g989 ( 
.A1(n_856),
.A2(n_315),
.B(n_14),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_808),
.A2(n_352),
.B(n_341),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_833),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_760),
.A2(n_334),
.B(n_330),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_894),
.A2(n_324),
.B1(n_315),
.B2(n_16),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_764),
.A2(n_203),
.B(n_199),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_751),
.A2(n_193),
.B(n_187),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_828),
.A2(n_182),
.B(n_176),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_883),
.A2(n_167),
.B(n_161),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_885),
.A2(n_159),
.B(n_154),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_894),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_870),
.A2(n_17),
.B(n_18),
.C(n_21),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_882),
.A2(n_133),
.B(n_131),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_893),
.A2(n_904),
.B(n_901),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_789),
.B(n_17),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_829),
.A2(n_18),
.B(n_21),
.C(n_27),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_791),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_847),
.B(n_34),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_803),
.A2(n_130),
.B(n_124),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_902),
.B(n_104),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_888),
.B(n_36),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_886),
.A2(n_37),
.B1(n_39),
.B2(n_44),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_895),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_817),
.B(n_39),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_839),
.A2(n_123),
.B(n_115),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_779),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_899),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_779),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_866),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_909),
.A2(n_112),
.B(n_108),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_880),
.B(n_101),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_818),
.B(n_47),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_781),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_781),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_794),
.A2(n_99),
.B(n_95),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_768),
.B(n_48),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_823),
.B(n_49),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_865),
.B(n_49),
.Y(n_1026)
);

OAI21xp33_ASAP7_75t_L g1027 ( 
.A1(n_857),
.A2(n_51),
.B(n_52),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_793),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_793),
.Y(n_1029)
);

NAND2x1p5_ASAP7_75t_L g1030 ( 
.A(n_833),
.B(n_86),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_833),
.B(n_54),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_819),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_902),
.B(n_54),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_851),
.B(n_55),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_898),
.B(n_55),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_821),
.B(n_56),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_820),
.B(n_56),
.Y(n_1037)
);

CKINVDCx10_ASAP7_75t_R g1038 ( 
.A(n_821),
.Y(n_1038)
);

OAI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_863),
.A2(n_58),
.B(n_59),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_837),
.B(n_58),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_763),
.B(n_74),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_848),
.B(n_59),
.Y(n_1042)
);

OR2x6_ASAP7_75t_SL g1043 ( 
.A(n_831),
.B(n_62),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_797),
.A2(n_63),
.B(n_64),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_850),
.B(n_66),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_799),
.A2(n_68),
.B(n_72),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_852),
.B(n_68),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_864),
.B(n_73),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_875),
.B(n_811),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_800),
.A2(n_807),
.B(n_854),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_833),
.A2(n_756),
.B(n_774),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_L g1052 ( 
.A(n_855),
.B(n_911),
.C(n_880),
.Y(n_1052)
);

AOI21xp33_ASAP7_75t_L g1053 ( 
.A1(n_911),
.A2(n_766),
.B(n_773),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_802),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_784),
.B(n_903),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_795),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_903),
.A2(n_871),
.B(n_842),
.C(n_826),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_795),
.A2(n_853),
.B(n_869),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_878),
.A2(n_834),
.B(n_869),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_796),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_796),
.A2(n_815),
.B(n_853),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_827),
.A2(n_838),
.B1(n_776),
.B2(n_844),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_838),
.A2(n_825),
.B1(n_843),
.B2(n_834),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_798),
.A2(n_867),
.B(n_809),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_798),
.A2(n_867),
.B(n_809),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_825),
.A2(n_830),
.B(n_900),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_881),
.Y(n_1067)
);

BUFx2_ASAP7_75t_SL g1068 ( 
.A(n_790),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_838),
.A2(n_830),
.B1(n_900),
.B2(n_873),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_897),
.A2(n_873),
.B1(n_890),
.B2(n_862),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_765),
.B(n_889),
.C(n_892),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_897),
.A2(n_859),
.B(n_862),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_836),
.A2(n_891),
.B(n_859),
.C(n_868),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_SL g1074 ( 
.A1(n_778),
.A2(n_868),
.B1(n_876),
.B2(n_891),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_876),
.B(n_653),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_877),
.B(n_653),
.Y(n_1076)
);

O2A1O1Ixp5_ASAP7_75t_L g1077 ( 
.A1(n_824),
.A2(n_832),
.B(n_856),
.C(n_858),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_753),
.B(n_858),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_753),
.A2(n_755),
.B(n_805),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_801),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_L g1081 ( 
.A(n_833),
.B(n_606),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_753),
.B(n_858),
.Y(n_1082)
);

AND3x4_ASAP7_75t_L g1083 ( 
.A(n_923),
.B(n_1033),
.C(n_1008),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_913),
.B(n_1078),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_951),
.B(n_1079),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_982),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_963),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1079),
.B(n_914),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1075),
.B(n_1076),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_L g1090 ( 
.A(n_940),
.B(n_1052),
.C(n_939),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1050),
.B(n_928),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_1009),
.B(n_946),
.C(n_1003),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1050),
.B(n_968),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_953),
.B(n_1011),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_912),
.B(n_1068),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1081),
.A2(n_952),
.B(n_1002),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_922),
.A2(n_935),
.B(n_1024),
.C(n_1025),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1015),
.B(n_954),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1077),
.A2(n_930),
.B(n_925),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_941),
.B(n_919),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_926),
.A2(n_918),
.B(n_959),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_991),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_SL g1103 ( 
.A1(n_973),
.A2(n_1057),
.B(n_993),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_936),
.B(n_937),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_963),
.B(n_979),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_925),
.A2(n_932),
.B(n_948),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_945),
.A2(n_934),
.B(n_943),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_917),
.B(n_938),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_947),
.A2(n_967),
.B(n_961),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1058),
.A2(n_1065),
.B(n_1064),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_957),
.A2(n_1055),
.B(n_916),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1032),
.Y(n_1112)
);

OAI22x1_ASAP7_75t_L g1113 ( 
.A1(n_1026),
.A2(n_1041),
.B1(n_944),
.B2(n_1035),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1063),
.A2(n_1069),
.B(n_1053),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1061),
.A2(n_1066),
.B(n_1070),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1063),
.A2(n_1069),
.B(n_1062),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1070),
.A2(n_1072),
.B(n_1051),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1062),
.A2(n_966),
.B(n_1019),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_924),
.B(n_965),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1034),
.B(n_1067),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1033),
.B(n_1017),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_969),
.B(n_1049),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_963),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1049),
.B(n_1006),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_SL g1125 ( 
.A1(n_973),
.A2(n_993),
.B(n_1073),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_920),
.A2(n_927),
.B(n_964),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1056),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1016),
.B(n_1021),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1029),
.B(n_929),
.Y(n_1129)
);

OA22x2_ASAP7_75t_L g1130 ( 
.A1(n_999),
.A2(n_1010),
.B1(n_1005),
.B2(n_1039),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_950),
.B(n_1014),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1022),
.B(n_1028),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1060),
.Y(n_1133)
);

OR2x6_ASAP7_75t_L g1134 ( 
.A(n_912),
.B(n_976),
.Y(n_1134)
);

NAND2x1p5_ASAP7_75t_L g1135 ( 
.A(n_979),
.B(n_988),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_912),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_971),
.A2(n_985),
.B(n_921),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_985),
.A2(n_1013),
.B(n_994),
.Y(n_1138)
);

CKINVDCx8_ASAP7_75t_R g1139 ( 
.A(n_1038),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_L g1140 ( 
.A(n_980),
.B(n_958),
.C(n_1074),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1054),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1008),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1031),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_1036),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1031),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_981),
.B(n_987),
.Y(n_1146)
);

OAI21xp33_ASAP7_75t_L g1147 ( 
.A1(n_949),
.A2(n_1027),
.B(n_1037),
.Y(n_1147)
);

AND2x6_ASAP7_75t_L g1148 ( 
.A(n_979),
.B(n_1080),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1012),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_942),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_955),
.A2(n_977),
.B(n_962),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_942),
.Y(n_1152)
);

OR2x6_ASAP7_75t_L g1153 ( 
.A(n_988),
.B(n_1080),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_989),
.A2(n_915),
.A3(n_977),
.B(n_975),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1013),
.A2(n_995),
.B(n_1071),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_1043),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1018),
.A2(n_998),
.B(n_997),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1001),
.A2(n_1080),
.B(n_988),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1020),
.B(n_1040),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1023),
.A2(n_1030),
.B(n_996),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1042),
.A2(n_1048),
.B(n_1047),
.C(n_1045),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_991),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1001),
.A2(n_972),
.B(n_992),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_991),
.B(n_999),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1010),
.B(n_1007),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_972),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1030),
.A2(n_1007),
.B(n_1046),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1044),
.A2(n_984),
.B(n_986),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_990),
.A2(n_974),
.B(n_975),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_970),
.B(n_1004),
.Y(n_1170)
);

AND2x6_ASAP7_75t_L g1171 ( 
.A(n_1005),
.B(n_1000),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_960),
.A2(n_974),
.B(n_978),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_978),
.B(n_983),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_983),
.A2(n_951),
.B(n_1078),
.C(n_913),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_913),
.B(n_1078),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_989),
.A2(n_915),
.A3(n_858),
.B(n_1057),
.Y(n_1176)
);

OAI22x1_ASAP7_75t_L g1177 ( 
.A1(n_1003),
.A2(n_763),
.B1(n_1026),
.B2(n_1009),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1056),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_963),
.Y(n_1179)
);

INVx5_ASAP7_75t_L g1180 ( 
.A(n_963),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_L g1181 ( 
.A1(n_931),
.A2(n_1078),
.B(n_1082),
.C(n_913),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_913),
.B(n_1078),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_913),
.B(n_1078),
.Y(n_1183)
);

NOR2x1_ASAP7_75t_L g1184 ( 
.A(n_1052),
.B(n_790),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1079),
.A2(n_933),
.B(n_913),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_951),
.A2(n_913),
.B(n_1082),
.C(n_1078),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_965),
.Y(n_1187)
);

AOI21x1_ASAP7_75t_SL g1188 ( 
.A1(n_930),
.A2(n_1078),
.B(n_913),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1079),
.A2(n_933),
.B(n_913),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_989),
.A2(n_915),
.A3(n_858),
.B(n_1057),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1076),
.B(n_941),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_933),
.A2(n_761),
.B(n_1081),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_951),
.A2(n_913),
.B(n_1082),
.C(n_1078),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1032),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_913),
.B(n_1078),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_913),
.B(n_1078),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1076),
.B(n_941),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1079),
.A2(n_933),
.B(n_913),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1059),
.A2(n_933),
.B(n_956),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_963),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_913),
.B(n_1078),
.Y(n_1201)
);

OAI22x1_ASAP7_75t_L g1202 ( 
.A1(n_1003),
.A2(n_763),
.B1(n_1026),
.B2(n_1009),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_963),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1059),
.A2(n_933),
.B(n_956),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1059),
.A2(n_933),
.B(n_956),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_973),
.B(n_1049),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1079),
.A2(n_933),
.B(n_913),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1032),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_913),
.B(n_1078),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_933),
.A2(n_761),
.B(n_1081),
.Y(n_1210)
);

BUFx4_ASAP7_75t_SL g1211 ( 
.A(n_912),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1056),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_913),
.B(n_1078),
.Y(n_1213)
);

OR2x6_ASAP7_75t_L g1214 ( 
.A(n_912),
.B(n_770),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_963),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_913),
.B(n_1078),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_941),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_933),
.A2(n_761),
.B(n_1081),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_951),
.B(n_913),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_933),
.A2(n_761),
.B(n_1081),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1079),
.A2(n_933),
.B(n_913),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_963),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_933),
.A2(n_761),
.B(n_1081),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1059),
.A2(n_933),
.B(n_956),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_963),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1076),
.B(n_874),
.Y(n_1226)
);

O2A1O1Ixp5_ASAP7_75t_L g1227 ( 
.A1(n_931),
.A2(n_1078),
.B(n_1082),
.C(n_913),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_941),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1155),
.A2(n_1096),
.B(n_1138),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1107),
.A2(n_1189),
.B(n_1185),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1086),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1175),
.B(n_1182),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1185),
.A2(n_1198),
.B(n_1189),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1112),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1140),
.A2(n_1173),
.B1(n_1171),
.B2(n_1130),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1206),
.B(n_1166),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1206),
.B(n_1166),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1084),
.B(n_1183),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1191),
.B(n_1197),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1097),
.A2(n_1092),
.B(n_1174),
.C(n_1186),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1198),
.A2(n_1221),
.B(n_1207),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1100),
.B(n_1228),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1175),
.B(n_1182),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1166),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1195),
.B(n_1196),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1217),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1116),
.A2(n_1099),
.B(n_1114),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1228),
.B(n_1124),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1180),
.Y(n_1249)
);

BUFx12f_ASAP7_75t_L g1250 ( 
.A(n_1134),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1226),
.B(n_1090),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1195),
.A2(n_1216),
.B1(n_1213),
.B2(n_1196),
.Y(n_1252)
);

OR2x2_ASAP7_75t_SL g1253 ( 
.A(n_1165),
.B(n_1108),
.Y(n_1253)
);

NAND2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1180),
.B(n_1203),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1194),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1089),
.B(n_1201),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1150),
.B(n_1152),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1201),
.B(n_1209),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1187),
.Y(n_1259)
);

NOR2xp67_ASAP7_75t_SL g1260 ( 
.A(n_1139),
.B(n_1125),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1181),
.A2(n_1227),
.B(n_1193),
.Y(n_1261)
);

AOI221xp5_ASAP7_75t_L g1262 ( 
.A1(n_1219),
.A2(n_1165),
.B1(n_1202),
.B2(n_1177),
.C(n_1209),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1121),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1142),
.B(n_1122),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1171),
.A2(n_1130),
.B1(n_1113),
.B2(n_1083),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1136),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1213),
.A2(n_1216),
.B1(n_1103),
.B2(n_1164),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1203),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1208),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1161),
.A2(n_1144),
.B(n_1159),
.C(n_1146),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1119),
.B(n_1149),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1108),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1133),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1211),
.Y(n_1274)
);

OR2x2_ASAP7_75t_SL g1275 ( 
.A(n_1141),
.B(n_1089),
.Y(n_1275)
);

AOI21xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1156),
.A2(n_1120),
.B(n_1095),
.Y(n_1276)
);

INVx4_ASAP7_75t_L g1277 ( 
.A(n_1180),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1134),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1159),
.A2(n_1172),
.B(n_1147),
.C(n_1170),
.Y(n_1279)
);

NAND2x1p5_ASAP7_75t_L g1280 ( 
.A(n_1180),
.B(n_1215),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1215),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1095),
.Y(n_1282)
);

AO21x1_ASAP7_75t_L g1283 ( 
.A1(n_1118),
.A2(n_1085),
.B(n_1170),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1127),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1094),
.B(n_1093),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1143),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1171),
.A2(n_1145),
.B1(n_1184),
.B2(n_1093),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1087),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1192),
.A2(n_1218),
.B(n_1210),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1214),
.B(n_1095),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1214),
.B(n_1153),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1094),
.B(n_1098),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1098),
.B(n_1088),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1111),
.A2(n_1163),
.B(n_1169),
.C(n_1167),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1129),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1153),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1178),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1128),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1214),
.B(n_1153),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1220),
.A2(n_1223),
.B(n_1104),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1087),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1162),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1164),
.A2(n_1151),
.B(n_1106),
.C(n_1099),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1087),
.Y(n_1305)
);

NOR2x1_ASAP7_75t_L g1306 ( 
.A(n_1102),
.B(n_1225),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1091),
.B(n_1106),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1212),
.B(n_1102),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1123),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1171),
.A2(n_1137),
.B1(n_1128),
.B2(n_1131),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1123),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1123),
.B(n_1225),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1151),
.A2(n_1158),
.B(n_1126),
.C(n_1109),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1131),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1179),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1179),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1132),
.A2(n_1135),
.B1(n_1105),
.B2(n_1222),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1132),
.A2(n_1225),
.B1(n_1222),
.B2(n_1200),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1154),
.B(n_1190),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1179),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1200),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1200),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1115),
.A2(n_1110),
.B(n_1117),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1154),
.B(n_1190),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_SL g1325 ( 
.A1(n_1157),
.A2(n_1148),
.B1(n_1160),
.B2(n_1222),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1148),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1135),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1154),
.B(n_1176),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1188),
.A2(n_1190),
.B1(n_1176),
.B2(n_1148),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1168),
.B(n_1148),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1176),
.Y(n_1331)
);

INVx3_ASAP7_75t_SL g1332 ( 
.A(n_1199),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1204),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1205),
.A2(n_951),
.B1(n_923),
.B2(n_1092),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1101),
.B(n_1224),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1175),
.B(n_913),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1086),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1175),
.A2(n_913),
.B1(n_1082),
.B2(n_1078),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1092),
.A2(n_951),
.B1(n_923),
.B2(n_1173),
.Y(n_1339)
);

CKINVDCx8_ASAP7_75t_R g1340 ( 
.A(n_1086),
.Y(n_1340)
);

INVx3_ASAP7_75t_SL g1341 ( 
.A(n_1086),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1226),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1175),
.B(n_913),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1166),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_SL g1345 ( 
.A1(n_1111),
.A2(n_1165),
.B(n_1094),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1226),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1166),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1112),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1206),
.B(n_1166),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_SL g1350 ( 
.A(n_1150),
.Y(n_1350)
);

OR2x6_ASAP7_75t_L g1351 ( 
.A(n_1125),
.B(n_1103),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1166),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1133),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1166),
.Y(n_1354)
);

O2A1O1Ixp5_ASAP7_75t_L g1355 ( 
.A1(n_1097),
.A2(n_931),
.B(n_1078),
.C(n_913),
.Y(n_1355)
);

CKINVDCx6p67_ASAP7_75t_R g1356 ( 
.A(n_1150),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_R g1357 ( 
.A(n_1166),
.B(n_710),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1155),
.A2(n_1096),
.B(n_1138),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1175),
.B(n_913),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1206),
.B(n_1166),
.Y(n_1360)
);

BUFx4_ASAP7_75t_SL g1361 ( 
.A(n_1086),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1191),
.B(n_1197),
.Y(n_1362)
);

NAND2x1p5_ASAP7_75t_L g1363 ( 
.A(n_1180),
.B(n_963),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1112),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1166),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1219),
.A2(n_951),
.B(n_1078),
.C(n_913),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1086),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1086),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1133),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1092),
.A2(n_951),
.B1(n_923),
.B2(n_1173),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1175),
.B(n_913),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1175),
.B(n_913),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1133),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1191),
.B(n_1197),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1112),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1175),
.B(n_913),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1175),
.B(n_913),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1175),
.A2(n_913),
.B1(n_1082),
.B2(n_1078),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1133),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1155),
.A2(n_1096),
.B(n_1138),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1226),
.Y(n_1381)
);

INVx3_ASAP7_75t_SL g1382 ( 
.A(n_1086),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1155),
.A2(n_1096),
.B(n_1163),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1175),
.B(n_913),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1175),
.B(n_913),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1155),
.A2(n_1096),
.B(n_1138),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1191),
.B(n_1197),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1260),
.A2(n_1238),
.B1(n_1251),
.B2(n_1339),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1291),
.B(n_1290),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1351),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1239),
.B(n_1362),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1255),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1351),
.A2(n_1265),
.B1(n_1235),
.B2(n_1370),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1291),
.B(n_1300),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1267),
.A2(n_1262),
.B1(n_1287),
.B2(n_1387),
.Y(n_1395)
);

OR2x6_ASAP7_75t_L g1396 ( 
.A(n_1351),
.B(n_1240),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1346),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1269),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1232),
.B(n_1243),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1232),
.B(n_1243),
.Y(n_1400)
);

AO21x1_ASAP7_75t_L g1401 ( 
.A1(n_1329),
.A2(n_1304),
.B(n_1279),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1261),
.A2(n_1289),
.B(n_1301),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1245),
.A2(n_1258),
.B1(n_1384),
.B2(n_1371),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1381),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1229),
.A2(n_1380),
.B(n_1358),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1300),
.B(n_1282),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1257),
.Y(n_1407)
);

AO21x1_ASAP7_75t_SL g1408 ( 
.A1(n_1319),
.A2(n_1328),
.B(n_1324),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1348),
.Y(n_1409)
);

INVx8_ASAP7_75t_L g1410 ( 
.A(n_1300),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1245),
.A2(n_1258),
.B1(n_1385),
.B2(n_1377),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1364),
.Y(n_1412)
);

BUFx12f_ASAP7_75t_L g1413 ( 
.A(n_1321),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1336),
.A2(n_1371),
.B1(n_1385),
.B2(n_1384),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1259),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1336),
.A2(n_1359),
.B1(n_1377),
.B2(n_1376),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1262),
.A2(n_1267),
.B1(n_1374),
.B2(n_1338),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1326),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1338),
.A2(n_1378),
.B1(n_1252),
.B2(n_1343),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1375),
.Y(n_1420)
);

NAND2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1310),
.B(n_1247),
.Y(n_1421)
);

BUFx12f_ASAP7_75t_L g1422 ( 
.A(n_1250),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1246),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1256),
.B(n_1343),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1273),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1359),
.A2(n_1376),
.B1(n_1372),
.B2(n_1292),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1378),
.A2(n_1242),
.B1(n_1263),
.B2(n_1334),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1252),
.A2(n_1342),
.B1(n_1248),
.B2(n_1372),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1353),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1369),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1275),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1292),
.A2(n_1272),
.B1(n_1366),
.B2(n_1253),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1271),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1299),
.B(n_1295),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1285),
.B(n_1293),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1373),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1249),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1301),
.A2(n_1386),
.B(n_1380),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1379),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1261),
.A2(n_1323),
.B(n_1386),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1355),
.A2(n_1270),
.B(n_1383),
.C(n_1233),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1264),
.A2(n_1307),
.B1(n_1345),
.B2(n_1283),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1285),
.A2(n_1293),
.B1(n_1318),
.B2(n_1286),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1264),
.A2(n_1307),
.B1(n_1278),
.B2(n_1247),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1341),
.B(n_1382),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1249),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1303),
.Y(n_1447)
);

BUFx2_ASAP7_75t_SL g1448 ( 
.A(n_1337),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1284),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1308),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1361),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1309),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1340),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1298),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1296),
.B(n_1360),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1277),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1297),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1276),
.A2(n_1266),
.B1(n_1296),
.B2(n_1236),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1249),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1327),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1244),
.Y(n_1461)
);

OAI21xp33_ASAP7_75t_L g1462 ( 
.A1(n_1313),
.A2(n_1241),
.B(n_1230),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1244),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1237),
.A2(n_1349),
.B1(n_1350),
.B2(n_1331),
.Y(n_1464)
);

BUFx4f_ASAP7_75t_SL g1465 ( 
.A(n_1356),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1319),
.B(n_1328),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1317),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1306),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1326),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1349),
.A2(n_1350),
.B1(n_1274),
.B2(n_1347),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_1231),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1315),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1288),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1316),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1244),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1367),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1347),
.A2(n_1354),
.B1(n_1352),
.B2(n_1357),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1352),
.A2(n_1354),
.B1(n_1325),
.B2(n_1311),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1333),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1312),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1312),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1368),
.A2(n_1365),
.B1(n_1344),
.B2(n_1326),
.Y(n_1482)
);

CKINVDCx11_ASAP7_75t_R g1483 ( 
.A(n_1344),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1330),
.A2(n_1324),
.B(n_1363),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1344),
.Y(n_1485)
);

CKINVDCx11_ASAP7_75t_R g1486 ( 
.A(n_1365),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1302),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1302),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1322),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1365),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1320),
.A2(n_1268),
.B1(n_1281),
.B2(n_1305),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1294),
.A2(n_1335),
.B(n_1332),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1268),
.A2(n_1281),
.B1(n_1302),
.B2(n_1254),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1280),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1280),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1238),
.A2(n_1078),
.B1(n_1082),
.B2(n_913),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1346),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1234),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1238),
.B(n_1232),
.Y(n_1499)
);

INVx6_ASAP7_75t_L g1500 ( 
.A(n_1277),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1234),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1238),
.A2(n_1078),
.B1(n_1082),
.B2(n_913),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1234),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1351),
.A2(n_951),
.B1(n_1092),
.B2(n_923),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1257),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1275),
.Y(n_1506)
);

INVx4_ASAP7_75t_L g1507 ( 
.A(n_1249),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1275),
.Y(n_1508)
);

NAND2x1p5_ASAP7_75t_L g1509 ( 
.A(n_1310),
.B(n_1247),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1234),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1346),
.Y(n_1511)
);

BUFx4f_ASAP7_75t_SL g1512 ( 
.A(n_1337),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1234),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1351),
.A2(n_951),
.B1(n_1092),
.B2(n_923),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1337),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1238),
.A2(n_1078),
.B1(n_1082),
.B2(n_913),
.Y(n_1516)
);

NAND2x1p5_ASAP7_75t_L g1517 ( 
.A(n_1310),
.B(n_1247),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1234),
.Y(n_1518)
);

BUFx8_ASAP7_75t_L g1519 ( 
.A(n_1350),
.Y(n_1519)
);

INVx6_ASAP7_75t_L g1520 ( 
.A(n_1277),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1234),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1238),
.B(n_1232),
.Y(n_1522)
);

BUFx2_ASAP7_75t_SL g1523 ( 
.A(n_1277),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1314),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1238),
.A2(n_1078),
.B1(n_1082),
.B2(n_913),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1257),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1238),
.B(n_1232),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1361),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1466),
.B(n_1419),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1466),
.B(n_1421),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1396),
.B(n_1408),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1438),
.A2(n_1441),
.B(n_1401),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1450),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1453),
.Y(n_1534)
);

INVx4_ASAP7_75t_L g1535 ( 
.A(n_1410),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1410),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_SL g1537 ( 
.A1(n_1396),
.A2(n_1502),
.B(n_1496),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1438),
.A2(n_1401),
.B(n_1462),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1457),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1396),
.B(n_1408),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1421),
.B(n_1509),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1410),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1467),
.B(n_1417),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1457),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1391),
.B(n_1499),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1484),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1405),
.A2(n_1402),
.B(n_1516),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1525),
.A2(n_1527),
.B(n_1522),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1484),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1402),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1447),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1524),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1489),
.Y(n_1553)
);

NAND2x1p5_ASAP7_75t_L g1554 ( 
.A(n_1390),
.B(n_1492),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1406),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1433),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1440),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1453),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1406),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1392),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1421),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1509),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1424),
.B(n_1399),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1388),
.A2(n_1393),
.B1(n_1428),
.B2(n_1427),
.Y(n_1564)
);

INVxp67_ASAP7_75t_SL g1565 ( 
.A(n_1455),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1434),
.B(n_1442),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1434),
.B(n_1395),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1517),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1390),
.Y(n_1569)
);

CKINVDCx16_ASAP7_75t_R g1570 ( 
.A(n_1413),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1440),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1406),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1398),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1400),
.B(n_1414),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1431),
.B(n_1506),
.Y(n_1575)
);

INVx4_ASAP7_75t_SL g1576 ( 
.A(n_1500),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1394),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1409),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1416),
.B(n_1426),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1423),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1412),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1420),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1452),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1390),
.B(n_1479),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1498),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1501),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1444),
.B(n_1431),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1503),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1472),
.Y(n_1589)
);

NOR2xp67_ASAP7_75t_SL g1590 ( 
.A(n_1413),
.B(n_1523),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1506),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1515),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1394),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1492),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1394),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1508),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1492),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1510),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1508),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1513),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1389),
.B(n_1494),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1518),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1521),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1425),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1389),
.B(n_1435),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1432),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1397),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1389),
.B(n_1436),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1403),
.B(n_1411),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1443),
.B(n_1458),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1429),
.B(n_1430),
.Y(n_1611)
);

AO31x2_ASAP7_75t_L g1612 ( 
.A1(n_1478),
.A2(n_1460),
.A3(n_1439),
.B(n_1454),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1449),
.Y(n_1613)
);

OR2x6_ASAP7_75t_L g1614 ( 
.A(n_1523),
.B(n_1494),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1473),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1500),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1504),
.Y(n_1617)
);

BUFx3_ASAP7_75t_L g1618 ( 
.A(n_1407),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1480),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1514),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1481),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1474),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1456),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1468),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1497),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1594),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1530),
.B(n_1464),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1602),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1594),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1561),
.B(n_1505),
.Y(n_1630)
);

INVx4_ASAP7_75t_R g1631 ( 
.A(n_1618),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1530),
.B(n_1488),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1529),
.B(n_1511),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1554),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1529),
.B(n_1487),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1554),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1573),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1531),
.B(n_1477),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1540),
.B(n_1470),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1602),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1541),
.B(n_1415),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1579),
.B(n_1482),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1545),
.B(n_1471),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1574),
.B(n_1404),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1538),
.B(n_1469),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1609),
.B(n_1491),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1564),
.A2(n_1485),
.B1(n_1490),
.B2(n_1493),
.Y(n_1647)
);

BUFx2_ASAP7_75t_SL g1648 ( 
.A(n_1616),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1592),
.B(n_1476),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1609),
.B(n_1495),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1538),
.B(n_1418),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1557),
.B(n_1418),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1534),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1546),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1571),
.B(n_1532),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1565),
.B(n_1526),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1571),
.B(n_1418),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1571),
.B(n_1469),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1575),
.B(n_1526),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1575),
.B(n_1448),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1562),
.B(n_1437),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1554),
.Y(n_1662)
);

NAND3xp33_ASAP7_75t_SL g1663 ( 
.A(n_1617),
.B(n_1485),
.C(n_1490),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1625),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1569),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1606),
.B(n_1437),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_SL g1667 ( 
.A(n_1590),
.B(n_1519),
.Y(n_1667)
);

OR2x6_ASAP7_75t_L g1668 ( 
.A(n_1537),
.B(n_1500),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1553),
.B(n_1512),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1605),
.B(n_1459),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1566),
.B(n_1459),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1606),
.B(n_1446),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1569),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1566),
.B(n_1459),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1546),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1586),
.B(n_1588),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1532),
.B(n_1469),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1552),
.B(n_1446),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1539),
.Y(n_1679)
);

OAI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1617),
.A2(n_1465),
.B1(n_1507),
.B2(n_1422),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1563),
.B(n_1515),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1664),
.B(n_1533),
.Y(n_1682)
);

AND2x2_ASAP7_75t_SL g1683 ( 
.A(n_1667),
.B(n_1610),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1628),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1652),
.B(n_1562),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1664),
.B(n_1544),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1679),
.B(n_1556),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1679),
.B(n_1551),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1642),
.A2(n_1548),
.B1(n_1620),
.B2(n_1537),
.C(n_1589),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_L g1690 ( 
.A(n_1642),
.B(n_1620),
.C(n_1548),
.Y(n_1690)
);

OAI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1667),
.A2(n_1610),
.B1(n_1596),
.B2(n_1570),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1647),
.A2(n_1570),
.B1(n_1599),
.B2(n_1591),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1647),
.A2(n_1599),
.B1(n_1591),
.B2(n_1596),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1650),
.B(n_1641),
.Y(n_1694)
);

OAI221xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1644),
.A2(n_1547),
.B1(n_1567),
.B2(n_1587),
.C(n_1543),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1646),
.A2(n_1596),
.B1(n_1567),
.B2(n_1543),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1650),
.B(n_1641),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1656),
.B(n_1580),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1663),
.A2(n_1587),
.B1(n_1601),
.B2(n_1577),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1663),
.A2(n_1601),
.B1(n_1577),
.B2(n_1593),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1643),
.B(n_1607),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1656),
.B(n_1583),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1646),
.A2(n_1608),
.B1(n_1590),
.B2(n_1601),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1632),
.B(n_1622),
.Y(n_1704)
);

NOR3xp33_ASAP7_75t_L g1705 ( 
.A(n_1680),
.B(n_1535),
.C(n_1568),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1632),
.B(n_1604),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1644),
.A2(n_1555),
.B1(n_1572),
.B2(n_1559),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1657),
.B(n_1658),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1660),
.B(n_1558),
.Y(n_1709)
);

NAND3xp33_ASAP7_75t_L g1710 ( 
.A(n_1666),
.B(n_1625),
.C(n_1624),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1633),
.B(n_1604),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1633),
.B(n_1604),
.Y(n_1712)
);

OAI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1668),
.A2(n_1559),
.B1(n_1595),
.B2(n_1555),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1627),
.A2(n_1601),
.B1(n_1593),
.B2(n_1577),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1681),
.A2(n_1608),
.B1(n_1595),
.B2(n_1572),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1671),
.B(n_1560),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1658),
.B(n_1597),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1637),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1674),
.B(n_1578),
.Y(n_1719)
);

OAI21xp33_ASAP7_75t_SL g1720 ( 
.A1(n_1668),
.A2(n_1614),
.B(n_1600),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1678),
.B(n_1581),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_L g1722 ( 
.A(n_1666),
.B(n_1549),
.C(n_1624),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1680),
.B(n_1584),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1678),
.B(n_1581),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1670),
.B(n_1582),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1672),
.B(n_1549),
.C(n_1621),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1627),
.B(n_1665),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1660),
.A2(n_1559),
.B1(n_1593),
.B2(n_1536),
.Y(n_1728)
);

AOI221x1_ASAP7_75t_SL g1729 ( 
.A1(n_1672),
.A2(n_1603),
.B1(n_1600),
.B2(n_1613),
.C(n_1615),
.Y(n_1729)
);

NAND4xp25_ASAP7_75t_L g1730 ( 
.A(n_1635),
.B(n_1603),
.C(n_1613),
.D(n_1611),
.Y(n_1730)
);

OAI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1669),
.A2(n_1445),
.B1(n_1618),
.B2(n_1616),
.C(n_1542),
.Y(n_1731)
);

OAI221xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1668),
.A2(n_1614),
.B1(n_1451),
.B2(n_1621),
.C(n_1619),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1676),
.B(n_1582),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1673),
.B(n_1550),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1649),
.B(n_1422),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1661),
.B(n_1619),
.C(n_1623),
.Y(n_1736)
);

NAND4xp25_ASAP7_75t_L g1737 ( 
.A(n_1659),
.B(n_1611),
.C(n_1615),
.D(n_1598),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1676),
.B(n_1585),
.Y(n_1738)
);

OA211x2_ASAP7_75t_L g1739 ( 
.A1(n_1668),
.A2(n_1576),
.B(n_1519),
.C(n_1612),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1708),
.B(n_1655),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1708),
.B(n_1655),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1718),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1718),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1717),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1684),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1717),
.B(n_1727),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1710),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1729),
.B(n_1694),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1727),
.B(n_1645),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1734),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1706),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1685),
.B(n_1645),
.Y(n_1752)
);

INVx4_ASAP7_75t_L g1753 ( 
.A(n_1683),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1685),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1733),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1738),
.Y(n_1756)
);

NAND2x1p5_ASAP7_75t_L g1757 ( 
.A(n_1723),
.B(n_1634),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1720),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1683),
.B(n_1630),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1697),
.B(n_1626),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1721),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1711),
.B(n_1712),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1724),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1736),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1686),
.B(n_1626),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1682),
.B(n_1704),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1716),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1722),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1725),
.Y(n_1769)
);

NAND2xp33_ASAP7_75t_R g1770 ( 
.A(n_1709),
.B(n_1653),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1688),
.B(n_1629),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1723),
.B(n_1629),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1719),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1720),
.B(n_1651),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1726),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1702),
.B(n_1677),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1730),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1710),
.B(n_1628),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1687),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1749),
.B(n_1634),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1747),
.A2(n_1690),
.B(n_1695),
.C(n_1692),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1742),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1749),
.B(n_1740),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1749),
.B(n_1636),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1740),
.B(n_1636),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1742),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1743),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1772),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1740),
.B(n_1662),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1753),
.A2(n_1689),
.B1(n_1693),
.B2(n_1691),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1741),
.B(n_1662),
.Y(n_1791)
);

INVxp67_ASAP7_75t_SL g1792 ( 
.A(n_1768),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1741),
.B(n_1639),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1743),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1775),
.B(n_1698),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1741),
.B(n_1639),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1748),
.B(n_1696),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1766),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1775),
.B(n_1764),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1746),
.B(n_1673),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1743),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1746),
.B(n_1703),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1742),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1742),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1746),
.B(n_1703),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1779),
.B(n_1735),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1748),
.B(n_1701),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1760),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1760),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1772),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1775),
.B(n_1737),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1752),
.B(n_1677),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1760),
.Y(n_1813)
);

OAI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1747),
.A2(n_1731),
.B1(n_1715),
.B2(n_1699),
.C(n_1705),
.Y(n_1814)
);

NOR2xp67_ASAP7_75t_L g1815 ( 
.A(n_1753),
.B(n_1654),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1750),
.Y(n_1816)
);

OR2x2_ASAP7_75t_SL g1817 ( 
.A(n_1768),
.B(n_1659),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1750),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1764),
.A2(n_1715),
.B(n_1707),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1779),
.B(n_1640),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1750),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1777),
.B(n_1640),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1765),
.B(n_1654),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1771),
.Y(n_1824)
);

NOR2xp67_ASAP7_75t_L g1825 ( 
.A(n_1753),
.B(n_1675),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1798),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1807),
.B(n_1777),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1811),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1787),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1797),
.B(n_1777),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1787),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1794),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1792),
.B(n_1776),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1783),
.B(n_1757),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1794),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1783),
.B(n_1757),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1781),
.B(n_1753),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1799),
.B(n_1778),
.Y(n_1838)
);

INVx2_ASAP7_75t_SL g1839 ( 
.A(n_1788),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1801),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1811),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1806),
.B(n_1519),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1801),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1799),
.B(n_1778),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1782),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1817),
.B(n_1823),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1816),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1802),
.B(n_1757),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1816),
.Y(n_1849)
);

NOR2xp67_ASAP7_75t_L g1850 ( 
.A(n_1815),
.B(n_1753),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1822),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1820),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1818),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1802),
.B(n_1757),
.Y(n_1854)
);

NAND2x1_ASAP7_75t_L g1855 ( 
.A(n_1815),
.B(n_1758),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1818),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1805),
.B(n_1757),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1805),
.B(n_1758),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1795),
.B(n_1776),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1814),
.A2(n_1758),
.B1(n_1772),
.B2(n_1638),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1795),
.B(n_1776),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1817),
.B(n_1823),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1819),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1793),
.B(n_1755),
.Y(n_1864)
);

NAND2x1p5_ASAP7_75t_L g1865 ( 
.A(n_1825),
.B(n_1759),
.Y(n_1865)
);

AND2x2_ASAP7_75t_SL g1866 ( 
.A(n_1790),
.B(n_1700),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1824),
.B(n_1771),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1782),
.Y(n_1868)
);

OAI21xp33_ASAP7_75t_SL g1869 ( 
.A1(n_1825),
.A2(n_1759),
.B(n_1790),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1793),
.B(n_1774),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1796),
.B(n_1774),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1839),
.Y(n_1872)
);

NOR2x1_ASAP7_75t_L g1873 ( 
.A(n_1837),
.B(n_1788),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1838),
.B(n_1824),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_SL g1875 ( 
.A1(n_1863),
.A2(n_1770),
.B1(n_1528),
.B2(n_1788),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1838),
.B(n_1808),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1842),
.B(n_1528),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1839),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1845),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1826),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1829),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_SL g1882 ( 
.A(n_1869),
.B(n_1866),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1828),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_R g1884 ( 
.A(n_1866),
.B(n_1770),
.Y(n_1884)
);

INVx1_ASAP7_75t_SL g1885 ( 
.A(n_1841),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1829),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1831),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1845),
.Y(n_1888)
);

INVx2_ASAP7_75t_SL g1889 ( 
.A(n_1855),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1865),
.Y(n_1890)
);

AO21x2_ASAP7_75t_L g1891 ( 
.A1(n_1850),
.A2(n_1804),
.B(n_1803),
.Y(n_1891)
);

INVx1_ASAP7_75t_SL g1892 ( 
.A(n_1858),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1830),
.B(n_1766),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1827),
.B(n_1766),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1868),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1851),
.B(n_1796),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1844),
.B(n_1808),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1831),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1860),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1852),
.B(n_1833),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1834),
.B(n_1788),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1858),
.B(n_1844),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1846),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1832),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1848),
.B(n_1810),
.Y(n_1905)
);

INVx2_ASAP7_75t_SL g1906 ( 
.A(n_1855),
.Y(n_1906)
);

AOI21xp33_ASAP7_75t_L g1907 ( 
.A1(n_1846),
.A2(n_1813),
.B(n_1809),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1862),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1848),
.B(n_1810),
.Y(n_1909)
);

INVx2_ASAP7_75t_SL g1910 ( 
.A(n_1868),
.Y(n_1910)
);

OAI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1882),
.A2(n_1862),
.B1(n_1865),
.B2(n_1859),
.Y(n_1911)
);

AOI322xp5_ASAP7_75t_L g1912 ( 
.A1(n_1882),
.A2(n_1854),
.A3(n_1857),
.B1(n_1861),
.B2(n_1871),
.C1(n_1870),
.C2(n_1834),
.Y(n_1912)
);

NAND3xp33_ASAP7_75t_SL g1913 ( 
.A(n_1884),
.B(n_1865),
.C(n_1857),
.Y(n_1913)
);

OAI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1899),
.A2(n_1668),
.B1(n_1854),
.B2(n_1864),
.Y(n_1914)
);

AOI21xp33_ASAP7_75t_L g1915 ( 
.A1(n_1899),
.A2(n_1867),
.B(n_1835),
.Y(n_1915)
);

OAI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1880),
.A2(n_1668),
.B1(n_1810),
.B2(n_1867),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1883),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1885),
.B(n_1870),
.Y(n_1918)
);

INVx2_ASAP7_75t_SL g1919 ( 
.A(n_1910),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1881),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1903),
.B(n_1809),
.Y(n_1921)
);

A2O1A1Ixp33_ASAP7_75t_L g1922 ( 
.A1(n_1875),
.A2(n_1836),
.B(n_1810),
.C(n_1813),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1877),
.B(n_1836),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1889),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1881),
.Y(n_1925)
);

INVx1_ASAP7_75t_SL g1926 ( 
.A(n_1892),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1886),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1908),
.A2(n_1873),
.B1(n_1893),
.B2(n_1900),
.Y(n_1928)
);

OAI21xp5_ASAP7_75t_SL g1929 ( 
.A1(n_1873),
.A2(n_1907),
.B(n_1890),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1894),
.B(n_1871),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1902),
.B(n_1785),
.Y(n_1931)
);

OAI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1875),
.A2(n_1832),
.B1(n_1835),
.B2(n_1840),
.C(n_1843),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1890),
.A2(n_1739),
.B1(n_1772),
.B2(n_1638),
.Y(n_1933)
);

OAI32xp33_ASAP7_75t_L g1934 ( 
.A1(n_1889),
.A2(n_1856),
.A3(n_1849),
.B1(n_1847),
.B2(n_1853),
.Y(n_1934)
);

NOR4xp25_ASAP7_75t_L g1935 ( 
.A(n_1910),
.B(n_1843),
.C(n_1840),
.D(n_1847),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1896),
.B(n_1785),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1879),
.B(n_1789),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1886),
.Y(n_1938)
);

NOR2x1_ASAP7_75t_L g1939 ( 
.A(n_1891),
.B(n_1849),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1926),
.B(n_1879),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1939),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1917),
.B(n_1888),
.Y(n_1942)
);

INVx1_ASAP7_75t_SL g1943 ( 
.A(n_1918),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1921),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1923),
.B(n_1874),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1920),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1919),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1915),
.B(n_1888),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1936),
.B(n_1905),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1913),
.B(n_1874),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1924),
.B(n_1895),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1925),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1927),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1938),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1937),
.Y(n_1955)
);

NOR3xp33_ASAP7_75t_L g1956 ( 
.A(n_1911),
.B(n_1906),
.C(n_1895),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1934),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1931),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1911),
.A2(n_1906),
.B1(n_1909),
.B2(n_1905),
.Y(n_1959)
);

INVx1_ASAP7_75t_SL g1960 ( 
.A(n_1930),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1928),
.B(n_1872),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1935),
.B(n_1876),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1960),
.B(n_1932),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1962),
.A2(n_1929),
.B(n_1928),
.Y(n_1964)
);

AOI311xp33_ASAP7_75t_L g1965 ( 
.A1(n_1957),
.A2(n_1914),
.A3(n_1922),
.B(n_1916),
.C(n_1887),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_SL g1966 ( 
.A(n_1959),
.B(n_1914),
.Y(n_1966)
);

O2A1O1Ixp33_ASAP7_75t_L g1967 ( 
.A1(n_1962),
.A2(n_1916),
.B(n_1898),
.C(n_1904),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1961),
.A2(n_1878),
.B(n_1872),
.Y(n_1968)
);

O2A1O1Ixp33_ASAP7_75t_L g1969 ( 
.A1(n_1956),
.A2(n_1898),
.B(n_1887),
.C(n_1904),
.Y(n_1969)
);

OAI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1950),
.A2(n_1948),
.B1(n_1943),
.B2(n_1945),
.C(n_1912),
.Y(n_1970)
);

NAND2xp33_ASAP7_75t_R g1971 ( 
.A(n_1940),
.B(n_1876),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_SL g1972 ( 
.A1(n_1947),
.A2(n_1941),
.B1(n_1955),
.B2(n_1958),
.C(n_1944),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1949),
.B(n_1909),
.Y(n_1973)
);

OAI321xp33_ASAP7_75t_L g1974 ( 
.A1(n_1942),
.A2(n_1933),
.A3(n_1878),
.B1(n_1897),
.B2(n_1732),
.C(n_1728),
.Y(n_1974)
);

AOI221xp5_ASAP7_75t_L g1975 ( 
.A1(n_1941),
.A2(n_1891),
.B1(n_1897),
.B2(n_1901),
.C(n_1856),
.Y(n_1975)
);

A2O1A1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1944),
.A2(n_1901),
.B(n_1772),
.C(n_1774),
.Y(n_1976)
);

OAI211xp5_ASAP7_75t_L g1977 ( 
.A1(n_1964),
.A2(n_1951),
.B(n_1952),
.C(n_1954),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1970),
.B(n_1949),
.Y(n_1978)
);

NAND3xp33_ASAP7_75t_L g1979 ( 
.A(n_1972),
.B(n_1954),
.C(n_1952),
.Y(n_1979)
);

INVx1_ASAP7_75t_SL g1980 ( 
.A(n_1973),
.Y(n_1980)
);

OAI322xp33_ASAP7_75t_L g1981 ( 
.A1(n_1963),
.A2(n_1953),
.A3(n_1946),
.B1(n_1745),
.B2(n_1821),
.C1(n_1891),
.C2(n_1754),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1966),
.A2(n_1901),
.B1(n_1946),
.B2(n_1953),
.Y(n_1982)
);

NOR3xp33_ASAP7_75t_L g1983 ( 
.A(n_1967),
.B(n_1486),
.C(n_1483),
.Y(n_1983)
);

NOR2x1_ASAP7_75t_L g1984 ( 
.A(n_1969),
.B(n_1901),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1968),
.B(n_1789),
.Y(n_1985)
);

NAND5xp2_ASAP7_75t_L g1986 ( 
.A(n_1965),
.B(n_1714),
.C(n_1784),
.D(n_1780),
.E(n_1791),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1974),
.B(n_1976),
.Y(n_1987)
);

NOR3x1_ASAP7_75t_L g1988 ( 
.A(n_1971),
.B(n_1745),
.C(n_1821),
.Y(n_1988)
);

NAND2xp33_ASAP7_75t_L g1989 ( 
.A(n_1975),
.B(n_1780),
.Y(n_1989)
);

AOI211xp5_ASAP7_75t_L g1990 ( 
.A1(n_1986),
.A2(n_1713),
.B(n_1772),
.C(n_1784),
.Y(n_1990)
);

NOR3xp33_ASAP7_75t_L g1991 ( 
.A(n_1978),
.B(n_1486),
.C(n_1483),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1984),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1980),
.B(n_1791),
.Y(n_1993)
);

NAND4xp25_ASAP7_75t_L g1994 ( 
.A(n_1983),
.B(n_1739),
.C(n_1542),
.D(n_1536),
.Y(n_1994)
);

AOI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1982),
.A2(n_1979),
.B1(n_1989),
.B2(n_1987),
.C(n_1977),
.Y(n_1995)
);

OAI211xp5_ASAP7_75t_L g1996 ( 
.A1(n_1985),
.A2(n_1507),
.B(n_1463),
.C(n_1475),
.Y(n_1996)
);

NOR3xp33_ASAP7_75t_L g1997 ( 
.A(n_1981),
.B(n_1507),
.C(n_1475),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1993),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1995),
.A2(n_1988),
.B1(n_1804),
.B2(n_1803),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1991),
.A2(n_1786),
.B1(n_1812),
.B2(n_1800),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1992),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1997),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1990),
.B(n_1786),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1996),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_2001),
.B(n_1994),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1998),
.Y(n_2006)
);

NAND2x1p5_ASAP7_75t_L g2007 ( 
.A(n_2004),
.B(n_1463),
.Y(n_2007)
);

NOR2x1_ASAP7_75t_L g2008 ( 
.A(n_2002),
.B(n_1812),
.Y(n_2008)
);

AOI221xp5_ASAP7_75t_SL g2009 ( 
.A1(n_2003),
.A2(n_1754),
.B1(n_1761),
.B2(n_1763),
.C(n_1800),
.Y(n_2009)
);

INVxp33_ASAP7_75t_L g2010 ( 
.A(n_1999),
.Y(n_2010)
);

OAI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_2010),
.A2(n_2000),
.B(n_1763),
.Y(n_2011)
);

NOR2xp67_ASAP7_75t_L g2012 ( 
.A(n_2006),
.B(n_1461),
.Y(n_2012)
);

OAI211xp5_ASAP7_75t_L g2013 ( 
.A1(n_2005),
.A2(n_1763),
.B(n_1761),
.C(n_1771),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_2008),
.Y(n_2014)
);

AO22x1_ASAP7_75t_L g2015 ( 
.A1(n_2014),
.A2(n_2011),
.B1(n_2012),
.B2(n_2007),
.Y(n_2015)
);

NOR4xp25_ASAP7_75t_L g2016 ( 
.A(n_2015),
.B(n_2013),
.C(n_2009),
.D(n_1761),
.Y(n_2016)
);

AO22x2_ASAP7_75t_L g2017 ( 
.A1(n_2016),
.A2(n_1765),
.B1(n_1769),
.B2(n_1755),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2016),
.Y(n_2018)
);

OAI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_2018),
.A2(n_1461),
.B1(n_1769),
.B2(n_1765),
.Y(n_2019)
);

OAI21xp5_ASAP7_75t_SL g2020 ( 
.A1(n_2017),
.A2(n_1755),
.B(n_1756),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_2019),
.A2(n_1648),
.B1(n_1500),
.B2(n_1520),
.Y(n_2021)
);

OAI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_2020),
.A2(n_1762),
.B(n_1756),
.Y(n_2022)
);

NOR2x1_ASAP7_75t_L g2023 ( 
.A(n_2022),
.B(n_1648),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_2023),
.A2(n_2021),
.B1(n_1520),
.B2(n_1767),
.Y(n_2024)
);

OAI221xp5_ASAP7_75t_R g2025 ( 
.A1(n_2024),
.A2(n_1520),
.B1(n_1576),
.B2(n_1631),
.C(n_1744),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_2025),
.A2(n_1520),
.B1(n_1751),
.B2(n_1773),
.Y(n_2026)
);


endmodule