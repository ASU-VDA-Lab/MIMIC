module fake_jpeg_1708_n_534 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_534);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_55),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_56),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_21),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_57),
.A2(n_15),
.B1(n_31),
.B2(n_29),
.Y(n_125)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_69),
.B(n_40),
.Y(n_99)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_17),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_93),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_33),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_87),
.Y(n_97)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_95),
.Y(n_109)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_28),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_99),
.B(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_20),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_102),
.B(n_125),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_45),
.A2(n_44),
.B1(n_40),
.B2(n_35),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_113),
.A2(n_117),
.B1(n_126),
.B2(n_152),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_43),
.B1(n_17),
.B2(n_39),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_SL g122 ( 
.A(n_79),
.Y(n_122)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_54),
.A2(n_40),
.B1(n_43),
.B2(n_39),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_40),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_131),
.B(n_139),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_52),
.B(n_24),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_46),
.A2(n_64),
.B1(n_48),
.B2(n_80),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_76),
.Y(n_194)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_106),
.A2(n_29),
.B1(n_27),
.B2(n_31),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_162),
.A2(n_41),
.B1(n_131),
.B2(n_115),
.Y(n_221)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_47),
.B1(n_62),
.B2(n_55),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_165),
.A2(n_177),
.B1(n_142),
.B2(n_121),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_170),
.Y(n_219)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx4_ASAP7_75t_SL g218 ( 
.A(n_167),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_168),
.Y(n_214)
);

AOI32xp33_ASAP7_75t_L g169 ( 
.A1(n_106),
.A2(n_49),
.A3(n_81),
.B1(n_20),
.B2(n_38),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_194),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_97),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_174),
.Y(n_224)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_192),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_125),
.A2(n_38),
.B1(n_24),
.B2(n_37),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_111),
.B(n_103),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_196),
.Y(n_230)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_98),
.B(n_68),
.C(n_56),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_195),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g233 ( 
.A(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_113),
.A2(n_75),
.B1(n_61),
.B2(n_37),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_188),
.A2(n_197),
.B1(n_201),
.B2(n_135),
.Y(n_215)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_191),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_108),
.B(n_19),
.C(n_27),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_125),
.B(n_151),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_126),
.A2(n_15),
.B1(n_81),
.B2(n_33),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

INVx4_ASAP7_75t_SL g200 ( 
.A(n_105),
.Y(n_200)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_40),
.B1(n_15),
.B2(n_78),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_118),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_203),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_100),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_140),
.B(n_0),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_206),
.Y(n_234)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_114),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_128),
.B(n_0),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_215),
.A2(n_203),
.B1(n_168),
.B2(n_184),
.Y(n_269)
);

OAI21xp33_ASAP7_75t_SL g259 ( 
.A1(n_221),
.A2(n_168),
.B(n_187),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_165),
.B1(n_180),
.B2(n_185),
.Y(n_246)
);

AO22x1_ASAP7_75t_SL g227 ( 
.A1(n_160),
.A2(n_129),
.B1(n_112),
.B2(n_149),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_239),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_174),
.Y(n_235)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_166),
.B(n_134),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_238),
.B(n_230),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_242),
.A2(n_239),
.B(n_224),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_246),
.A2(n_267),
.B1(n_214),
.B2(n_218),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_248),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_199),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_256),
.C(n_260),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_210),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_251),
.Y(n_284)
);

AO21x2_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_196),
.B(n_178),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_254),
.B1(n_265),
.B2(n_268),
.Y(n_273)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_223),
.A2(n_172),
.B1(n_199),
.B2(n_173),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_216),
.C(n_226),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_257),
.Y(n_297)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_264),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_181),
.C(n_190),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_206),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_163),
.C(n_164),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_192),
.C(n_229),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_204),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_211),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_219),
.A2(n_172),
.B1(n_195),
.B2(n_193),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_211),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_270),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_215),
.A2(n_110),
.B1(n_146),
.B2(n_138),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_220),
.A2(n_170),
.B1(n_202),
.B2(n_198),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_269),
.A2(n_208),
.B(n_176),
.Y(n_302)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_212),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_274),
.B(n_200),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_212),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_286),
.Y(n_306)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_252),
.A2(n_227),
.B1(n_213),
.B2(n_229),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_285),
.A2(n_252),
.B1(n_267),
.B2(n_260),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_213),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_295),
.C(n_279),
.Y(n_307)
);

AOI32xp33_ASAP7_75t_L g290 ( 
.A1(n_247),
.A2(n_235),
.A3(n_227),
.B1(n_222),
.B2(n_179),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_242),
.B(n_237),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_292),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_241),
.B(n_207),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_250),
.A2(n_182),
.B1(n_218),
.B2(n_157),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_299),
.B1(n_233),
.B2(n_232),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_249),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_205),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_207),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_SL g296 ( 
.A(n_265),
.B(n_161),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_101),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_250),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_301),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_245),
.A2(n_218),
.B1(n_237),
.B2(n_217),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_254),
.B(n_214),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_270),
.B1(n_266),
.B2(n_264),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g349 ( 
.A(n_303),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_298),
.A2(n_252),
.B1(n_246),
.B2(n_245),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_309),
.B1(n_310),
.B2(n_319),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_307),
.B(n_312),
.C(n_328),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_308),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_301),
.A2(n_286),
.B1(n_282),
.B2(n_283),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_301),
.A2(n_253),
.B1(n_248),
.B2(n_257),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_262),
.C(n_271),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_321),
.C(n_300),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_209),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_314),
.B(n_318),
.Y(n_365)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_271),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_327),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_209),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_278),
.A2(n_258),
.B1(n_243),
.B2(n_240),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_275),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_320),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_287),
.B(n_240),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_273),
.A2(n_233),
.B1(n_157),
.B2(n_138),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_273),
.A2(n_233),
.B1(n_232),
.B2(n_167),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_285),
.A2(n_208),
.B1(n_175),
.B2(n_186),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_275),
.Y(n_325)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_278),
.B(n_101),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_289),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_334),
.Y(n_356)
);

AOI21xp33_ASAP7_75t_L g362 ( 
.A1(n_331),
.A2(n_191),
.B(n_200),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_189),
.C(n_171),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_332),
.B(n_333),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_274),
.B(n_291),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_191),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_272),
.A2(n_127),
.B1(n_116),
.B2(n_149),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_335),
.A2(n_277),
.B1(n_280),
.B2(n_297),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_367),
.Y(n_374)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_340),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_305),
.A2(n_272),
.B(n_302),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_341),
.A2(n_343),
.B(n_347),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_305),
.A2(n_272),
.B(n_292),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_326),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_345),
.B(n_358),
.Y(n_377)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_329),
.A2(n_272),
.B(n_290),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_309),
.Y(n_348)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_348),
.Y(n_378)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_306),
.Y(n_350)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_311),
.A2(n_299),
.B(n_280),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_353),
.B(n_362),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_311),
.A2(n_297),
.B(n_288),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_315),
.A2(n_288),
.B1(n_276),
.B2(n_277),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_354),
.A2(n_361),
.B1(n_346),
.B2(n_330),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_304),
.Y(n_357)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_306),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_310),
.Y(n_360)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_315),
.A2(n_276),
.B1(n_281),
.B2(n_142),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_308),
.A2(n_320),
.B1(n_323),
.B2(n_322),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_363),
.A2(n_366),
.B1(n_335),
.B2(n_328),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_324),
.A2(n_281),
.B1(n_136),
.B2(n_127),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_316),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_351),
.B(n_312),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_397),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_307),
.C(n_317),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_384),
.C(n_386),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_355),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_371),
.B(n_390),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_373),
.A2(n_380),
.B1(n_382),
.B2(n_385),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_354),
.Y(n_376)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_365),
.B(n_332),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_379),
.B(n_392),
.Y(n_408)
);

OAI22x1_ASAP7_75t_L g382 ( 
.A1(n_360),
.A2(n_333),
.B1(n_327),
.B2(n_281),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_334),
.C(n_143),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_367),
.A2(n_281),
.B1(n_143),
.B2(n_136),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_121),
.C(n_191),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_154),
.C(n_88),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_396),
.C(n_337),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_355),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_365),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_391),
.B(n_361),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_281),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_393),
.Y(n_419)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_338),
.Y(n_395)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_395),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_359),
.B(n_154),
.C(n_95),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_343),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_395),
.Y(n_398)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_398),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_374),
.A2(n_388),
.B(n_372),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_399),
.B(n_416),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_353),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_400),
.B(n_401),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_358),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_383),
.A2(n_363),
.B1(n_336),
.B2(n_357),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_402),
.A2(n_159),
.B1(n_33),
.B2(n_41),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_378),
.B(n_350),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_404),
.B(n_412),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_341),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_411),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_397),
.B(n_356),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_409),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_347),
.Y(n_409)
);

FAx1_ASAP7_75t_SL g412 ( 
.A(n_369),
.B(n_345),
.CI(n_357),
.CON(n_412),
.SN(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_352),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_413),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_337),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_414),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_338),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_417),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_388),
.A2(n_340),
.B(n_349),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_362),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_377),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_422),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_342),
.C(n_344),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_421),
.B(n_375),
.C(n_380),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_342),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_425),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_429),
.B(n_440),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_414),
.A2(n_377),
.B(n_383),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_436),
.B(n_417),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_394),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_431),
.B(n_432),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_375),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_406),
.A2(n_368),
.B(n_381),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_381),
.Y(n_439)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_439),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_368),
.C(n_373),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_415),
.A2(n_387),
.B(n_366),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_441),
.A2(n_12),
.B(n_11),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_385),
.C(n_33),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_442),
.B(n_449),
.Y(n_466)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_398),
.Y(n_443)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_443),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_405),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_444),
.B(n_413),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_402),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_445),
.B(n_414),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_446),
.A2(n_33),
.B1(n_42),
.B2(n_3),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_411),
.B(n_33),
.C(n_159),
.Y(n_449)
);

MAJx2_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_403),
.C(n_407),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_467),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_435),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_421),
.C(n_403),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_454),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_414),
.C(n_422),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_457),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_412),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_456),
.A2(n_459),
.B1(n_462),
.B2(n_463),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_420),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_448),
.A2(n_445),
.B1(n_447),
.B2(n_436),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_464),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_14),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_13),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_430),
.A2(n_13),
.B(n_12),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_465),
.A2(n_469),
.B1(n_468),
.B2(n_438),
.Y(n_479)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_12),
.C(n_11),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_468),
.B(n_441),
.Y(n_472)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_472),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_470),
.B(n_440),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_474),
.B(n_475),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_458),
.B(n_429),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_460),
.B(n_459),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_464),
.Y(n_488)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_479),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_452),
.C(n_437),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_433),
.C(n_455),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_SL g481 ( 
.A1(n_456),
.A2(n_438),
.B1(n_446),
.B2(n_428),
.Y(n_481)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_481),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_435),
.Y(n_482)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_482),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_483),
.B(n_486),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_463),
.B(n_442),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_484),
.A2(n_487),
.B(n_466),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_433),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_449),
.Y(n_487)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_488),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_490),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_492),
.B(n_497),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_473),
.A2(n_465),
.B(n_467),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_493),
.A2(n_496),
.B(n_3),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_462),
.Y(n_495)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_495),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_483),
.A2(n_36),
.B(n_2),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_0),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_36),
.Y(n_498)
);

AOI21x1_ASAP7_75t_L g505 ( 
.A1(n_498),
.A2(n_499),
.B(n_471),
.Y(n_505)
);

AO21x1_ASAP7_75t_L g499 ( 
.A1(n_481),
.A2(n_36),
.B(n_2),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_486),
.C(n_477),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_512),
.Y(n_520)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_505),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_500),
.A2(n_472),
.B(n_2),
.Y(n_508)
);

AOI31xp33_ASAP7_75t_L g517 ( 
.A1(n_508),
.A2(n_499),
.A3(n_498),
.B(n_6),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_489),
.B(n_0),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_511),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_4),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_489),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_5),
.C(n_6),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_494),
.B(n_4),
.Y(n_514)
);

NOR3xp33_ASAP7_75t_L g518 ( 
.A(n_514),
.B(n_4),
.C(n_5),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_507),
.A2(n_501),
.B(n_491),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_515),
.A2(n_522),
.B(n_506),
.Y(n_523)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_517),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_518),
.B(n_519),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_503),
.A2(n_5),
.B(n_6),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_524),
.C(n_525),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_516),
.A2(n_509),
.B(n_504),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_520),
.A2(n_513),
.B(n_521),
.Y(n_525)
);

OAI321xp33_ASAP7_75t_L g528 ( 
.A1(n_526),
.A2(n_517),
.A3(n_510),
.B1(n_7),
.B2(n_8),
.C(n_10),
.Y(n_528)
);

O2A1O1Ixp33_ASAP7_75t_SL g532 ( 
.A1(n_528),
.A2(n_529),
.B(n_5),
.C(n_7),
.Y(n_532)
);

OAI321xp33_ASAP7_75t_L g529 ( 
.A1(n_527),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_10),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g531 ( 
.A(n_530),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_532),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_8),
.Y(n_534)
);


endmodule