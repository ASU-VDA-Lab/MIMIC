module real_jpeg_5307_n_6 (n_46, n_5, n_4, n_43, n_0, n_1, n_47, n_2, n_45, n_44, n_3, n_6);

input n_46;
input n_5;
input n_4;
input n_43;
input n_0;
input n_1;
input n_47;
input n_2;
input n_45;
input n_44;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_40;
wire n_39;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_0),
.B(n_36),
.Y(n_38)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_1),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_4),
.B(n_11),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_18),
.B1(n_40),
.B2(n_41),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_16),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_21),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_23),
.B(n_39),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_22),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_35),
.B(n_38),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B(n_34),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_33),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_43),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_44),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_45),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_46),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_47),
.Y(n_37)
);


endmodule