module fake_aes_3262_n_517 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_517);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_517;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_84;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx5_ASAP7_75t_L g76 ( .A(n_9), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_18), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_44), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_60), .Y(n_79) );
BUFx10_ASAP7_75t_L g80 ( .A(n_48), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_70), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_4), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_75), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_62), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_25), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_14), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_69), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_41), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_13), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_39), .Y(n_90) );
BUFx2_ASAP7_75t_L g91 ( .A(n_56), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_59), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_13), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_49), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_15), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_4), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_28), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_17), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_14), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_11), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_55), .Y(n_101) );
CKINVDCx14_ASAP7_75t_R g102 ( .A(n_9), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_5), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_50), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_61), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_21), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_51), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_68), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_7), .Y(n_109) );
AND2x2_ASAP7_75t_L g110 ( .A(n_91), .B(n_0), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_76), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_91), .B(n_0), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_88), .Y(n_113) );
OAI22xp5_ASAP7_75t_SL g114 ( .A1(n_86), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_76), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_102), .B(n_1), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_76), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_76), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_76), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_86), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_80), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
BUFx12f_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_82), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_103), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_76), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_82), .B(n_6), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_76), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_78), .B(n_6), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_78), .B(n_7), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_119), .Y(n_133) );
INVx4_ASAP7_75t_L g134 ( .A(n_115), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_115), .B(n_81), .Y(n_135) );
INVx6_ASAP7_75t_L g136 ( .A(n_113), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_115), .B(n_103), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_126), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_115), .B(n_97), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_122), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_111), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_110), .B(n_109), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_126), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_122), .B(n_77), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_119), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_113), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
NAND2x1p5_ASAP7_75t_L g148 ( .A(n_110), .B(n_83), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_124), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_113), .Y(n_150) );
OR2x6_ASAP7_75t_L g151 ( .A(n_114), .B(n_109), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_113), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_122), .B(n_98), .Y(n_154) );
OAI21xp33_ASAP7_75t_SL g155 ( .A1(n_131), .A2(n_95), .B(n_89), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_119), .Y(n_156) );
INVx1_ASAP7_75t_SL g157 ( .A(n_124), .Y(n_157) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_110), .B(n_85), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_138), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_138), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_134), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_158), .B(n_112), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_149), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_134), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_134), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_143), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_149), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_142), .B(n_112), .Y(n_170) );
INVx5_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_158), .B(n_117), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_148), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_158), .B(n_122), .Y(n_176) );
BUFx2_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_140), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
INVxp67_ASAP7_75t_SL g180 ( .A(n_148), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_142), .B(n_125), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_140), .B(n_117), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_144), .B(n_125), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_141), .B(n_131), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_141), .B(n_117), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
CKINVDCx8_ASAP7_75t_R g190 ( .A(n_151), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_145), .Y(n_191) );
OR2x6_ASAP7_75t_L g192 ( .A(n_151), .B(n_114), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_184), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_174), .B(n_154), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_180), .A2(n_151), .B1(n_90), .B2(n_128), .Y(n_196) );
NOR2xp33_ASAP7_75t_SL g197 ( .A(n_174), .B(n_90), .Y(n_197) );
INVx8_ASAP7_75t_L g198 ( .A(n_171), .Y(n_198) );
BUFx2_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_162), .A2(n_151), .B1(n_128), .B2(n_137), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_171), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_171), .B(n_124), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_186), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_184), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_171), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_171), .Y(n_206) );
OAI22xp33_ASAP7_75t_L g207 ( .A1(n_192), .A2(n_151), .B1(n_98), .B2(n_139), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_171), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_170), .B(n_155), .Y(n_209) );
BUFx12f_ASAP7_75t_L g210 ( .A(n_165), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_184), .Y(n_211) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_177), .B(n_85), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_170), .B(n_135), .Y(n_213) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_168), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_177), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_170), .B(n_155), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_161), .A2(n_152), .B(n_147), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_173), .A2(n_121), .B1(n_130), .B2(n_132), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_173), .B(n_170), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_191), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_167), .Y(n_221) );
OAI22xp33_ASAP7_75t_L g222 ( .A1(n_192), .A2(n_93), .B1(n_100), .B2(n_99), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_159), .B(n_121), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_167), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_160), .B(n_147), .Y(n_225) );
OR2x6_ASAP7_75t_L g226 ( .A(n_198), .B(n_183), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_198), .Y(n_227) );
AOI222xp33_ASAP7_75t_L g228 ( .A1(n_223), .A2(n_181), .B1(n_162), .B2(n_163), .C1(n_176), .C2(n_175), .Y(n_228) );
OAI22xp33_ASAP7_75t_L g229 ( .A1(n_197), .A2(n_192), .B1(n_190), .B2(n_169), .Y(n_229) );
HB1xp67_ASAP7_75t_SL g230 ( .A(n_212), .Y(n_230) );
OR2x2_ASAP7_75t_L g231 ( .A(n_196), .B(n_176), .Y(n_231) );
INVxp67_ASAP7_75t_L g232 ( .A(n_197), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_224), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_224), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_196), .A2(n_192), .B1(n_183), .B2(n_161), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_203), .B(n_185), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_203), .A2(n_212), .B1(n_183), .B2(n_200), .Y(n_237) );
BUFx3_ASAP7_75t_L g238 ( .A(n_198), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_208), .B(n_167), .Y(n_239) );
OAI22xp33_ASAP7_75t_L g240 ( .A1(n_199), .A2(n_192), .B1(n_190), .B2(n_185), .Y(n_240) );
AND2x6_ASAP7_75t_L g241 ( .A(n_220), .B(n_167), .Y(n_241) );
BUFx12f_ASAP7_75t_L g242 ( .A(n_210), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_198), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_210), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_219), .B(n_187), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_198), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_207), .B(n_199), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_210), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_212), .B(n_208), .Y(n_249) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_217), .A2(n_189), .B(n_188), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_215), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_214), .Y(n_252) );
OAI221xp5_ASAP7_75t_L g253 ( .A1(n_235), .A2(n_200), .B1(n_218), .B2(n_209), .C(n_216), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_237), .A2(n_209), .B(n_193), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_240), .A2(n_222), .B1(n_219), .B2(n_195), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_250), .A2(n_186), .B(n_187), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_233), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_251), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_233), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_236), .B(n_215), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_236), .B(n_195), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_251), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
OAI22xp33_ASAP7_75t_L g264 ( .A1(n_229), .A2(n_218), .B1(n_213), .B2(n_225), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_247), .A2(n_195), .B1(n_220), .B2(n_221), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_228), .A2(n_195), .B1(n_220), .B2(n_221), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_228), .A2(n_220), .B1(n_221), .B2(n_202), .Y(n_267) );
INVx5_ASAP7_75t_SL g268 ( .A(n_226), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_245), .B(n_193), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_234), .Y(n_270) );
OAI222xp33_ASAP7_75t_L g271 ( .A1(n_230), .A2(n_96), .B1(n_108), .B2(n_87), .C1(n_92), .C2(n_94), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_231), .A2(n_208), .B1(n_204), .B2(n_194), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_252), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_227), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_253), .A2(n_232), .B(n_249), .C(n_266), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_264), .A2(n_231), .B1(n_226), .B2(n_246), .Y(n_276) );
INVx4_ASAP7_75t_L g277 ( .A(n_274), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_253), .A2(n_226), .B1(n_246), .B2(n_243), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_257), .Y(n_279) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_256), .B(n_113), .C(n_108), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_260), .B(n_238), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_260), .B(n_226), .Y(n_282) );
OAI31xp33_ASAP7_75t_L g283 ( .A1(n_271), .A2(n_238), .A3(n_239), .B(n_87), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_257), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_255), .A2(n_226), .B1(n_243), .B2(n_227), .Y(n_285) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_259), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_274), .B(n_243), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_274), .Y(n_288) );
OAI221xp5_ASAP7_75t_L g289 ( .A1(n_265), .A2(n_205), .B1(n_201), .B2(n_193), .C(n_206), .Y(n_289) );
OAI33xp33_ASAP7_75t_L g290 ( .A1(n_259), .A2(n_101), .A3(n_104), .B1(n_105), .B2(n_106), .B3(n_79), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_261), .B(n_227), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_261), .B(n_227), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_273), .A2(n_227), .B1(n_242), .B2(n_239), .Y(n_293) );
OAI21xp33_ASAP7_75t_L g294 ( .A1(n_267), .A2(n_256), .B(n_254), .Y(n_294) );
BUFx12f_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_269), .B(n_239), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_277), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_283), .A2(n_285), .B1(n_276), .B2(n_278), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_284), .B(n_263), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_284), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_277), .B(n_274), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_279), .B(n_286), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_279), .B(n_258), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_292), .B(n_263), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_295), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
NAND4xp25_ASAP7_75t_L g307 ( .A(n_275), .B(n_84), .C(n_107), .D(n_79), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_288), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_294), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_294), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_280), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_280), .Y(n_312) );
AOI22xp33_ASAP7_75t_SL g313 ( .A1(n_282), .A2(n_268), .B1(n_262), .B2(n_242), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_277), .Y(n_314) );
AOI222xp33_ASAP7_75t_L g315 ( .A1(n_290), .A2(n_268), .B1(n_269), .B2(n_270), .C1(n_248), .C2(n_244), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_276), .B(n_270), .Y(n_317) );
OAI21xp5_ASAP7_75t_L g318 ( .A1(n_289), .A2(n_272), .B(n_250), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_292), .B(n_268), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_287), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_282), .B(n_268), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_296), .B(n_268), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_287), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
OR2x2_ASAP7_75t_SL g325 ( .A(n_291), .B(n_84), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_287), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_293), .Y(n_327) );
OAI322xp33_ASAP7_75t_L g328 ( .A1(n_303), .A2(n_113), .A3(n_129), .B1(n_127), .B2(n_123), .C1(n_118), .C2(n_116), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_300), .B(n_113), .Y(n_329) );
CKINVDCx6p67_ASAP7_75t_R g330 ( .A(n_314), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_303), .B(n_8), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_300), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_300), .B(n_88), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_324), .B(n_8), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_299), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_314), .Y(n_336) );
OAI31xp33_ASAP7_75t_L g337 ( .A1(n_307), .A2(n_239), .A3(n_205), .B(n_201), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_302), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_297), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_313), .A2(n_206), .B1(n_201), .B2(n_208), .Y(n_340) );
NAND4xp25_ASAP7_75t_L g341 ( .A(n_298), .B(n_118), .C(n_123), .D(n_129), .Y(n_341) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_302), .B(n_206), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_299), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_308), .Y(n_344) );
NAND4xp25_ASAP7_75t_L g345 ( .A(n_315), .B(n_120), .C(n_150), .D(n_12), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_304), .B(n_10), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_306), .B(n_10), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_308), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_306), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_323), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_327), .B(n_11), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_323), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_327), .B(n_12), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_320), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_306), .B(n_15), .Y(n_355) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_297), .B(n_120), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_317), .B(n_16), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_320), .B(n_16), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_316), .Y(n_360) );
AOI31xp33_ASAP7_75t_L g361 ( .A1(n_313), .A2(n_17), .A3(n_120), .B(n_211), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_326), .Y(n_362) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_297), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_317), .B(n_150), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_305), .B(n_241), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_319), .B(n_241), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_345), .A2(n_307), .B1(n_322), .B2(n_319), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_335), .B(n_309), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_338), .B(n_311), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_335), .B(n_309), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_344), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_338), .B(n_312), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_344), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_330), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_330), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_336), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_360), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_361), .A2(n_316), .B1(n_297), .B2(n_325), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_348), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_343), .B(n_312), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_343), .B(n_346), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_350), .Y(n_384) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_356), .B(n_301), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_332), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_346), .B(n_310), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_350), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_352), .B(n_310), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_354), .B(n_321), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_354), .B(n_321), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_334), .B(n_316), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_352), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_347), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_332), .Y(n_396) );
AO21x2_ASAP7_75t_L g397 ( .A1(n_329), .A2(n_318), .B(n_301), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_367), .B(n_318), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_342), .B(n_301), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_363), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_367), .B(n_301), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_359), .B(n_322), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_359), .B(n_146), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_339), .Y(n_404) );
OAI21x1_ASAP7_75t_SL g405 ( .A1(n_339), .A2(n_325), .B(n_211), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_337), .A2(n_241), .B(n_204), .Y(n_406) );
AND2x4_ASAP7_75t_SL g407 ( .A(n_358), .B(n_204), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_349), .B(n_146), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_362), .B(n_146), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_342), .A2(n_194), .B1(n_224), .B2(n_191), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_362), .B(n_146), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g412 ( .A1(n_356), .A2(n_241), .B(n_194), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_331), .B(n_19), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_331), .B(n_20), .Y(n_414) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_333), .Y(n_415) );
AOI211x1_ASAP7_75t_SL g416 ( .A1(n_351), .A2(n_22), .B(n_23), .C(n_24), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_357), .B(n_26), .Y(n_417) );
INVxp33_ASAP7_75t_L g418 ( .A(n_355), .Y(n_418) );
AOI322xp5_ASAP7_75t_L g419 ( .A1(n_380), .A2(n_342), .A3(n_353), .B1(n_355), .B2(n_358), .C1(n_333), .C2(n_349), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g420 ( .A(n_392), .B(n_357), .C(n_364), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_387), .B(n_329), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_368), .A2(n_365), .B1(n_366), .B2(n_364), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_377), .A2(n_341), .B1(n_328), .B2(n_340), .C(n_194), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_372), .Y(n_424) );
INVx3_ASAP7_75t_SL g425 ( .A(n_376), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_383), .B(n_27), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_374), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_402), .B(n_29), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_400), .B(n_30), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_379), .B(n_31), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_390), .B(n_32), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_378), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_384), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_369), .B(n_136), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_400), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_369), .B(n_136), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_375), .B(n_33), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_388), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_386), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_371), .B(n_136), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_393), .Y(n_442) );
AOI221xp5_ASAP7_75t_SL g443 ( .A1(n_399), .A2(n_34), .B1(n_35), .B2(n_36), .C(n_37), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_382), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_386), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_371), .B(n_136), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_370), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_390), .B(n_391), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_373), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_396), .Y(n_450) );
NOR2x1_ASAP7_75t_L g451 ( .A(n_406), .B(n_191), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_391), .Y(n_452) );
AND2x4_ASAP7_75t_SL g453 ( .A(n_404), .B(n_191), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_401), .B(n_38), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_407), .Y(n_455) );
NOR3xp33_ASAP7_75t_L g456 ( .A(n_417), .B(n_189), .C(n_188), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_405), .B(n_188), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_398), .Y(n_458) );
XOR2xp5_ASAP7_75t_L g459 ( .A(n_418), .B(n_40), .Y(n_459) );
XNOR2x1_ASAP7_75t_L g460 ( .A(n_410), .B(n_42), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_389), .Y(n_461) );
NOR2xp33_ASAP7_75t_R g462 ( .A(n_394), .B(n_43), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_413), .A2(n_189), .B(n_182), .C(n_179), .Y(n_463) );
OR2x6_ASAP7_75t_L g464 ( .A(n_399), .B(n_45), .Y(n_464) );
AOI221x1_ASAP7_75t_L g465 ( .A1(n_414), .A2(n_46), .B1(n_47), .B2(n_52), .C(n_53), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_395), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_415), .Y(n_467) );
OA22x2_ASAP7_75t_L g468 ( .A1(n_407), .A2(n_54), .B1(n_57), .B2(n_58), .Y(n_468) );
AO22x1_ASAP7_75t_L g469 ( .A1(n_418), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_398), .B(n_66), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_412), .B(n_145), .C(n_179), .Y(n_471) );
NAND2xp33_ASAP7_75t_SL g472 ( .A(n_397), .B(n_67), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_408), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_408), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_397), .B(n_71), .Y(n_475) );
XOR2x2_ASAP7_75t_L g476 ( .A(n_385), .B(n_72), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_397), .B(n_73), .Y(n_477) );
AOI211xp5_ASAP7_75t_L g478 ( .A1(n_403), .A2(n_74), .B(n_178), .C(n_172), .Y(n_478) );
OA21x2_ASAP7_75t_SL g479 ( .A1(n_385), .A2(n_416), .B(n_411), .Y(n_479) );
OAI21xp33_ASAP7_75t_SL g480 ( .A1(n_411), .A2(n_178), .B(n_166), .Y(n_480) );
XOR2x2_ASAP7_75t_L g481 ( .A(n_403), .B(n_152), .Y(n_481) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_409), .B(n_145), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_425), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_458), .A2(n_422), .B1(n_420), .B2(n_444), .Y(n_484) );
AOI31xp33_ASAP7_75t_L g485 ( .A1(n_438), .A2(n_443), .A3(n_459), .B(n_436), .Y(n_485) );
INVx6_ASAP7_75t_L g486 ( .A(n_464), .Y(n_486) );
AOI22x1_ASAP7_75t_L g487 ( .A1(n_436), .A2(n_429), .B1(n_467), .B2(n_455), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_480), .A2(n_476), .B(n_419), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_480), .A2(n_438), .B1(n_464), .B2(n_449), .C(n_447), .Y(n_489) );
AOI211xp5_ASAP7_75t_L g490 ( .A1(n_469), .A2(n_462), .B(n_426), .C(n_472), .Y(n_490) );
O2A1O1Ixp5_ASAP7_75t_L g491 ( .A1(n_461), .A2(n_457), .B(n_466), .C(n_429), .Y(n_491) );
AOI21xp33_ASAP7_75t_L g492 ( .A1(n_426), .A2(n_475), .B(n_477), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_468), .A2(n_457), .B(n_481), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_452), .A2(n_421), .B1(n_431), .B2(n_427), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_424), .A2(n_433), .B1(n_432), .B2(n_442), .C(n_439), .Y(n_495) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_434), .A2(n_448), .B1(n_473), .B2(n_474), .C(n_423), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_491), .A2(n_453), .B(n_451), .C(n_478), .Y(n_497) );
NOR4xp25_ASAP7_75t_L g498 ( .A(n_483), .B(n_463), .C(n_430), .D(n_470), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_485), .A2(n_453), .B(n_482), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g500 ( .A1(n_488), .A2(n_460), .B1(n_471), .B2(n_479), .C(n_437), .Y(n_500) );
NAND4xp25_ASAP7_75t_SL g501 ( .A(n_493), .B(n_479), .C(n_465), .D(n_428), .Y(n_501) );
OAI211xp5_ASAP7_75t_SL g502 ( .A1(n_496), .A2(n_446), .B(n_435), .C(n_441), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_487), .A2(n_454), .B(n_456), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_495), .A2(n_440), .B1(n_450), .B2(n_445), .C(n_454), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_500), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_501), .A2(n_490), .B(n_489), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_502), .A2(n_486), .B1(n_492), .B2(n_484), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_503), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g509 ( .A1(n_506), .A2(n_498), .B1(n_499), .B2(n_486), .C(n_504), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_505), .A2(n_497), .B1(n_494), .B2(n_456), .C(n_445), .Y(n_510) );
OAI221xp5_ASAP7_75t_L g511 ( .A1(n_509), .A2(n_507), .B1(n_508), .B2(n_133), .C(n_156), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_510), .A2(n_133), .B1(n_156), .B2(n_164), .C(n_182), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_511), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_512), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_513), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_515), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_516), .A2(n_513), .B(n_514), .Y(n_517) );
endmodule