module fake_jpeg_4102_n_245 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_245);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_0),
.B(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_7),
.CON(n_33),
.SN(n_33)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_27),
.B1(n_15),
.B2(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_14),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_27),
.B1(n_18),
.B2(n_20),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_52),
.B1(n_23),
.B2(n_17),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_18),
.B1(n_27),
.B2(n_14),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_17),
.B1(n_16),
.B2(n_25),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_54),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_30),
.A2(n_15),
.B1(n_17),
.B2(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_31),
.B(n_26),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_60),
.B(n_65),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_28),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_29),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_71),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_38),
.C(n_36),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_43),
.B(n_46),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_68),
.Y(n_85)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_80),
.B1(n_57),
.B2(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_79),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_20),
.B1(n_19),
.B2(n_28),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_16),
.B1(n_57),
.B2(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_19),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_42),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_90),
.B1(n_96),
.B2(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_59),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_89),
.A2(n_95),
.B1(n_53),
.B2(n_62),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_50),
.B1(n_57),
.B2(n_58),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_75),
.B1(n_72),
.B2(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_103),
.Y(n_117)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_100),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_53),
.B1(n_49),
.B2(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_81),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_66),
.B(n_65),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_63),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_83),
.C(n_85),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_76),
.B(n_61),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_29),
.B(n_25),
.Y(n_145)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_121),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_69),
.B1(n_76),
.B2(n_61),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_122),
.B1(n_95),
.B2(n_103),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_64),
.B1(n_53),
.B2(n_62),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_49),
.B1(n_29),
.B2(n_25),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_65),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_132),
.B1(n_143),
.B2(n_107),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_130),
.B(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_93),
.B1(n_82),
.B2(n_84),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_135),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_136),
.C(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_90),
.C(n_102),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_142),
.B(n_144),
.Y(n_161)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_66),
.B(n_99),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_91),
.B1(n_100),
.B2(n_49),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_0),
.B(n_1),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_105),
.B(n_138),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_118),
.B1(n_126),
.B2(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_107),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_151),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_121),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_158),
.B1(n_94),
.B2(n_108),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_105),
.Y(n_151)
);

NOR2xp67_ASAP7_75t_R g152 ( 
.A(n_140),
.B(n_125),
.Y(n_152)
);

OAI322xp33_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_11),
.A3(n_13),
.B1(n_12),
.B2(n_4),
.C1(n_6),
.C2(n_8),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_114),
.C(n_118),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_163),
.B1(n_169),
.B2(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_114),
.B(n_111),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_0),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_144),
.B(n_130),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_134),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_184),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_174),
.C(n_179),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_159),
.A2(n_128),
.B1(n_94),
.B2(n_108),
.Y(n_172)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_38),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_176),
.B(n_180),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_162),
.C(n_6),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_186),
.B(n_169),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_108),
.C(n_56),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_162),
.C(n_160),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_56),
.B1(n_70),
.B2(n_3),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_155),
.B1(n_157),
.B2(n_164),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_56),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_187),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_179),
.B1(n_168),
.B2(n_173),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_153),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_201),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_166),
.Y(n_193)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_193),
.B(n_182),
.CI(n_180),
.CON(n_206),
.SN(n_206)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_149),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_196),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_153),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_202),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_161),
.B(n_165),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_151),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_208),
.C(n_200),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_189),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_204),
.B(n_212),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_193),
.B(n_195),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_214),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_171),
.C(n_178),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_174),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_211),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_184),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_158),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_197),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_222),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_224),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_198),
.B(n_191),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_206),
.A2(n_197),
.B1(n_191),
.B2(n_163),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_209),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_213),
.A2(n_163),
.B(n_9),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_221),
.Y(n_226)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_205),
.B(n_210),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_228),
.A2(n_229),
.B(n_230),
.Y(n_235)
);

AOI21x1_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_8),
.B(n_13),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_0),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_231),
.B(n_1),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_220),
.B(n_70),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_233),
.B(n_9),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_4),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_8),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_236),
.A2(n_235),
.B(n_225),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_238),
.B(n_239),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_9),
.C(n_12),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_1),
.B(n_3),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_241),
.C(n_3),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_3),
.Y(n_245)
);


endmodule