module fake_netlist_6_4381_n_1189 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_342, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1189);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1189;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_465;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1079;
wire n_362;
wire n_828;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_419;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_703;
wire n_578;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_595;
wire n_627;
wire n_524;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_1164;
wire n_509;
wire n_575;
wire n_368;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_840;
wire n_392;
wire n_568;
wire n_442;
wire n_874;
wire n_480;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_898;
wire n_617;
wire n_698;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_1095;
wire n_573;
wire n_769;
wire n_639;
wire n_963;
wire n_676;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_718;
wire n_517;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_742;
wire n_532;
wire n_535;
wire n_691;
wire n_901;
wire n_544;
wire n_372;
wire n_468;
wire n_1078;
wire n_504;
wire n_923;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_948;
wire n_522;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_1119;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_516;
wire n_1163;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_838;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_1176;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_638;
wire n_1181;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_1183;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_1054;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_492;
wire n_972;
wire n_699;
wire n_551;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_624;
wire n_451;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_796;
wire n_686;
wire n_1041;
wire n_757;
wire n_719;
wire n_594;
wire n_565;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_855;
wire n_513;
wire n_776;
wire n_645;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_608;
wire n_811;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_1110;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_993;
wire n_409;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_1155;
wire n_756;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_1051;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_1125;
wire n_652;
wire n_553;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_1111;
wire n_511;
wire n_715;
wire n_467;
wire n_359;
wire n_973;
wire n_1053;
wire n_416;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_1167;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_651;
wire n_404;
wire n_1153;
wire n_439;
wire n_518;
wire n_679;
wire n_1069;
wire n_1185;
wire n_612;
wire n_453;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_588;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_1175;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_743;
wire n_766;
wire n_816;
wire n_1157;
wire n_430;
wire n_527;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_825;
wire n_636;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_1124;
wire n_784;
wire n_434;
wire n_515;
wire n_983;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_1077;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_1082;
wire n_1154;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_736;
wire n_613;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_827;
wire n_531;
wire n_1001;
wire n_361;
wire n_663;
wire n_508;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_891;
wire n_1150;
wire n_410;
wire n_398;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_214),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_20),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_153),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_21),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_34),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_134),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_4),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_6),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_4),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_238),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_270),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_11),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_45),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_251),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_159),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_236),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_78),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_321),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_164),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_151),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_149),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_209),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_347),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_312),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_182),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_115),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_146),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_327),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_277),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_125),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_127),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_63),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_147),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_76),
.Y(n_385)
);

INVxp33_ASAP7_75t_SL g386 ( 
.A(n_160),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_93),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_328),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_53),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_323),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_272),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_118),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_73),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_203),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_124),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_6),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g397 ( 
.A(n_217),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_46),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_305),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_204),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_216),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_56),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_2),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_319),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_190),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_260),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_36),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_111),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_79),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_324),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_222),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_104),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_110),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_144),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_310),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_280),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_171),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_213),
.Y(n_419)
);

INVxp33_ASAP7_75t_SL g420 ( 
.A(n_334),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_228),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_218),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_212),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_175),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_35),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_307),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_48),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_220),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_136),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_139),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_193),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_52),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_84),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_18),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_259),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_14),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_83),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_1),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_223),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_131),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_287),
.B(n_186),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_257),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_51),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_126),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_261),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_234),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_62),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_121),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_227),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_254),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_174),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_140),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_316),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g454 ( 
.A(n_313),
.B(n_142),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_264),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_90),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_335),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_263),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_1),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_99),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_348),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_304),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_101),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_47),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_308),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_243),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_293),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_198),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_177),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_66),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_332),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_345),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_100),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_183),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_86),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_75),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_26),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_290),
.Y(n_478)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_43),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_31),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_267),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_114),
.Y(n_482)
);

BUFx2_ASAP7_75t_SL g483 ( 
.A(n_232),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_128),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_245),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_137),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_94),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_30),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_279),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_130),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_70),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_338),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_342),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_339),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_306),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_8),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_150),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_33),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_258),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_19),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_276),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_141),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_275),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_314),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_15),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_71),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_81),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_239),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_237),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_246),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_69),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_133),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_303),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_162),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_207),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_22),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_318),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_61),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_325),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_288),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_309),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_269),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_252),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_315),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_300),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_291),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_336),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_113),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_341),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_49),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_120),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_286),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_157),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_15),
.Y(n_534)
);

INVxp33_ASAP7_75t_L g535 ( 
.A(n_337),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_322),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_311),
.Y(n_537)
);

INVxp33_ASAP7_75t_L g538 ( 
.A(n_156),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_196),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_230),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_271),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_16),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_3),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_283),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_255),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_7),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_122),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_158),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_329),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_72),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_330),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_67),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_168),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_29),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_2),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_221),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_16),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_195),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_10),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_320),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_74),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_265),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_59),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_343),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_38),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_64),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_331),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_28),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_192),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_184),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_0),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_14),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_197),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_152),
.Y(n_574)
);

BUFx5_ASAP7_75t_L g575 ( 
.A(n_266),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_248),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_229),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_262),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_422),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_356),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_529),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_358),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_349),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_403),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_361),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_430),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_469),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_575),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_351),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_474),
.B(n_0),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_436),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_438),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_505),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_575),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_575),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_427),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_534),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_397),
.B(n_3),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_401),
.B(n_5),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_575),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_401),
.B(n_17),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_430),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_543),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_575),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_396),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_559),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_353),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_492),
.B(n_503),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_496),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_479),
.B(n_9),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_429),
.Y(n_611)
);

CKINVDCx16_ASAP7_75t_R g612 ( 
.A(n_377),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_571),
.Y(n_613)
);

OA21x2_ASAP7_75t_L g614 ( 
.A1(n_350),
.A2(n_9),
.B(n_10),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_501),
.B(n_11),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_430),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_406),
.B(n_12),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_572),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_352),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_409),
.B(n_12),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_379),
.B(n_13),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_354),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_500),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_555),
.B(n_13),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_500),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_357),
.B(n_23),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_359),
.B(n_24),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_360),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_445),
.B(n_25),
.Y(n_629)
);

AND2x2_ASAP7_75t_SL g630 ( 
.A(n_392),
.B(n_27),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_500),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_450),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_457),
.B(n_32),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_362),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_459),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_363),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_364),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_366),
.B(n_37),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_458),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_365),
.Y(n_640)
);

CKINVDCx16_ASAP7_75t_R g641 ( 
.A(n_407),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_466),
.B(n_39),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_L g643 ( 
.A(n_542),
.B(n_40),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_412),
.B(n_41),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_471),
.B(n_42),
.Y(n_645)
);

OR2x6_ASAP7_75t_L g646 ( 
.A(n_483),
.B(n_44),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_367),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_476),
.A2(n_498),
.B1(n_538),
.B2(n_535),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_368),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_369),
.B(n_50),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_370),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_371),
.B(n_54),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_433),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_SL g654 ( 
.A1(n_355),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_373),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_375),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_376),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_380),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_381),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_372),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_481),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_518),
.B(n_60),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_383),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_SL g664 ( 
.A1(n_546),
.A2(n_65),
.B1(n_68),
.B2(n_77),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_386),
.B(n_80),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_384),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_528),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_385),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_387),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_389),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_378),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_390),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_393),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_561),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_395),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_399),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_400),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_404),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_405),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_410),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_411),
.B(n_82),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_382),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_414),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_388),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_415),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_416),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_418),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_574),
.B(n_85),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_419),
.Y(n_689)
);

NOR2x1_ASAP7_75t_L g690 ( 
.A(n_454),
.B(n_87),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_421),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_602),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_579),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_602),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_589),
.B(n_423),
.Y(n_695)
);

INVx8_ASAP7_75t_L g696 ( 
.A(n_607),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_584),
.B(n_557),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_640),
.Y(n_698)
);

INVxp33_ASAP7_75t_L g699 ( 
.A(n_635),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_623),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_660),
.B(n_424),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_671),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_612),
.B(n_398),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_641),
.B(n_420),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_616),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_581),
.B(n_452),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_605),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_616),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_682),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_684),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_632),
.Y(n_711)
);

AND2x2_ASAP7_75t_SL g712 ( 
.A(n_630),
.B(n_644),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_632),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_625),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_631),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_605),
.B(n_428),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_583),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_636),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_596),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_587),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_639),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_610),
.B(n_523),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_639),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_586),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_637),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_647),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_648),
.A2(n_470),
.B1(n_502),
.B2(n_460),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_608),
.B(n_495),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_656),
.Y(n_729)
);

OAI22xp33_ASAP7_75t_L g730 ( 
.A1(n_609),
.A2(n_570),
.B1(n_441),
.B2(n_544),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_661),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_645),
.B(n_485),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_580),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_661),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_590),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_582),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_667),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_SL g738 ( 
.A1(n_654),
.A2(n_539),
.B1(n_570),
.B2(n_432),
.Y(n_738)
);

AND2x6_ASAP7_75t_L g739 ( 
.A(n_690),
.B(n_431),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_611),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_667),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_653),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_659),
.B(n_391),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_674),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_674),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_591),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_621),
.B(n_434),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_601),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_598),
.A2(n_408),
.B1(n_446),
.B2(n_374),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_666),
.B(n_394),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_689),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_624),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_689),
.Y(n_753)
);

OR2x4_ASAP7_75t_L g754 ( 
.A(n_697),
.B(n_592),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_752),
.B(n_706),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_752),
.B(n_722),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_721),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_736),
.A2(n_599),
.B(n_615),
.C(n_617),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_723),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_744),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_748),
.A2(n_601),
.B(n_626),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_720),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_709),
.B(n_646),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_722),
.B(n_627),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_743),
.B(n_638),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_745),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_750),
.B(n_650),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_753),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_712),
.A2(n_601),
.B1(n_614),
.B2(n_652),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_737),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_732),
.B(n_665),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_695),
.B(n_646),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_735),
.B(n_669),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_728),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_701),
.B(n_681),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_730),
.A2(n_614),
.B1(n_620),
.B2(n_619),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_735),
.B(n_749),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_710),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_700),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_719),
.Y(n_780)
);

BUFx8_ASAP7_75t_L g781 ( 
.A(n_693),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_714),
.A2(n_643),
.B(n_633),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_696),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_711),
.Y(n_784)
);

AND2x6_ASAP7_75t_SL g785 ( 
.A(n_716),
.B(n_597),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_747),
.B(n_622),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_699),
.B(n_727),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_707),
.A2(n_664),
.B1(n_642),
.B2(n_662),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_746),
.Y(n_789)
);

BUFx5_ASAP7_75t_L g790 ( 
.A(n_739),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_698),
.B(n_628),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_737),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_739),
.B(n_634),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_741),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_739),
.B(n_657),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_724),
.B(n_718),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_725),
.B(n_663),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_702),
.B(n_670),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_741),
.B(n_402),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_713),
.B(n_672),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_726),
.B(n_675),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_703),
.B(n_678),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_731),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_734),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_708),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_775),
.B(n_696),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_776),
.A2(n_688),
.B1(n_629),
.B2(n_738),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_800),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_756),
.A2(n_679),
.B(n_687),
.C(n_680),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_794),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_765),
.A2(n_482),
.B(n_464),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_780),
.Y(n_812)
);

INVx5_ASAP7_75t_L g813 ( 
.A(n_794),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_783),
.Y(n_814)
);

BUFx12f_ASAP7_75t_L g815 ( 
.A(n_785),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_767),
.A2(n_573),
.B(n_553),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_805),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_779),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_772),
.B(n_704),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_805),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_789),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_774),
.B(n_733),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_755),
.B(n_716),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_759),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_769),
.B(n_578),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_802),
.B(n_717),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_758),
.A2(n_437),
.B(n_439),
.C(n_435),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_784),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_791),
.B(n_729),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_766),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_798),
.B(n_440),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_777),
.A2(n_691),
.B(n_677),
.C(n_685),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_773),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_754),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_757),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_778),
.B(n_740),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_781),
.Y(n_837)
);

O2A1O1Ixp5_ASAP7_75t_SL g838 ( 
.A1(n_771),
.A2(n_651),
.B(n_655),
.C(n_649),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_768),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_762),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_764),
.A2(n_761),
.B1(n_788),
.B2(n_786),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_796),
.A2(n_594),
.B(n_588),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_763),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_763),
.B(n_751),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_790),
.B(n_413),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_790),
.B(n_442),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_770),
.B(n_742),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_782),
.A2(n_600),
.B(n_595),
.Y(n_848)
);

BUFx12f_ASAP7_75t_L g849 ( 
.A(n_799),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_760),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_848),
.A2(n_795),
.B(n_793),
.Y(n_851)
);

AO21x2_ASAP7_75t_L g852 ( 
.A1(n_846),
.A2(n_825),
.B(n_841),
.Y(n_852)
);

OR2x6_ASAP7_75t_L g853 ( 
.A(n_837),
.B(n_787),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_807),
.A2(n_790),
.B1(n_447),
.B2(n_448),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_838),
.A2(n_804),
.B(n_803),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_818),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_821),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_812),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_819),
.A2(n_790),
.B1(n_831),
.B2(n_833),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_808),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_811),
.A2(n_449),
.B1(n_451),
.B2(n_444),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_834),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_842),
.A2(n_801),
.B(n_797),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_829),
.B(n_453),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_830),
.Y(n_865)
);

OAI21x1_ASAP7_75t_L g866 ( 
.A1(n_845),
.A2(n_792),
.B(n_461),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_850),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_824),
.Y(n_868)
);

BUFx2_ASAP7_75t_R g869 ( 
.A(n_840),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_828),
.B(n_708),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_835),
.Y(n_871)
);

AOI21xp33_ASAP7_75t_L g872 ( 
.A1(n_826),
.A2(n_823),
.B(n_806),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_843),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_843),
.B(n_736),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_817),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_810),
.Y(n_876)
);

BUFx10_ASAP7_75t_L g877 ( 
.A(n_836),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_839),
.B(n_692),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_SL g879 ( 
.A1(n_849),
.A2(n_847),
.B1(n_814),
.B2(n_828),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_810),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_820),
.Y(n_881)
);

OAI21x1_ASAP7_75t_L g882 ( 
.A1(n_816),
.A2(n_462),
.B(n_455),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_877),
.B(n_844),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_853),
.B(n_815),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_877),
.B(n_822),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_872),
.B(n_832),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_871),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_852),
.A2(n_827),
.B(n_813),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_873),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_871),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_851),
.A2(n_809),
.B(n_465),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_853),
.B(n_603),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_860),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_869),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_864),
.B(n_683),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_SL g896 ( 
.A1(n_874),
.A2(n_813),
.B1(n_425),
.B2(n_426),
.Y(n_896)
);

AOI221xp5_ASAP7_75t_L g897 ( 
.A1(n_854),
.A2(n_677),
.B1(n_691),
.B2(n_606),
.C(n_618),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_R g898 ( 
.A(n_858),
.B(n_876),
.Y(n_898)
);

AOI221xp5_ASAP7_75t_L g899 ( 
.A1(n_874),
.A2(n_593),
.B1(n_585),
.B2(n_582),
.C(n_613),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_852),
.A2(n_813),
.B(n_467),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_856),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_859),
.A2(n_468),
.B(n_463),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_881),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_862),
.B(n_876),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_880),
.B(n_694),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_856),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_863),
.A2(n_857),
.B(n_867),
.Y(n_907)
);

AOI222xp33_ASAP7_75t_L g908 ( 
.A1(n_857),
.A2(n_585),
.B1(n_613),
.B2(n_686),
.C1(n_676),
.C2(n_673),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_865),
.B(n_658),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_865),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_SL g911 ( 
.A1(n_868),
.A2(n_443),
.B1(n_456),
.B2(n_417),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_861),
.A2(n_473),
.B1(n_477),
.B2(n_475),
.Y(n_912)
);

OAI211xp5_ASAP7_75t_L g913 ( 
.A1(n_879),
.A2(n_478),
.B(n_484),
.C(n_480),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_887),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_889),
.B(n_875),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_890),
.Y(n_916)
);

NAND3xp33_ASAP7_75t_L g917 ( 
.A(n_886),
.B(n_878),
.C(n_489),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_893),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_907),
.A2(n_882),
.B(n_855),
.Y(n_919)
);

OAI22xp33_ASAP7_75t_L g920 ( 
.A1(n_892),
.A2(n_870),
.B1(n_486),
.B2(n_488),
.Y(n_920)
);

BUFx2_ASAP7_75t_R g921 ( 
.A(n_909),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_904),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_901),
.B(n_866),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_885),
.B(n_472),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_892),
.B(n_883),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_903),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_906),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_910),
.A2(n_487),
.B1(n_491),
.B2(n_517),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_903),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_895),
.B(n_493),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_896),
.B(n_705),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_908),
.Y(n_932)
);

INVxp67_ASAP7_75t_SL g933 ( 
.A(n_905),
.Y(n_933)
);

OR2x6_ASAP7_75t_L g934 ( 
.A(n_884),
.B(n_705),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_891),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_902),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_897),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_898),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_894),
.B(n_715),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_884),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_913),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_899),
.B(n_715),
.Y(n_942)
);

OAI211xp5_ASAP7_75t_SL g943 ( 
.A1(n_912),
.A2(n_668),
.B(n_533),
.C(n_577),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_911),
.B(n_490),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_888),
.B(n_494),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_900),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_889),
.B(n_497),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_887),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_889),
.B(n_510),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_887),
.B(n_499),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_889),
.B(n_512),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_889),
.B(n_504),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_889),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_889),
.B(n_513),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_889),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_887),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_887),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_887),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_887),
.Y(n_959)
);

AO31x2_ASAP7_75t_L g960 ( 
.A1(n_900),
.A2(n_536),
.A3(n_576),
.B(n_568),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_889),
.B(n_519),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_887),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_887),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_903),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_889),
.B(n_525),
.Y(n_965)
);

INVxp67_ASAP7_75t_SL g966 ( 
.A(n_889),
.Y(n_966)
);

AOI221xp5_ASAP7_75t_SL g967 ( 
.A1(n_932),
.A2(n_506),
.B1(n_507),
.B2(n_567),
.C(n_566),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_916),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_914),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_948),
.Y(n_970)
);

AO21x2_ASAP7_75t_L g971 ( 
.A1(n_919),
.A2(n_509),
.B(n_508),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_953),
.B(n_511),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_957),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_963),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_956),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_953),
.B(n_514),
.Y(n_976)
);

AOI221xp5_ASAP7_75t_L g977 ( 
.A1(n_937),
.A2(n_547),
.B1(n_516),
.B2(n_520),
.C(n_564),
.Y(n_977)
);

NAND3xp33_ASAP7_75t_L g978 ( 
.A(n_917),
.B(n_521),
.C(n_515),
.Y(n_978)
);

AOI211xp5_ASAP7_75t_SL g979 ( 
.A1(n_941),
.A2(n_522),
.B(n_524),
.C(n_526),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_955),
.Y(n_980)
);

AO21x2_ASAP7_75t_L g981 ( 
.A1(n_919),
.A2(n_935),
.B(n_946),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_966),
.B(n_527),
.Y(n_982)
);

INVxp67_ASAP7_75t_SL g983 ( 
.A(n_915),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_952),
.B(n_530),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_925),
.B(n_531),
.Y(n_985)
);

CKINVDCx6p67_ASAP7_75t_R g986 ( 
.A(n_929),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_918),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_947),
.B(n_540),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_922),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_924),
.B(n_532),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_L g991 ( 
.A(n_917),
.B(n_548),
.C(n_545),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_921),
.B(n_537),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_949),
.B(n_550),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_958),
.Y(n_994)
);

NOR2x1_ASAP7_75t_R g995 ( 
.A(n_938),
.B(n_541),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_959),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_936),
.A2(n_554),
.B(n_551),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_962),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_926),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_951),
.B(n_558),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_927),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_950),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_923),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_950),
.Y(n_1004)
);

OAI211xp5_ASAP7_75t_L g1005 ( 
.A1(n_944),
.A2(n_560),
.B(n_563),
.C(n_565),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_954),
.B(n_549),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_964),
.Y(n_1007)
);

OAI211xp5_ASAP7_75t_L g1008 ( 
.A1(n_933),
.A2(n_569),
.B(n_562),
.C(n_556),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_920),
.A2(n_552),
.B1(n_604),
.B2(n_91),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_928),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_960),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_940),
.A2(n_88),
.B1(n_89),
.B2(n_92),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_960),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_961),
.B(n_95),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_965),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_945),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_945),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_930),
.B(n_96),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_939),
.B(n_97),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_931),
.B(n_942),
.Y(n_1020)
);

AOI33xp33_ASAP7_75t_L g1021 ( 
.A1(n_928),
.A2(n_98),
.A3(n_102),
.B1(n_103),
.B2(n_105),
.B3(n_106),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_930),
.B(n_107),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_934),
.B(n_960),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_934),
.B(n_108),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_934),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_SL g1026 ( 
.A1(n_943),
.A2(n_109),
.B1(n_112),
.B2(n_116),
.Y(n_1026)
);

OAI31xp33_ASAP7_75t_SL g1027 ( 
.A1(n_917),
.A2(n_117),
.A3(n_119),
.B(n_123),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_916),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_914),
.Y(n_1029)
);

AOI222xp33_ASAP7_75t_L g1030 ( 
.A1(n_932),
.A2(n_129),
.B1(n_132),
.B2(n_135),
.C1(n_138),
.C2(n_143),
.Y(n_1030)
);

INVxp67_ASAP7_75t_L g1031 ( 
.A(n_955),
.Y(n_1031)
);

AO21x2_ASAP7_75t_L g1032 ( 
.A1(n_919),
.A2(n_145),
.B(n_148),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_914),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_953),
.B(n_154),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_929),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_915),
.B(n_155),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_SL g1037 ( 
.A(n_1005),
.B(n_992),
.C(n_1008),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1020),
.B(n_161),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_983),
.B(n_163),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_1025),
.B(n_165),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_1003),
.B(n_166),
.Y(n_1041)
);

CKINVDCx16_ASAP7_75t_R g1042 ( 
.A(n_1015),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_980),
.B(n_167),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_969),
.Y(n_1044)
);

NOR2xp67_ASAP7_75t_L g1045 ( 
.A(n_1031),
.B(n_169),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1002),
.B(n_170),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_969),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_1030),
.A2(n_172),
.B1(n_173),
.B2(n_176),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_994),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_L g1050 ( 
.A(n_1007),
.B(n_178),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_994),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1029),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_989),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1004),
.B(n_179),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_999),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_985),
.B(n_180),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_975),
.B(n_181),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_968),
.B(n_970),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_1001),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1036),
.B(n_185),
.Y(n_1060)
);

AOI211xp5_ASAP7_75t_L g1061 ( 
.A1(n_990),
.A2(n_1027),
.B(n_977),
.C(n_991),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1029),
.Y(n_1062)
);

AND2x2_ASAP7_75t_SL g1063 ( 
.A(n_1021),
.B(n_187),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1033),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_995),
.B(n_1006),
.Y(n_1065)
);

CKINVDCx16_ASAP7_75t_R g1066 ( 
.A(n_1035),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_973),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1033),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_1017),
.B(n_188),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_988),
.B(n_189),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1011),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_974),
.B(n_191),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_996),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_993),
.B(n_194),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1028),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_L g1076 ( 
.A(n_979),
.B(n_199),
.C(n_200),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_998),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_986),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1011),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1013),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1000),
.B(n_201),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1019),
.B(n_202),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_1042),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_1077),
.B(n_1013),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1068),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1044),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1061),
.A2(n_1009),
.B1(n_967),
.B2(n_1017),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_1059),
.B(n_981),
.Y(n_1088)
);

NAND3xp33_ASAP7_75t_L g1089 ( 
.A(n_1037),
.B(n_978),
.C(n_997),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_1053),
.B(n_981),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1073),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1055),
.B(n_987),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1051),
.B(n_1023),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1067),
.B(n_1010),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_1049),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1047),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_1052),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1071),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1062),
.Y(n_1099)
);

NOR2xp67_ASAP7_75t_SL g1100 ( 
.A(n_1076),
.B(n_1018),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1064),
.B(n_1016),
.Y(n_1101)
);

OAI21xp33_ASAP7_75t_L g1102 ( 
.A1(n_1063),
.A2(n_1048),
.B(n_1046),
.Y(n_1102)
);

NAND2xp33_ASAP7_75t_SL g1103 ( 
.A(n_1078),
.B(n_1034),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_1066),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1075),
.B(n_972),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1058),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1038),
.B(n_1024),
.Y(n_1107)
);

NAND2xp33_ASAP7_75t_L g1108 ( 
.A(n_1054),
.B(n_1014),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1065),
.B(n_1070),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1043),
.B(n_982),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1071),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_1079),
.B(n_976),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1074),
.B(n_984),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1081),
.B(n_1032),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1079),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_1040),
.Y(n_1116)
);

INVxp67_ASAP7_75t_SL g1117 ( 
.A(n_1090),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1106),
.B(n_1080),
.Y(n_1118)
);

OAI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1087),
.A2(n_1039),
.B1(n_1045),
.B2(n_1041),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1098),
.Y(n_1120)
);

NAND2x1_ASAP7_75t_L g1121 ( 
.A(n_1085),
.B(n_1080),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1098),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1095),
.B(n_1057),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1091),
.B(n_1040),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1093),
.B(n_1056),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1096),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1092),
.B(n_1032),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1102),
.A2(n_1022),
.B1(n_1026),
.B2(n_1069),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1112),
.B(n_971),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_1115),
.B(n_1069),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1127),
.B(n_1097),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1120),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1125),
.B(n_1083),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1128),
.A2(n_1089),
.B1(n_1116),
.B2(n_1113),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1122),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1117),
.B(n_1086),
.Y(n_1136)
);

XNOR2x1_ASAP7_75t_L g1137 ( 
.A(n_1119),
.B(n_1107),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1126),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_R g1139 ( 
.A(n_1123),
.B(n_1103),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_L g1140 ( 
.A(n_1121),
.B(n_1088),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1129),
.B(n_1099),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1130),
.B(n_1104),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1118),
.B(n_1114),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1124),
.A2(n_1109),
.B1(n_1105),
.B2(n_1094),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_1130),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1130),
.Y(n_1146)
);

OAI21xp33_ASAP7_75t_L g1147 ( 
.A1(n_1128),
.A2(n_1108),
.B(n_1100),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1125),
.B(n_1110),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1147),
.A2(n_1101),
.B(n_1050),
.Y(n_1149)
);

NAND5xp2_ASAP7_75t_L g1150 ( 
.A(n_1147),
.B(n_1082),
.C(n_1060),
.D(n_1072),
.E(n_1111),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1145),
.B(n_1101),
.Y(n_1151)
);

XNOR2x1_ASAP7_75t_L g1152 ( 
.A(n_1137),
.B(n_1012),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1134),
.A2(n_1084),
.B(n_1111),
.C(n_971),
.Y(n_1153)
);

NOR2x1_ASAP7_75t_L g1154 ( 
.A(n_1140),
.B(n_1141),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1144),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_1155)
);

OAI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1131),
.A2(n_210),
.B1(n_211),
.B2(n_215),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_SL g1157 ( 
.A(n_1139),
.B(n_219),
.C(n_224),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1142),
.A2(n_225),
.B1(n_226),
.B2(n_231),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_1133),
.Y(n_1159)
);

AOI322xp5_ASAP7_75t_L g1160 ( 
.A1(n_1148),
.A2(n_233),
.A3(n_235),
.B1(n_240),
.B2(n_241),
.C1(n_242),
.C2(n_244),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1149),
.B(n_1146),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1151),
.Y(n_1162)
);

AOI221xp5_ASAP7_75t_L g1163 ( 
.A1(n_1153),
.A2(n_1136),
.B1(n_1143),
.B2(n_1138),
.C(n_1135),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1159),
.B(n_1152),
.Y(n_1164)
);

AND3x2_ASAP7_75t_L g1165 ( 
.A(n_1157),
.B(n_1132),
.C(n_1154),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1155),
.Y(n_1166)
);

NAND4xp25_ASAP7_75t_L g1167 ( 
.A(n_1150),
.B(n_247),
.C(n_249),
.D(n_250),
.Y(n_1167)
);

NOR2x1p5_ASAP7_75t_L g1168 ( 
.A(n_1167),
.B(n_1162),
.Y(n_1168)
);

AND3x4_ASAP7_75t_L g1169 ( 
.A(n_1161),
.B(n_1160),
.C(n_1156),
.Y(n_1169)
);

AOI211xp5_ASAP7_75t_L g1170 ( 
.A1(n_1166),
.A2(n_1158),
.B(n_256),
.C(n_268),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1165),
.Y(n_1171)
);

AND3x4_ASAP7_75t_L g1172 ( 
.A(n_1169),
.B(n_1164),
.C(n_1163),
.Y(n_1172)
);

AO21x1_ASAP7_75t_L g1173 ( 
.A1(n_1171),
.A2(n_346),
.B(n_273),
.Y(n_1173)
);

OAI222xp33_ASAP7_75t_L g1174 ( 
.A1(n_1168),
.A2(n_253),
.B1(n_274),
.B2(n_278),
.C1(n_281),
.C2(n_282),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_L g1175 ( 
.A(n_1170),
.B(n_284),
.C(n_285),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1172),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1173),
.Y(n_1177)
);

AOI221xp5_ASAP7_75t_L g1178 ( 
.A1(n_1174),
.A2(n_289),
.B1(n_292),
.B2(n_294),
.C(n_295),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1175),
.A2(n_296),
.B(n_297),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1172),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1177),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1176),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1180),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1182),
.Y(n_1184)
);

XOR2xp5_ASAP7_75t_L g1185 ( 
.A(n_1183),
.B(n_1179),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1185),
.A2(n_1181),
.B1(n_1178),
.B2(n_299),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1184),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1186),
.A2(n_344),
.B(n_298),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1188),
.A2(n_1187),
.B1(n_301),
.B2(n_302),
.Y(n_1189)
);


endmodule