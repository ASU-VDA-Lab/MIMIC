module fake_ariane_1372_n_761 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_761);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_761;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_445;
wire n_515;
wire n_379;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_455;
wire n_429;
wire n_365;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_3),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_0),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_47),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_2),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_136),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_105),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_86),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_10),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_7),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_32),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_73),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_58),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_107),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_56),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_90),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_13),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_6),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_22),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_111),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_65),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_63),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_8),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_60),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_49),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_78),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_22),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_30),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_137),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_51),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_66),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_34),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_71),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_43),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_27),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_2),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_0),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_149),
.B(n_1),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_1),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

BUFx8_ASAP7_75t_SL g206 ( 
.A(n_144),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_3),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_4),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_4),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_5),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_142),
.B(n_194),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_5),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_157),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_6),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_192),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_7),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_8),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_151),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_9),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_148),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_147),
.B(n_9),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_169),
.B(n_10),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_147),
.B(n_11),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_141),
.B(n_11),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_158),
.B(n_12),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_201),
.B(n_156),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_144),
.B1(n_165),
.B2(n_171),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_208),
.A2(n_176),
.B1(n_150),
.B2(n_167),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_233),
.A2(n_165),
.B1(n_156),
.B2(n_164),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_206),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_183),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_164),
.B1(n_171),
.B2(n_145),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_160),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_193),
.B1(n_191),
.B2(n_189),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_217),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g245 ( 
.A1(n_208),
.A2(n_188),
.B1(n_187),
.B2(n_186),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_185),
.B1(n_181),
.B2(n_180),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_163),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_179),
.B1(n_178),
.B2(n_173),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_172),
.B1(n_166),
.B2(n_14),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_26),
.Y(n_252)
);

AO22x2_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_15),
.Y(n_254)
);

OR2x6_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_15),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_16),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_16),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_R g258 ( 
.A1(n_199),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_209),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_210),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_210),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_230),
.A2(n_232),
.B1(n_221),
.B2(n_202),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_231),
.A2(n_227),
.B1(n_224),
.B2(n_215),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_218),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_207),
.A2(n_220),
.B1(n_218),
.B2(n_234),
.Y(n_268)
);

AO22x2_ASAP7_75t_L g269 ( 
.A1(n_213),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_218),
.B(n_31),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_213),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_218),
.B(n_37),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_218),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_226),
.B(n_41),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_218),
.B(n_140),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_198),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_195),
.Y(n_278)
);

AO22x2_ASAP7_75t_L g279 ( 
.A1(n_226),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_198),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_223),
.A2(n_198),
.B1(n_200),
.B2(n_216),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_280),
.Y(n_282)
);

BUFx8_ASAP7_75t_L g283 ( 
.A(n_240),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_239),
.B(n_228),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_200),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_241),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_249),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_259),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_255),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_205),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_255),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_248),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_200),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_257),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_244),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_247),
.A2(n_229),
.B(n_228),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_238),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_253),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_267),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_246),
.B(n_228),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_273),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_235),
.B(n_205),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_243),
.B(n_228),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_266),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_271),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_271),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_228),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_261),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_252),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_262),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_237),
.B(n_205),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_250),
.B(n_211),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_277),
.B(n_274),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_245),
.B(n_229),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_258),
.B(n_229),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_280),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_280),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_280),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_242),
.B(n_211),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_317),
.B(n_294),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_289),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_292),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_291),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_211),
.Y(n_351)
);

AND2x2_ASAP7_75t_SL g352 ( 
.A(n_329),
.B(n_204),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

AND2x2_ASAP7_75t_SL g355 ( 
.A(n_311),
.B(n_204),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_328),
.B(n_216),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_299),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g358 ( 
.A(n_302),
.B(n_195),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_296),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_229),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_283),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_229),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_283),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_310),
.B(n_223),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

AND2x2_ASAP7_75t_SL g366 ( 
.A(n_312),
.B(n_195),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_296),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_223),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_225),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_296),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_325),
.B(n_225),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_296),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_303),
.B(n_225),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_282),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_304),
.B(n_225),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_305),
.B(n_225),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_302),
.B(n_225),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_195),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_301),
.B(n_195),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_316),
.B(n_52),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_286),
.Y(n_384)
);

OAI21xp33_ASAP7_75t_L g385 ( 
.A1(n_335),
.A2(n_212),
.B(n_196),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_301),
.B(n_196),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_340),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_317),
.B(n_197),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_334),
.B(n_196),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_320),
.B(n_196),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_337),
.A2(n_197),
.B(n_212),
.Y(n_393)
);

NAND2x1p5_ASAP7_75t_L g394 ( 
.A(n_318),
.B(n_197),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_334),
.B(n_196),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_320),
.B(n_212),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_315),
.B(n_212),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_295),
.B(n_212),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_332),
.B(n_197),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g403 ( 
.A(n_322),
.B(n_327),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_288),
.B(n_197),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_298),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_331),
.B(n_197),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_332),
.B(n_53),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_297),
.B(n_300),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_313),
.B(n_54),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_314),
.Y(n_410)
);

AND2x2_ASAP7_75t_SL g411 ( 
.A(n_339),
.B(n_55),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_298),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_333),
.B(n_57),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_351),
.B(n_321),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_410),
.B(n_321),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_358),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_351),
.B(n_330),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_357),
.B(n_285),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_381),
.B(n_330),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_288),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_403),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_411),
.B(n_306),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_352),
.B(n_306),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_348),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_352),
.B(n_309),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_405),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_405),
.Y(n_429)
);

NAND2x1p5_ASAP7_75t_L g430 ( 
.A(n_354),
.B(n_307),
.Y(n_430)
);

BUFx12f_ASAP7_75t_L g431 ( 
.A(n_353),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_375),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_352),
.B(n_309),
.Y(n_434)
);

NAND2x1_ASAP7_75t_SL g435 ( 
.A(n_368),
.B(n_339),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_358),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_411),
.B(n_284),
.Y(n_437)
);

BUFx12f_ASAP7_75t_L g438 ( 
.A(n_353),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_357),
.B(n_338),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_403),
.B(n_356),
.Y(n_440)
);

NOR2x1_ASAP7_75t_L g441 ( 
.A(n_361),
.B(n_363),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_375),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_326),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_337),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_356),
.B(n_287),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_399),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_324),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_355),
.B(n_287),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_355),
.B(n_285),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_347),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_347),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_350),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_409),
.B(n_324),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_358),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_364),
.B(n_290),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_355),
.B(n_319),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_380),
.B(n_319),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_349),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_349),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_364),
.B(n_308),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_411),
.B(n_59),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_350),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_375),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_368),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_361),
.B(n_61),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_401),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_358),
.Y(n_469)
);

NAND2x1_ASAP7_75t_SL g470 ( 
.A(n_383),
.B(n_62),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_417),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_421),
.B(n_366),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_423),
.A2(n_383),
.B1(n_409),
.B2(n_382),
.Y(n_474)
);

INVx6_ASAP7_75t_L g475 ( 
.A(n_431),
.Y(n_475)
);

INVx6_ASAP7_75t_L g476 ( 
.A(n_438),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_438),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_425),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

CKINVDCx11_ASAP7_75t_R g480 ( 
.A(n_432),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_419),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_444),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_459),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_432),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_467),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_441),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_469),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_432),
.Y(n_489)
);

CKINVDCx6p67_ASAP7_75t_R g490 ( 
.A(n_469),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_445),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_451),
.Y(n_492)
);

NAND2x1p5_ASAP7_75t_L g493 ( 
.A(n_436),
.B(n_455),
.Y(n_493)
);

BUFx12f_ASAP7_75t_L g494 ( 
.A(n_467),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_435),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_432),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_442),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_416),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_448),
.B(n_383),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_445),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_442),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_452),
.Y(n_502)
);

BUFx12f_ASAP7_75t_L g503 ( 
.A(n_445),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_442),
.Y(n_504)
);

BUFx2_ASAP7_75t_SL g505 ( 
.A(n_416),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_453),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_421),
.B(n_366),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_462),
.A2(n_383),
.B1(n_409),
.B2(n_363),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_459),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_450),
.B(n_446),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_442),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_415),
.B(n_440),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_428),
.Y(n_513)
);

NAND2x1p5_ASAP7_75t_L g514 ( 
.A(n_428),
.B(n_354),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_466),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_478),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_474),
.A2(n_462),
.B1(n_463),
.B2(n_420),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_494),
.A2(n_437),
.B1(n_434),
.B2(n_426),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_474),
.A2(n_416),
.B1(n_424),
.B2(n_456),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_494),
.A2(n_426),
.B1(n_434),
.B2(n_449),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_491),
.Y(n_521)
);

BUFx8_ASAP7_75t_SL g522 ( 
.A(n_473),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_508),
.A2(n_418),
.B1(n_414),
.B2(n_422),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_481),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_483),
.Y(n_525)
);

INVx6_ASAP7_75t_L g526 ( 
.A(n_479),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_481),
.A2(n_443),
.B1(n_439),
.B2(n_366),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_511),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_499),
.A2(n_454),
.B1(n_448),
.B2(n_433),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_428),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_499),
.A2(n_448),
.B1(n_454),
.B2(n_447),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_483),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_499),
.A2(n_454),
.B1(n_413),
.B2(n_464),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_473),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_485),
.A2(n_461),
.B1(n_430),
.B2(n_468),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_509),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_479),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_515),
.A2(n_430),
.B1(n_369),
.B2(n_354),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_SL g539 ( 
.A1(n_499),
.A2(n_413),
.B1(n_389),
.B2(n_393),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_515),
.A2(n_369),
.B1(n_354),
.B2(n_387),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_480),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_509),
.Y(n_542)
);

HB1xp67_ASAP7_75t_SL g543 ( 
.A(n_477),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_499),
.A2(n_427),
.B1(n_429),
.B2(n_460),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_492),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_480),
.Y(n_546)
);

BUFx4f_ASAP7_75t_SL g547 ( 
.A(n_477),
.Y(n_547)
);

OAI22xp33_ASAP7_75t_L g548 ( 
.A1(n_512),
.A2(n_457),
.B1(n_369),
.B2(n_360),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_472),
.A2(n_360),
.B1(n_386),
.B2(n_382),
.Y(n_549)
);

INVx11_ASAP7_75t_L g550 ( 
.A(n_503),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_503),
.A2(n_498),
.B1(n_505),
.B2(n_510),
.Y(n_551)
);

CKINVDCx11_ASAP7_75t_R g552 ( 
.A(n_496),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_502),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_490),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_506),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_500),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_491),
.A2(n_429),
.B1(n_427),
.B2(n_460),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_513),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_527),
.A2(n_507),
.B1(n_495),
.B2(n_386),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_541),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_SL g561 ( 
.A1(n_527),
.A2(n_486),
.B1(n_479),
.B2(n_475),
.Y(n_561)
);

AOI222xp33_ASAP7_75t_L g562 ( 
.A1(n_517),
.A2(n_519),
.B1(n_518),
.B2(n_523),
.C1(n_520),
.C2(n_533),
.Y(n_562)
);

OA222x2_ASAP7_75t_L g563 ( 
.A1(n_517),
.A2(n_470),
.B1(n_362),
.B2(n_407),
.C1(n_497),
.C2(n_489),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_524),
.B(n_475),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_541),
.A2(n_486),
.B1(n_475),
.B2(n_476),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_530),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_516),
.B(n_487),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_539),
.A2(n_349),
.B1(n_365),
.B2(n_362),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_535),
.A2(n_551),
.B1(n_556),
.B2(n_545),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_525),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_521),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_532),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_556),
.A2(n_365),
.B1(n_404),
.B2(n_395),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_524),
.A2(n_490),
.B1(n_486),
.B2(n_369),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_521),
.Y(n_576)
);

BUFx4f_ASAP7_75t_SL g577 ( 
.A(n_541),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_554),
.B(n_511),
.Y(n_578)
);

BUFx5_ASAP7_75t_L g579 ( 
.A(n_530),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_536),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_545),
.B(n_513),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_553),
.B(n_513),
.Y(n_582)
);

BUFx4f_ASAP7_75t_SL g583 ( 
.A(n_546),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_532),
.Y(n_584)
);

AOI222xp33_ASAP7_75t_L g585 ( 
.A1(n_553),
.A2(n_408),
.B1(n_393),
.B2(n_395),
.C1(n_390),
.C2(n_396),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_L g586 ( 
.A(n_555),
.B(n_390),
.C(n_387),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_534),
.B(n_476),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_555),
.A2(n_365),
.B1(n_370),
.B2(n_372),
.Y(n_588)
);

NOR2x1_ASAP7_75t_L g589 ( 
.A(n_554),
.B(n_484),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_534),
.B(n_476),
.Y(n_590)
);

OAI21xp33_ASAP7_75t_L g591 ( 
.A1(n_546),
.A2(n_407),
.B(n_396),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_536),
.Y(n_592)
);

BUFx4f_ASAP7_75t_SL g593 ( 
.A(n_546),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_542),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_542),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_549),
.A2(n_380),
.B1(n_358),
.B2(n_488),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_530),
.B(n_484),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_529),
.A2(n_531),
.B1(n_549),
.B2(n_544),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_558),
.B(n_513),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_557),
.A2(n_370),
.B1(n_372),
.B2(n_471),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_558),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_SL g602 ( 
.A1(n_554),
.A2(n_526),
.B1(n_486),
.B2(n_540),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_526),
.A2(n_471),
.B1(n_482),
.B2(n_488),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_530),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_SL g605 ( 
.A1(n_526),
.A2(n_471),
.B1(n_482),
.B2(n_493),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_562),
.A2(n_482),
.B1(n_471),
.B2(n_548),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_559),
.A2(n_538),
.B1(n_543),
.B2(n_358),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_591),
.B(n_537),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_568),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_SL g610 ( 
.A(n_590),
.B(n_388),
.C(n_547),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_598),
.A2(n_482),
.B1(n_375),
.B2(n_397),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_561),
.A2(n_375),
.B1(n_397),
.B2(n_458),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_585),
.A2(n_397),
.B1(n_392),
.B2(n_384),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_570),
.A2(n_574),
.B1(n_586),
.B2(n_588),
.Y(n_614)
);

AOI222xp33_ASAP7_75t_L g615 ( 
.A1(n_569),
.A2(n_388),
.B1(n_406),
.B2(n_376),
.C1(n_400),
.C2(n_384),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_573),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_563),
.A2(n_526),
.B1(n_537),
.B2(n_358),
.Y(n_617)
);

NOR3xp33_ASAP7_75t_L g618 ( 
.A(n_575),
.B(n_552),
.C(n_528),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_596),
.A2(n_493),
.B1(n_379),
.B2(n_537),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_596),
.A2(n_550),
.B1(n_514),
.B2(n_465),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_581),
.B(n_528),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_600),
.A2(n_397),
.B1(n_392),
.B2(n_384),
.Y(n_622)
);

OAI221xp5_ASAP7_75t_SL g623 ( 
.A1(n_563),
.A2(n_565),
.B1(n_602),
.B2(n_572),
.C(n_560),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_587),
.A2(n_528),
.B(n_522),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_581),
.A2(n_397),
.B1(n_392),
.B2(n_376),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_SL g626 ( 
.A1(n_560),
.A2(n_537),
.B1(n_489),
.B2(n_497),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_577),
.A2(n_550),
.B1(n_514),
.B2(n_465),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_582),
.A2(n_397),
.B1(n_400),
.B2(n_376),
.Y(n_628)
);

OAI222xp33_ASAP7_75t_L g629 ( 
.A1(n_605),
.A2(n_400),
.B1(n_394),
.B2(n_378),
.C1(n_377),
.C2(n_374),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_583),
.A2(n_465),
.B1(n_511),
.B2(n_394),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_573),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_584),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_SL g633 ( 
.A1(n_593),
.A2(n_394),
.B1(n_511),
.B2(n_501),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_582),
.A2(n_412),
.B1(n_377),
.B2(n_378),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_576),
.B(n_496),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_594),
.A2(n_412),
.B1(n_374),
.B2(n_371),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_594),
.A2(n_412),
.B1(n_371),
.B2(n_373),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_595),
.A2(n_371),
.B1(n_373),
.B2(n_406),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_584),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_579),
.A2(n_501),
.B1(n_496),
.B2(n_504),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_623),
.B(n_589),
.C(n_601),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_621),
.B(n_567),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_609),
.B(n_604),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_618),
.B(n_589),
.C(n_601),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_621),
.B(n_567),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_635),
.B(n_599),
.C(n_564),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_607),
.A2(n_567),
.B1(n_578),
.B2(n_595),
.Y(n_647)
);

NAND4xp25_ASAP7_75t_L g648 ( 
.A(n_610),
.B(n_599),
.C(n_597),
.D(n_603),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_617),
.A2(n_597),
.B(n_391),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_616),
.B(n_579),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_608),
.B(n_597),
.C(n_391),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_631),
.B(n_579),
.Y(n_652)
);

OAI21xp33_ASAP7_75t_L g653 ( 
.A1(n_608),
.A2(n_398),
.B(n_402),
.Y(n_653)
);

OAI221xp5_ASAP7_75t_L g654 ( 
.A1(n_614),
.A2(n_398),
.B1(n_385),
.B2(n_580),
.C(n_571),
.Y(n_654)
);

AND2x2_ASAP7_75t_SL g655 ( 
.A(n_616),
.B(n_579),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_632),
.B(n_579),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_632),
.B(n_579),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_606),
.B(n_501),
.C(n_496),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_639),
.B(n_579),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_624),
.B(n_579),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_L g661 ( 
.A(n_627),
.B(n_504),
.C(n_367),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_639),
.B(n_566),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_620),
.B(n_566),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_626),
.B(n_501),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_634),
.B(n_592),
.C(n_580),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_611),
.A2(n_367),
.B1(n_359),
.B2(n_373),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_619),
.B(n_571),
.Y(n_667)
);

AOI221xp5_ASAP7_75t_L g668 ( 
.A1(n_613),
.A2(n_385),
.B1(n_592),
.B2(n_402),
.C(n_367),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_645),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_645),
.B(n_640),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_642),
.B(n_612),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_655),
.B(n_625),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_655),
.B(n_650),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_646),
.B(n_628),
.C(n_615),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_643),
.B(n_636),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_SL g676 ( 
.A(n_660),
.B(n_629),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_657),
.B(n_633),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_662),
.Y(n_678)
);

OA211x2_ASAP7_75t_L g679 ( 
.A1(n_653),
.A2(n_664),
.B(n_644),
.C(n_651),
.Y(n_679)
);

AOI211xp5_ASAP7_75t_L g680 ( 
.A1(n_647),
.A2(n_630),
.B(n_367),
.C(n_359),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_656),
.B(n_638),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_658),
.A2(n_622),
.B1(n_637),
.B2(n_359),
.Y(n_682)
);

AND2x6_ASAP7_75t_L g683 ( 
.A(n_659),
.B(n_359),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_652),
.B(n_663),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_667),
.B(n_661),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_641),
.A2(n_64),
.B1(n_68),
.B2(n_69),
.Y(n_686)
);

XNOR2xp5_ASAP7_75t_L g687 ( 
.A(n_670),
.B(n_648),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_678),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_676),
.A2(n_679),
.B1(n_674),
.B2(n_672),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_684),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_670),
.B(n_664),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_685),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_685),
.B(n_647),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_669),
.B(n_661),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_673),
.B(n_649),
.Y(n_695)
);

XOR2x2_ASAP7_75t_L g696 ( 
.A(n_677),
.B(n_665),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_681),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_697),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_690),
.Y(n_699)
);

XNOR2xp5_ASAP7_75t_L g700 ( 
.A(n_687),
.B(n_671),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_688),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_701),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_700),
.A2(n_689),
.B1(n_696),
.B2(n_691),
.Y(n_703)
);

OA22x2_ASAP7_75t_L g704 ( 
.A1(n_700),
.A2(n_691),
.B1(n_693),
.B2(n_692),
.Y(n_704)
);

OA22x2_ASAP7_75t_L g705 ( 
.A1(n_699),
.A2(n_693),
.B1(n_690),
.B2(n_694),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_698),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_702),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_706),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_705),
.Y(n_709)
);

BUFx4f_ASAP7_75t_SL g710 ( 
.A(n_704),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_707),
.Y(n_711)
);

AO22x2_ASAP7_75t_L g712 ( 
.A1(n_709),
.A2(n_698),
.B1(n_703),
.B2(n_675),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_707),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_SL g714 ( 
.A1(n_711),
.A2(n_708),
.B(n_686),
.C(n_695),
.Y(n_714)
);

OA22x2_ASAP7_75t_L g715 ( 
.A1(n_713),
.A2(n_710),
.B1(n_673),
.B2(n_672),
.Y(n_715)
);

AOI221xp5_ASAP7_75t_L g716 ( 
.A1(n_712),
.A2(n_686),
.B1(n_671),
.B2(n_680),
.C(n_654),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_711),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_717),
.B(n_682),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_715),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_716),
.A2(n_683),
.B1(n_682),
.B2(n_666),
.Y(n_720)
);

AOI221xp5_ASAP7_75t_L g721 ( 
.A1(n_714),
.A2(n_668),
.B1(n_683),
.B2(n_79),
.C(n_80),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_715),
.A2(n_683),
.B1(n_74),
.B2(n_81),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_715),
.A2(n_683),
.B1(n_82),
.B2(n_84),
.Y(n_723)
);

NOR2x1_ASAP7_75t_L g724 ( 
.A(n_714),
.B(n_683),
.Y(n_724)
);

NOR2x1_ASAP7_75t_L g725 ( 
.A(n_719),
.B(n_683),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_718),
.B(n_72),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_724),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_721),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_720),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_722),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_723),
.Y(n_731)
);

OAI211xp5_ASAP7_75t_L g732 ( 
.A1(n_727),
.A2(n_728),
.B(n_731),
.C(n_725),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_726),
.Y(n_733)
);

AND4x1_ASAP7_75t_L g734 ( 
.A(n_729),
.B(n_94),
.C(n_95),
.D(n_96),
.Y(n_734)
);

OAI211xp5_ASAP7_75t_L g735 ( 
.A1(n_730),
.A2(n_98),
.B(n_99),
.C(n_100),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_726),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_729),
.Y(n_737)
);

AND4x1_ASAP7_75t_L g738 ( 
.A(n_728),
.B(n_101),
.C(n_102),
.D(n_103),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_733),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_736),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_737),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_734),
.B(n_106),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_732),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_732),
.B(n_108),
.Y(n_744)
);

AO22x2_ASAP7_75t_L g745 ( 
.A1(n_743),
.A2(n_735),
.B1(n_738),
.B2(n_112),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_739),
.Y(n_746)
);

AO22x2_ASAP7_75t_L g747 ( 
.A1(n_740),
.A2(n_109),
.B1(n_110),
.B2(n_113),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_741),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_744),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_742),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_748),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_749),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_746),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_745),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_754),
.A2(n_750),
.B1(n_747),
.B2(n_120),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_752),
.A2(n_751),
.B1(n_753),
.B2(n_121),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_756),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_757),
.A2(n_755),
.B1(n_119),
.B2(n_124),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_758),
.Y(n_759)
);

AOI221xp5_ASAP7_75t_L g760 ( 
.A1(n_759),
.A2(n_117),
.B1(n_125),
.B2(n_126),
.C(n_127),
.Y(n_760)
);

AOI211xp5_ASAP7_75t_L g761 ( 
.A1(n_760),
.A2(n_128),
.B(n_129),
.C(n_132),
.Y(n_761)
);


endmodule