module fake_jpeg_17637_n_88 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_88);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_88;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx10_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_17),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_18),
.B1(n_10),
.B2(n_16),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_10),
.B1(n_22),
.B2(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_20),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_26),
.C(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_12),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

AND2x6_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_0),
.Y(n_41)
);

NOR2xp67_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_10),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_50),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_35),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_9),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_36),
.B(n_38),
.C(n_33),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_16),
.B(n_13),
.Y(n_68)
);

NAND4xp25_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_40),
.C(n_23),
.D(n_9),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_54),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_35),
.B1(n_15),
.B2(n_11),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_14),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_12),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_47),
.B(n_43),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_68),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_51),
.C(n_46),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_66),
.C(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_35),
.Y(n_67)
);

OAI321xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_52),
.A3(n_55),
.B1(n_58),
.B2(n_54),
.C(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_58),
.B1(n_13),
.B2(n_9),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_64),
.C(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_76),
.C(n_72),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_72),
.B(n_7),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_79),
.B(n_6),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_82),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_75),
.B1(n_6),
.B2(n_2),
.Y(n_83)
);

AOI322xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_4),
.C1(n_5),
.C2(n_82),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_5),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_85),
.C(n_0),
.Y(n_87)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_4),
.CI(n_82),
.CON(n_88),
.SN(n_88)
);


endmodule