module fake_netlist_5_846_n_1841 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1841);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1841;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_10),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_118),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_158),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_47),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_42),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_64),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_94),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_59),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_122),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_72),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_74),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_7),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_134),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_26),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_6),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_33),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_12),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_31),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_65),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_97),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_71),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_38),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_103),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_138),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_33),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_110),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_75),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_53),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_5),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_46),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_93),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_132),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_147),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_60),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_151),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_91),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_26),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_67),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_121),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_41),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_17),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_69),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_43),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_2),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_7),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_68),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_79),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_100),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_61),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_130),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_34),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_135),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_57),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_5),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_87),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_36),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_131),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_39),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_58),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_47),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_85),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_150),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_11),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_62),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_96),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_10),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_13),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_24),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_137),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_29),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_54),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_144),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_55),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_88),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_29),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_111),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_25),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_159),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_31),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_129),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_51),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_125),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_119),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_25),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_99),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_90),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_145),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_46),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_83),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_49),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_44),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_126),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_32),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_37),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_44),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_52),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_27),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_73),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_14),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_36),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_32),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_89),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_49),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_19),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_38),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_0),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_1),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_84),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_81),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_80),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_43),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_112),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_50),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_149),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_148),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_143),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_105),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_22),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_133),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_66),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_19),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_52),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_17),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_24),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_34),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_37),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_77),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_127),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_2),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_16),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_53),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_120),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_136),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_11),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_123),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_155),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_35),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_35),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_15),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_142),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_102),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_42),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_28),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_6),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_22),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_41),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_108),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_174),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_297),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_191),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_178),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_168),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_297),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_162),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_297),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_250),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_167),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_169),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_297),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_177),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_179),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_191),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_314),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_181),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_225),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_250),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_233),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_184),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_233),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_303),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_185),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_192),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_189),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_235),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_185),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_189),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_204),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_204),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_323),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_255),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_323),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_185),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_255),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_317),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_243),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_317),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_243),
.Y(n_371)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_163),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_243),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_276),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_276),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_193),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_276),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_165),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_194),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_195),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_165),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_180),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_170),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_232),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_197),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_170),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_190),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_190),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_317),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_196),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_232),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_213),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_198),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_196),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_217),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_200),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_163),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_298),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_217),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_202),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_221),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_206),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_166),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_221),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_227),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_331),
.B(n_284),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_397),
.B(n_284),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_354),
.B(n_298),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_325),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_335),
.B(n_175),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_336),
.B(n_338),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_325),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_339),
.B(n_262),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_344),
.B(n_350),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_326),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_391),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_397),
.B(n_175),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_355),
.B(n_376),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_379),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_373),
.B(n_211),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_332),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_333),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_337),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_337),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g435 ( 
.A(n_341),
.B(n_211),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_380),
.B(n_285),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_347),
.B(n_282),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_343),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_396),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_247),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_343),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_348),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_349),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_356),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_373),
.B(n_247),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_327),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_356),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_403),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_382),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_402),
.B(n_268),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_353),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

BUFx8_ASAP7_75t_L g458 ( 
.A(n_340),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_385),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_378),
.Y(n_461)
);

BUFx8_ASAP7_75t_L g462 ( 
.A(n_340),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_353),
.Y(n_463)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_372),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_372),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_334),
.B(n_268),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_381),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_381),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_324),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_383),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_393),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_346),
.B(n_207),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_386),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_386),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_351),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_387),
.Y(n_478)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_372),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_417),
.B(n_365),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_436),
.B(n_329),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_418),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_409),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_422),
.B(n_384),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_L g486 ( 
.A(n_414),
.B(n_208),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_460),
.Y(n_487)
);

AND3x2_ASAP7_75t_L g488 ( 
.A(n_422),
.B(n_216),
.C(n_164),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_409),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_418),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_424),
.Y(n_491)
);

INVx5_ASAP7_75t_L g492 ( 
.A(n_408),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_437),
.A2(n_313),
.B1(n_272),
.B2(n_321),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_420),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_451),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_463),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_412),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_412),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_430),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_413),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_430),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_463),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_432),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_451),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_416),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_426),
.B(n_392),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_415),
.A2(n_352),
.B1(n_389),
.B2(n_359),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_416),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_443),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_463),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_443),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_SL g515 ( 
.A(n_411),
.B(n_257),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_469),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_406),
.B(n_366),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_410),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_440),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_455),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_428),
.B(n_368),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_474),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_441),
.B(n_210),
.Y(n_525)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_460),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_453),
.B(n_370),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_421),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_431),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_410),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_431),
.Y(n_531)
);

OAI22xp33_ASAP7_75t_L g532 ( 
.A1(n_449),
.A2(n_289),
.B1(n_277),
.B2(n_251),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_431),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_439),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_411),
.B(n_214),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_439),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_424),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_473),
.B(n_369),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_407),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_432),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_439),
.Y(n_542)
);

AO22x2_ASAP7_75t_L g543 ( 
.A1(n_407),
.A2(n_257),
.B1(n_230),
.B2(n_234),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_434),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g545 ( 
.A1(n_458),
.A2(n_244),
.B1(n_328),
.B2(n_345),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_447),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_424),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_428),
.A2(n_372),
.B1(n_306),
.B2(n_230),
.Y(n_548)
);

NOR2xp67_ASAP7_75t_L g549 ( 
.A(n_455),
.B(n_215),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_460),
.B(n_166),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g551 ( 
.A(n_474),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_419),
.B(n_369),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_447),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_425),
.B(n_371),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_466),
.B(n_371),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_434),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_438),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_407),
.B(n_222),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_451),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_SL g560 ( 
.A(n_477),
.B(n_171),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_438),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_435),
.B(n_223),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_455),
.B(n_224),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_447),
.Y(n_564)
);

CKINVDCx6p67_ASAP7_75t_R g565 ( 
.A(n_452),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_455),
.B(n_374),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_455),
.B(n_228),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_442),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_442),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_455),
.B(n_229),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_428),
.A2(n_372),
.B1(n_270),
.B2(n_271),
.Y(n_571)
);

CKINVDCx6p67_ASAP7_75t_R g572 ( 
.A(n_452),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_460),
.B(n_374),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_424),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_427),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_458),
.B(n_231),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_427),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_445),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_445),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_427),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_427),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_423),
.B(n_428),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_457),
.B(n_375),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_427),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_423),
.B(n_377),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_479),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_427),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_429),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_446),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_L g590 ( 
.A1(n_457),
.A2(n_242),
.B1(n_269),
.B2(n_273),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_451),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_423),
.B(n_377),
.Y(n_592)
);

CKINVDCx14_ASAP7_75t_R g593 ( 
.A(n_459),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_446),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_450),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_448),
.B(n_237),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_450),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_451),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_461),
.B(n_467),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_448),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_472),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_448),
.B(n_238),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_458),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_454),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_448),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_454),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_454),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_454),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_461),
.B(n_358),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_454),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_456),
.B(n_465),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_429),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_435),
.B(n_240),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_456),
.B(n_248),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_429),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_458),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_467),
.B(n_387),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_429),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_454),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_468),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_429),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_468),
.B(n_183),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_464),
.Y(n_623)
);

AOI21x1_ASAP7_75t_L g624 ( 
.A1(n_470),
.A2(n_173),
.B(n_172),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_462),
.B(n_252),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_470),
.A2(n_227),
.B1(n_322),
.B2(n_234),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_471),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_471),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_552),
.B(n_465),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_600),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_554),
.B(n_465),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_540),
.B(n_408),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_551),
.B(n_186),
.Y(n_633)
);

BUFx5_ASAP7_75t_L g634 ( 
.A(n_586),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_540),
.A2(n_292),
.B1(n_288),
.B2(n_254),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_517),
.B(n_462),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_550),
.A2(n_275),
.B1(n_283),
.B2(n_306),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_539),
.B(n_408),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_483),
.Y(n_639)
);

NOR3xp33_ASAP7_75t_L g640 ( 
.A(n_509),
.B(n_590),
.C(n_515),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_600),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_480),
.B(n_481),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_603),
.B(n_236),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_599),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_527),
.B(n_462),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_523),
.B(n_408),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_497),
.B(n_475),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_605),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_524),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_523),
.A2(n_290),
.B1(n_258),
.B2(n_259),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_536),
.B(n_188),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_603),
.B(n_236),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_503),
.B(n_462),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_523),
.B(n_433),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_503),
.B(n_261),
.Y(n_655)
);

NOR3xp33_ASAP7_75t_L g656 ( 
.A(n_609),
.B(n_173),
.C(n_172),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_605),
.Y(n_657)
);

AND2x4_ASAP7_75t_SL g658 ( 
.A(n_565),
.B(n_176),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_523),
.B(n_433),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_524),
.B(n_475),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g661 ( 
.A(n_521),
.B(n_265),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_532),
.B(n_182),
.C(n_176),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_582),
.A2(n_263),
.B1(n_291),
.B2(n_286),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_620),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_617),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_497),
.B(n_274),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_483),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_487),
.B(n_433),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_483),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_620),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_512),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_526),
.B(n_555),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_525),
.B(n_199),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_L g674 ( 
.A1(n_493),
.A2(n_283),
.B1(n_281),
.B2(n_280),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_617),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_627),
.B(n_433),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_512),
.B(n_295),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_622),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_492),
.B(n_296),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_611),
.A2(n_464),
.B(n_478),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_592),
.B(n_476),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_492),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_592),
.B(n_476),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_627),
.B(n_479),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_628),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_628),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_484),
.B(n_203),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_550),
.A2(n_322),
.B1(n_281),
.B2(n_280),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_585),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_482),
.B(n_490),
.Y(n_690)
);

NOR2xp67_ASAP7_75t_L g691 ( 
.A(n_601),
.B(n_478),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_493),
.B(n_388),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_593),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_583),
.A2(n_388),
.B(n_390),
.C(n_405),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_489),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_596),
.B(n_308),
.Y(n_696)
);

O2A1O1Ixp5_ASAP7_75t_L g697 ( 
.A1(n_573),
.A2(n_241),
.B(n_182),
.C(n_187),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_482),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_602),
.B(n_309),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_489),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_558),
.B(n_205),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_490),
.A2(n_390),
.B(n_394),
.C(n_405),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_494),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_489),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_486),
.B(n_219),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_550),
.A2(n_246),
.B1(n_270),
.B2(n_271),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_494),
.B(n_479),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_514),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_495),
.B(n_312),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_520),
.B(n_394),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_495),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_500),
.B(n_316),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_500),
.B(n_479),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_614),
.A2(n_560),
.B1(n_550),
.B2(n_576),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_502),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_626),
.B(n_220),
.C(n_239),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_530),
.B(n_395),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_502),
.B(n_505),
.Y(n_718)
);

OAI22xp33_ASAP7_75t_L g719 ( 
.A1(n_505),
.A2(n_246),
.B1(n_275),
.B2(n_241),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_514),
.Y(n_720)
);

A2O1A1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_541),
.A2(n_212),
.B(n_209),
.C(n_201),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_544),
.B(n_429),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_544),
.Y(n_723)
);

INVx8_ASAP7_75t_L g724 ( 
.A(n_550),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_616),
.B(n_508),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_516),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_556),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_556),
.B(n_395),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_557),
.B(n_561),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_543),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_557),
.B(n_444),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_625),
.B(n_253),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_514),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_496),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_561),
.Y(n_735)
);

OAI221xp5_ASAP7_75t_L g736 ( 
.A1(n_548),
.A2(n_209),
.B1(n_212),
.B2(n_218),
.C(n_226),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_578),
.B(n_444),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_578),
.A2(n_399),
.B(n_401),
.C(n_404),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_579),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_565),
.B(n_399),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_589),
.B(n_218),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_589),
.A2(n_226),
.B(n_245),
.C(n_249),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_594),
.B(n_260),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_518),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_594),
.B(n_401),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_571),
.B(n_245),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_518),
.Y(n_747)
);

AO22x2_ASAP7_75t_L g748 ( 
.A1(n_543),
.A2(n_304),
.B1(n_293),
.B2(n_291),
.Y(n_748)
);

INVx8_ASAP7_75t_L g749 ( 
.A(n_550),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_586),
.B(n_444),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_568),
.Y(n_751)
);

INVxp33_ASAP7_75t_L g752 ( 
.A(n_545),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_562),
.A2(n_404),
.B(n_362),
.C(n_367),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_572),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_518),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_488),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_586),
.B(n_568),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_543),
.Y(n_758)
);

AO22x2_ASAP7_75t_L g759 ( 
.A1(n_543),
.A2(n_293),
.B1(n_286),
.B2(n_278),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_569),
.Y(n_760)
);

OAI221xp5_ASAP7_75t_L g761 ( 
.A1(n_569),
.A2(n_311),
.B1(n_304),
.B2(n_249),
.C(n_278),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_595),
.B(n_444),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_595),
.B(n_444),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_597),
.B(n_444),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_550),
.B(n_256),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_485),
.B(n_256),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_485),
.B(n_263),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_485),
.B(n_491),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_572),
.B(n_264),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_607),
.B(n_266),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_485),
.B(n_311),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_607),
.A2(n_464),
.B(n_357),
.Y(n_772)
);

NOR2xp67_ASAP7_75t_L g773 ( 
.A(n_566),
.B(n_56),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_624),
.B(n_287),
.C(n_279),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_501),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_491),
.B(n_435),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_619),
.B(n_267),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_501),
.A2(n_435),
.B1(n_318),
.B2(n_315),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_496),
.Y(n_779)
);

OR2x6_ASAP7_75t_L g780 ( 
.A(n_624),
.B(n_357),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_504),
.B(n_367),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_491),
.B(n_435),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_598),
.B(n_310),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_491),
.B(n_435),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_528),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_533),
.B(n_435),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_504),
.B(n_364),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_533),
.B(n_464),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_533),
.B(n_464),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_528),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_507),
.A2(n_510),
.B(n_511),
.C(n_513),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_717),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_671),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_630),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_710),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_641),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_678),
.B(n_619),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_685),
.B(n_621),
.Y(n_798)
);

OAI22xp33_ASAP7_75t_L g799 ( 
.A1(n_644),
.A2(n_320),
.B1(n_319),
.B2(n_307),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_685),
.B(n_621),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_685),
.B(n_574),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_734),
.Y(n_802)
);

BUFx4f_ASAP7_75t_SL g803 ( 
.A(n_754),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_648),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_649),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_657),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_639),
.Y(n_807)
);

BUFx12f_ASAP7_75t_L g808 ( 
.A(n_726),
.Y(n_808)
);

AND2x6_ASAP7_75t_L g809 ( 
.A(n_714),
.B(n_598),
.Y(n_809)
);

OAI22xp33_ASAP7_75t_L g810 ( 
.A1(n_644),
.A2(n_678),
.B1(n_729),
.B2(n_690),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_672),
.B(n_533),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_649),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_646),
.A2(n_623),
.B(n_464),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_681),
.B(n_604),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_671),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_671),
.B(n_538),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_693),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_689),
.B(n_538),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_629),
.B(n_538),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_R g820 ( 
.A(n_633),
.B(n_613),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_667),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_631),
.B(n_638),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_654),
.B(n_574),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_751),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_659),
.A2(n_623),
.B(n_496),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_640),
.B(n_574),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_681),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_658),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_665),
.Y(n_829)
);

AND2x6_ASAP7_75t_L g830 ( 
.A(n_740),
.B(n_664),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_675),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_647),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_660),
.Y(n_833)
);

OR2x6_ASAP7_75t_L g834 ( 
.A(n_756),
.B(n_360),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_683),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_640),
.B(n_577),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_728),
.B(n_604),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_634),
.B(n_577),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_634),
.B(n_577),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_642),
.A2(n_570),
.B1(n_563),
.B2(n_567),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_734),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_760),
.Y(n_842)
);

CKINVDCx8_ASAP7_75t_R g843 ( 
.A(n_643),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_670),
.A2(n_608),
.B1(n_606),
.B2(n_615),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_781),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_669),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_634),
.B(n_580),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_692),
.B(n_294),
.Y(n_848)
);

BUFx12f_ASAP7_75t_L g849 ( 
.A(n_643),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_662),
.A2(n_511),
.B1(n_507),
.B2(n_510),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_758),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_686),
.B(n_547),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_734),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_695),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_698),
.B(n_547),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_634),
.B(n_580),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_703),
.B(n_575),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_711),
.B(n_575),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_728),
.B(n_606),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_634),
.B(n_580),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_787),
.Y(n_861)
);

NOR3xp33_ASAP7_75t_SL g862 ( 
.A(n_674),
.B(n_299),
.C(n_300),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_715),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_779),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_634),
.B(n_581),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_691),
.B(n_581),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_700),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_723),
.B(n_575),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_730),
.A2(n_513),
.B(n_553),
.C(n_546),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_727),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_704),
.Y(n_871)
);

BUFx4f_ASAP7_75t_L g872 ( 
.A(n_643),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_SL g873 ( 
.A(n_656),
.B(n_301),
.C(n_302),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_662),
.A2(n_498),
.B1(n_499),
.B2(n_564),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_730),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_769),
.B(n_305),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_735),
.B(n_608),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_739),
.B(n_581),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_743),
.B(n_718),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_SL g880 ( 
.A1(n_636),
.A2(n_651),
.B1(n_732),
.B2(n_687),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_708),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_720),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_779),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_733),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_632),
.B(n_584),
.Y(n_885)
);

NAND2x1p5_ASAP7_75t_L g886 ( 
.A(n_745),
.B(n_584),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_745),
.B(n_584),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_775),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_655),
.B(n_360),
.Y(n_889)
);

AND2x6_ASAP7_75t_SL g890 ( 
.A(n_652),
.B(n_651),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_722),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_676),
.B(n_587),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_731),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_770),
.B(n_777),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_653),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_R g896 ( 
.A(n_661),
.B(n_70),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_737),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_705),
.B(n_587),
.Y(n_898)
);

INVx4_ASAP7_75t_R g899 ( 
.A(n_725),
.Y(n_899)
);

BUFx12f_ASAP7_75t_L g900 ( 
.A(n_652),
.Y(n_900)
);

OR2x6_ASAP7_75t_L g901 ( 
.A(n_652),
.B(n_361),
.Y(n_901)
);

AO22x1_ASAP7_75t_L g902 ( 
.A1(n_656),
.A2(n_361),
.B1(n_362),
.B2(n_364),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_673),
.B(n_668),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_768),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_744),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_783),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_701),
.B(n_588),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_736),
.A2(n_637),
.B1(n_688),
.B2(n_706),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_SL g909 ( 
.A1(n_724),
.A2(n_588),
.B1(n_618),
.B2(n_615),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_716),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_752),
.B(n_588),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_747),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_755),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_757),
.B(n_612),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_785),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_790),
.B(n_612),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_645),
.B(n_498),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_724),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_SL g919 ( 
.A(n_674),
.B(n_0),
.C(n_1),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_736),
.A2(n_637),
.B1(n_688),
.B2(n_706),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_766),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_684),
.B(n_707),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_767),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_724),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_748),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_771),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_748),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_791),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_748),
.A2(n_499),
.B1(n_546),
.B2(n_553),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_709),
.B(n_618),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_762),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_759),
.B(n_542),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_763),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_780),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_780),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_764),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_749),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_712),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_776),
.Y(n_939)
);

BUFx8_ASAP7_75t_L g940 ( 
.A(n_719),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_741),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_666),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_782),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_713),
.B(n_615),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_784),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_650),
.B(n_496),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_677),
.Y(n_947)
);

INVxp67_ASAP7_75t_SL g948 ( 
.A(n_750),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_759),
.A2(n_542),
.B1(n_564),
.B2(n_529),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_786),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_765),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_749),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_759),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_696),
.B(n_534),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_697),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_682),
.B(n_623),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_774),
.A2(n_534),
.B1(n_528),
.B2(n_529),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_699),
.B(n_496),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_635),
.B(n_506),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_774),
.B(n_746),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_702),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_697),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_788),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_778),
.B(n_535),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_749),
.A2(n_506),
.B1(n_610),
.B2(n_591),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_773),
.A2(n_506),
.B1(n_610),
.B2(n_591),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_789),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_761),
.A2(n_535),
.B1(n_529),
.B2(n_531),
.Y(n_968)
);

INVx5_ASAP7_75t_L g969 ( 
.A(n_682),
.Y(n_969)
);

INVxp67_ASAP7_75t_L g970 ( 
.A(n_719),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_680),
.B(n_623),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_761),
.A2(n_506),
.B1(n_591),
.B2(n_559),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_663),
.B(n_506),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_L g974 ( 
.A(n_694),
.B(n_549),
.C(n_531),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_679),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_808),
.B(n_738),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_851),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_851),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_805),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_880),
.B(n_894),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_822),
.B(n_694),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_908),
.A2(n_738),
.B(n_702),
.C(n_753),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_875),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_903),
.B(n_680),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_875),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_794),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_802),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_969),
.A2(n_753),
.B(n_559),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_826),
.A2(n_772),
.B(n_549),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_817),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_810),
.B(n_742),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_810),
.A2(n_721),
.B(n_772),
.C(n_537),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_795),
.B(n_3),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_805),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_797),
.B(n_537),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_803),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_802),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_802),
.Y(n_998)
);

BUFx4f_ASAP7_75t_L g999 ( 
.A(n_830),
.Y(n_999)
);

HAxp5_ASAP7_75t_L g1000 ( 
.A(n_940),
.B(n_3),
.CON(n_1000),
.SN(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_835),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_792),
.B(n_531),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_803),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_797),
.B(n_537),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_908),
.B(n_610),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_898),
.A2(n_559),
.B(n_519),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_911),
.B(n_534),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_812),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_836),
.A2(n_522),
.B(n_559),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_920),
.B(n_559),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_802),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_948),
.A2(n_519),
.B(n_522),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_920),
.B(n_519),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_833),
.B(n_4),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_841),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_796),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_863),
.Y(n_1017)
);

NAND2xp33_ASAP7_75t_SL g1018 ( 
.A(n_896),
.B(n_519),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_881),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_841),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_970),
.B(n_4),
.Y(n_1021)
);

AO21x1_ASAP7_75t_L g1022 ( 
.A1(n_836),
.A2(n_907),
.B(n_946),
.Y(n_1022)
);

O2A1O1Ixp5_ASAP7_75t_L g1023 ( 
.A1(n_866),
.A2(n_161),
.B(n_160),
.C(n_156),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_841),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_884),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_879),
.B(n_152),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_841),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_960),
.B(n_141),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_SL g1029 ( 
.A1(n_943),
.A2(n_8),
.B(n_9),
.C(n_12),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_835),
.B(n_8),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_909),
.A2(n_117),
.B1(n_116),
.B2(n_113),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_812),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_870),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_SL g1034 ( 
.A1(n_895),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_819),
.A2(n_109),
.B(n_104),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_919),
.A2(n_911),
.B(n_862),
.C(n_961),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_966),
.A2(n_98),
.B(n_92),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_946),
.A2(n_15),
.B(n_16),
.C(n_18),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_845),
.B(n_18),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_817),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_953),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_832),
.A2(n_86),
.B1(n_82),
.B2(n_78),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_861),
.B(n_891),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_825),
.A2(n_76),
.B(n_21),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_922),
.A2(n_20),
.B(n_23),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_846),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_922),
.A2(n_27),
.B(n_28),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_893),
.B(n_30),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_883),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_848),
.B(n_829),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_R g1051 ( 
.A(n_828),
.B(n_873),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_883),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_804),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_806),
.A2(n_30),
.B(n_40),
.C(n_45),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_811),
.A2(n_51),
.B(n_45),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_897),
.B(n_50),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_960),
.B(n_40),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_890),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_912),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_934),
.B(n_48),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_934),
.B(n_48),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_829),
.B(n_831),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_830),
.B(n_827),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_830),
.B(n_827),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_838),
.A2(n_860),
.B(n_839),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_910),
.A2(n_799),
.B(n_938),
.C(n_927),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_SL g1067 ( 
.A(n_896),
.B(n_820),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_831),
.B(n_832),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_888),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_912),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_913),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_830),
.B(n_936),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_876),
.B(n_834),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_799),
.A2(n_927),
.B(n_925),
.C(n_889),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_824),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_925),
.A2(n_842),
.B(n_941),
.C(n_869),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_838),
.A2(n_865),
.B(n_860),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_932),
.A2(n_940),
.B1(n_951),
.B2(n_939),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_883),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_959),
.A2(n_935),
.B1(n_926),
.B2(n_921),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_928),
.A2(n_959),
.B(n_973),
.C(n_950),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_935),
.B(n_840),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_913),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_830),
.B(n_936),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_905),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_L g1086 ( 
.A(n_849),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_931),
.B(n_933),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_882),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_837),
.B(n_859),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_SL g1090 ( 
.A(n_866),
.B(n_887),
.C(n_973),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_878),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_901),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_SL g1093 ( 
.A(n_820),
.B(n_843),
.C(n_917),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_906),
.A2(n_942),
.B(n_947),
.C(n_834),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_877),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_807),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_964),
.A2(n_823),
.B(n_818),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_837),
.B(n_859),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_793),
.B(n_815),
.Y(n_1099)
);

AOI21x1_ASAP7_75t_L g1100 ( 
.A1(n_885),
.A2(n_823),
.B(n_865),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_900),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_904),
.B(n_923),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_915),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_939),
.A2(n_945),
.B(n_930),
.C(n_962),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_834),
.B(n_975),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_899),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_883),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_901),
.Y(n_1108)
);

O2A1O1Ixp5_ASAP7_75t_L g1109 ( 
.A1(n_958),
.A2(n_955),
.B(n_971),
.C(n_885),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_814),
.B(n_967),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_901),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_821),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_904),
.B(n_923),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_814),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_854),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_872),
.A2(n_902),
.B1(n_929),
.B2(n_949),
.C(n_850),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_963),
.B(n_867),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_872),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_954),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_924),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_852),
.B(n_855),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_886),
.B(n_871),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_886),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_916),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1065),
.A2(n_944),
.B(n_856),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_984),
.A2(n_965),
.B(n_958),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1016),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1120),
.Y(n_1128)
);

AOI31xp67_ASAP7_75t_L g1129 ( 
.A1(n_980),
.A2(n_984),
.A3(n_1026),
.B(n_1082),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1017),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_1040),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1018),
.A2(n_956),
.B(n_914),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1100),
.A2(n_944),
.B(n_847),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_987),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_SL g1135 ( 
.A1(n_980),
.A2(n_801),
.B(n_800),
.C(n_798),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_1118),
.B(n_952),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1119),
.B(n_1087),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1081),
.A2(n_956),
.B(n_892),
.Y(n_1138)
);

NOR3xp33_ASAP7_75t_L g1139 ( 
.A(n_1093),
.B(n_930),
.C(n_974),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_981),
.A2(n_918),
.B1(n_952),
.B2(n_924),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1081),
.A2(n_809),
.B(n_957),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1043),
.B(n_850),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_SL g1143 ( 
.A1(n_1036),
.A2(n_801),
.B(n_798),
.C(n_800),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1041),
.A2(n_949),
.B1(n_929),
.B2(n_968),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1033),
.Y(n_1145)
);

AO32x2_ASAP7_75t_L g1146 ( 
.A1(n_1080),
.A2(n_844),
.A3(n_972),
.B1(n_853),
.B2(n_809),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_1111),
.B(n_952),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1022),
.A2(n_892),
.B(n_856),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1109),
.A2(n_809),
.B(n_957),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1077),
.A2(n_847),
.B(n_839),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1062),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1082),
.A2(n_971),
.B(n_868),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1095),
.B(n_809),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_986),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_990),
.Y(n_1155)
);

AOI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_1066),
.A2(n_1050),
.B(n_1074),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_SL g1157 ( 
.A1(n_1076),
.A2(n_858),
.B(n_857),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1104),
.A2(n_809),
.B(n_874),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1069),
.Y(n_1159)
);

AOI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_1094),
.A2(n_1113),
.B(n_1102),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1006),
.A2(n_989),
.B(n_988),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1097),
.A2(n_816),
.B(n_813),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1005),
.A2(n_937),
.B(n_952),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1075),
.Y(n_1164)
);

OA21x2_ASAP7_75t_L g1165 ( 
.A1(n_1104),
.A2(n_1090),
.B(n_1009),
.Y(n_1165)
);

CKINVDCx11_ASAP7_75t_R g1166 ( 
.A(n_996),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_987),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1001),
.B(n_924),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_SL g1169 ( 
.A1(n_1116),
.A2(n_924),
.B(n_853),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1001),
.B(n_864),
.Y(n_1170)
);

AOI21xp33_ASAP7_75t_L g1171 ( 
.A1(n_1073),
.A2(n_874),
.B(n_1105),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1005),
.A2(n_1013),
.B(n_1010),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_982),
.A2(n_991),
.A3(n_1036),
.B(n_1121),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_996),
.B(n_1003),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_L g1175 ( 
.A(n_1057),
.B(n_1038),
.C(n_1021),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1091),
.B(n_1021),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1090),
.A2(n_1028),
.B(n_982),
.C(n_1105),
.Y(n_1177)
);

AOI221xp5_ASAP7_75t_L g1178 ( 
.A1(n_993),
.A2(n_1057),
.B1(n_1041),
.B2(n_1038),
.C(n_1034),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1078),
.A2(n_1114),
.B1(n_1098),
.B2(n_1089),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1124),
.B(n_1114),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_SL g1181 ( 
.A1(n_1028),
.A2(n_1026),
.B(n_1013),
.C(n_1010),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_992),
.A2(n_1121),
.B(n_1007),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1044),
.A2(n_1045),
.B(n_1047),
.C(n_1056),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_1031),
.A2(n_1055),
.B(n_1037),
.Y(n_1184)
);

CKINVDCx6p67_ASAP7_75t_R g1185 ( 
.A(n_1003),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_995),
.A2(n_1004),
.A3(n_1054),
.B(n_1072),
.Y(n_1186)
);

AOI21xp33_ASAP7_75t_L g1187 ( 
.A1(n_1078),
.A2(n_1068),
.B(n_1110),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_983),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_987),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_985),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1012),
.A2(n_999),
.B(n_1084),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_979),
.B(n_994),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1000),
.B(n_1030),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1054),
.A2(n_1048),
.A3(n_1035),
.B(n_1063),
.Y(n_1194)
);

OA21x2_ASAP7_75t_L g1195 ( 
.A1(n_1023),
.A2(n_1117),
.B(n_1064),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1110),
.A2(n_1025),
.B(n_1046),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1002),
.B(n_1053),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1089),
.A2(n_1098),
.B1(n_999),
.B2(n_1068),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1019),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1008),
.B(n_1032),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1067),
.A2(n_1123),
.B(n_1122),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1099),
.A2(n_1085),
.B(n_1020),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1106),
.B(n_1051),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1088),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1060),
.A2(n_1061),
.B(n_1120),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_987),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_L g1207 ( 
.A(n_1060),
.B(n_1061),
.C(n_1030),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1039),
.A2(n_1115),
.B(n_1096),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1015),
.B(n_1107),
.Y(n_1209)
);

BUFx8_ASAP7_75t_L g1210 ( 
.A(n_1092),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1042),
.A2(n_1049),
.B(n_1027),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_998),
.A2(n_1079),
.B(n_1052),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_977),
.B(n_978),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_1014),
.A2(n_1112),
.A3(n_1059),
.B(n_1083),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_1108),
.B(n_976),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_L g1216 ( 
.A(n_993),
.B(n_1014),
.C(n_1103),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_1070),
.A2(n_1071),
.A3(n_1107),
.B(n_1024),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_998),
.A2(n_1020),
.B(n_1052),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1079),
.B(n_1051),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_997),
.A2(n_1027),
.B(n_1049),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1015),
.B(n_1024),
.Y(n_1221)
);

NAND2xp33_ASAP7_75t_L g1222 ( 
.A(n_997),
.B(n_1011),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_997),
.A2(n_1049),
.B(n_1011),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1029),
.A2(n_1000),
.A3(n_997),
.B(n_1027),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1029),
.A2(n_976),
.B(n_1058),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1011),
.B(n_1027),
.Y(n_1226)
);

OA22x2_ASAP7_75t_L g1227 ( 
.A1(n_976),
.A2(n_1086),
.B1(n_1101),
.B2(n_1011),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1049),
.A2(n_822),
.B(n_903),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1086),
.A2(n_1065),
.B(n_1100),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1016),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_990),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1065),
.A2(n_1100),
.B(n_1077),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1119),
.B(n_644),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_984),
.A2(n_822),
.B(n_903),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1081),
.A2(n_952),
.B(n_924),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1065),
.A2(n_1100),
.B(n_1077),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1016),
.Y(n_1237)
);

AO21x2_ASAP7_75t_L g1238 ( 
.A1(n_980),
.A2(n_1022),
.B(n_984),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1119),
.B(n_644),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1050),
.B(n_516),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_984),
.A2(n_822),
.B(n_903),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1119),
.B(n_644),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1065),
.A2(n_1100),
.B(n_1077),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1022),
.A2(n_1081),
.A3(n_1104),
.B(n_982),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_987),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_984),
.A2(n_822),
.B(n_903),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1065),
.A2(n_1100),
.B(n_1077),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_SL g1248 ( 
.A1(n_1076),
.A2(n_1074),
.B(n_1047),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1016),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1016),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1062),
.Y(n_1251)
);

BUFx10_ASAP7_75t_L g1252 ( 
.A(n_993),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1081),
.A2(n_1109),
.B(n_980),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1065),
.A2(n_1100),
.B(n_1077),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1050),
.B(n_516),
.Y(n_1255)
);

INVxp67_ASAP7_75t_SL g1256 ( 
.A(n_1114),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_984),
.A2(n_822),
.B(n_903),
.Y(n_1257)
);

NAND3xp33_ASAP7_75t_SL g1258 ( 
.A(n_980),
.B(n_880),
.C(n_636),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1016),
.Y(n_1259)
);

OA21x2_ASAP7_75t_L g1260 ( 
.A1(n_1109),
.A2(n_1081),
.B(n_1097),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_986),
.Y(n_1261)
);

CKINVDCx14_ASAP7_75t_R g1262 ( 
.A(n_990),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1065),
.A2(n_1100),
.B(n_1077),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_984),
.A2(n_822),
.B(n_903),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_SL g1265 ( 
.A(n_999),
.B(n_940),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1022),
.A2(n_1081),
.A3(n_1104),
.B(n_982),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1065),
.A2(n_1100),
.B(n_1077),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1065),
.A2(n_1100),
.B(n_1077),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_996),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1065),
.A2(n_1100),
.B(n_1077),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_990),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_984),
.A2(n_822),
.B(n_903),
.Y(n_1272)
);

INVx5_ASAP7_75t_L g1273 ( 
.A(n_987),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_984),
.A2(n_822),
.B(n_903),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_980),
.A2(n_880),
.B1(n_894),
.B2(n_644),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1109),
.A2(n_1081),
.B(n_1097),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_984),
.A2(n_822),
.B(n_903),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_996),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1248),
.A2(n_1258),
.B(n_1126),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1137),
.B(n_1176),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1134),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1275),
.A2(n_1156),
.B(n_1225),
.C(n_1177),
.Y(n_1282)
);

AO21x2_ASAP7_75t_L g1283 ( 
.A1(n_1182),
.A2(n_1253),
.B(n_1149),
.Y(n_1283)
);

OR2x6_ASAP7_75t_L g1284 ( 
.A(n_1235),
.B(n_1169),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1134),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1184),
.A2(n_1183),
.A3(n_1148),
.B(n_1172),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1225),
.A2(n_1178),
.B(n_1193),
.C(n_1187),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1168),
.B(n_1147),
.Y(n_1288)
);

AO21x2_ASAP7_75t_L g1289 ( 
.A1(n_1182),
.A2(n_1253),
.B(n_1149),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1127),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1273),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1175),
.A2(n_1207),
.B1(n_1141),
.B2(n_1144),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1175),
.A2(n_1207),
.B1(n_1141),
.B2(n_1144),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1243),
.A2(n_1254),
.B(n_1247),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1130),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1273),
.B(n_1128),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1233),
.A2(n_1239),
.B1(n_1242),
.B2(n_1216),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1228),
.A2(n_1139),
.B(n_1277),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1145),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1238),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1138),
.A2(n_1234),
.A3(n_1257),
.B(n_1246),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1269),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1159),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1238),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1241),
.A2(n_1264),
.B(n_1274),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1154),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1261),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1155),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1251),
.B(n_1151),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1272),
.A2(n_1216),
.B(n_1160),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1205),
.A2(n_1208),
.B(n_1191),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_SL g1312 ( 
.A1(n_1208),
.A2(n_1158),
.B(n_1157),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1158),
.A2(n_1270),
.B(n_1268),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1263),
.A2(n_1267),
.B(n_1162),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1164),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1171),
.B(n_1179),
.C(n_1198),
.Y(n_1316)
);

NOR2x1_ASAP7_75t_SL g1317 ( 
.A(n_1215),
.B(n_1140),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1196),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1132),
.A2(n_1181),
.B(n_1163),
.Y(n_1319)
);

INVxp67_ASAP7_75t_SL g1320 ( 
.A(n_1213),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1230),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1125),
.A2(n_1229),
.B(n_1133),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1240),
.B(n_1255),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1152),
.A2(n_1150),
.B(n_1202),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1265),
.A2(n_1142),
.B1(n_1227),
.B2(n_1215),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1199),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_L g1327 ( 
.A(n_1153),
.B(n_1273),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1180),
.B(n_1197),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1211),
.A2(n_1276),
.B(n_1260),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1200),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1201),
.A2(n_1129),
.B(n_1212),
.Y(n_1331)
);

INVxp67_ASAP7_75t_SL g1332 ( 
.A(n_1256),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1252),
.B(n_1192),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1237),
.Y(n_1334)
);

CKINVDCx9p33_ASAP7_75t_R g1335 ( 
.A(n_1231),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1218),
.A2(n_1260),
.B(n_1276),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1195),
.A2(n_1165),
.B(n_1220),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1252),
.B(n_1204),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1128),
.B(n_1168),
.Y(n_1339)
);

NAND2x1p5_ASAP7_75t_L g1340 ( 
.A(n_1134),
.B(n_1167),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1215),
.B(n_1174),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1195),
.A2(n_1165),
.B(n_1223),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1249),
.A2(n_1250),
.B(n_1259),
.Y(n_1343)
);

AO22x2_ASAP7_75t_L g1344 ( 
.A1(n_1188),
.A2(n_1190),
.B1(n_1219),
.B2(n_1266),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1244),
.Y(n_1345)
);

BUFx2_ASAP7_75t_SL g1346 ( 
.A(n_1271),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1278),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1210),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1244),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1226),
.A2(n_1221),
.B(n_1209),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1214),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1167),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1244),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1266),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1214),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1135),
.A2(n_1170),
.B(n_1203),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_L g1357 ( 
.A(n_1131),
.B(n_1147),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1174),
.A2(n_1136),
.B1(n_1185),
.B2(n_1262),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1143),
.A2(n_1265),
.B(n_1222),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1166),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1136),
.A2(n_1245),
.B1(n_1167),
.B2(n_1206),
.Y(n_1361)
);

INVx4_ASAP7_75t_SL g1362 ( 
.A(n_1224),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1146),
.A2(n_1194),
.B(n_1173),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1186),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1210),
.A2(n_1136),
.B1(n_1245),
.B2(n_1189),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1146),
.A2(n_1194),
.B(n_1186),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1189),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1194),
.A2(n_1186),
.B(n_1146),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1217),
.A2(n_1224),
.B(n_1206),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1224),
.B(n_1217),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1189),
.B(n_1206),
.Y(n_1371)
);

CKINVDCx16_ASAP7_75t_R g1372 ( 
.A(n_1245),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1269),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1161),
.A2(n_1236),
.B(n_1232),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1253),
.A2(n_1161),
.B(n_1149),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1234),
.A2(n_1246),
.B(n_1241),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1161),
.A2(n_1236),
.B(n_1232),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1178),
.A2(n_1175),
.B1(n_980),
.B2(n_880),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1253),
.A2(n_1161),
.B(n_1149),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1161),
.A2(n_1236),
.B(n_1232),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1240),
.Y(n_1381)
);

OAI21xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1178),
.A2(n_920),
.B(n_908),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1269),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1161),
.A2(n_1236),
.B(n_1232),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1193),
.B(n_1050),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1127),
.Y(n_1386)
);

INVxp67_ASAP7_75t_SL g1387 ( 
.A(n_1251),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1127),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1137),
.B(n_1176),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1161),
.A2(n_1236),
.B(n_1232),
.Y(n_1390)
);

NAND2x1p5_ASAP7_75t_L g1391 ( 
.A(n_1273),
.B(n_999),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1127),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1161),
.A2(n_1236),
.B(n_1232),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1141),
.A2(n_1178),
.B(n_908),
.C(n_920),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1127),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1127),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1176),
.A2(n_880),
.B1(n_1078),
.B2(n_894),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1240),
.Y(n_1398)
);

NAND2x1_ASAP7_75t_L g1399 ( 
.A(n_1169),
.B(n_1235),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1127),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1161),
.A2(n_1236),
.B(n_1232),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_SL g1402 ( 
.A1(n_1208),
.A2(n_1205),
.B(n_1248),
.Y(n_1402)
);

OR2x6_ASAP7_75t_L g1403 ( 
.A(n_1235),
.B(n_1169),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1248),
.A2(n_1258),
.B(n_1126),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1258),
.A2(n_880),
.B(n_894),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1251),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_1240),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1273),
.Y(n_1408)
);

NAND2x1p5_ASAP7_75t_L g1409 ( 
.A(n_1273),
.B(n_999),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1155),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1251),
.Y(n_1411)
);

NOR2xp67_ASAP7_75t_SL g1412 ( 
.A(n_1169),
.B(n_808),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1248),
.A2(n_1258),
.B(n_1126),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1176),
.A2(n_880),
.B1(n_1078),
.B2(n_894),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1161),
.A2(n_1236),
.B(n_1232),
.Y(n_1415)
);

NAND2x1p5_ASAP7_75t_L g1416 ( 
.A(n_1273),
.B(n_999),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1385),
.B(n_1338),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1309),
.B(n_1323),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1410),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1280),
.B(n_1389),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1320),
.B(n_1328),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1394),
.A2(n_1403),
.B(n_1284),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1297),
.B(n_1398),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1394),
.A2(n_1382),
.B(n_1282),
.C(n_1287),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1305),
.A2(n_1376),
.B(n_1310),
.Y(n_1425)
);

AOI21x1_ASAP7_75t_SL g1426 ( 
.A1(n_1300),
.A2(n_1304),
.B(n_1351),
.Y(n_1426)
);

AOI21x1_ASAP7_75t_SL g1427 ( 
.A1(n_1300),
.A2(n_1351),
.B(n_1371),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1381),
.B(n_1407),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1335),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1308),
.Y(n_1430)
);

AND2x2_ASAP7_75t_SL g1431 ( 
.A(n_1292),
.B(n_1293),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1343),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1405),
.A2(n_1397),
.B(n_1414),
.C(n_1378),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_SL g1434 ( 
.A1(n_1298),
.A2(n_1378),
.B(n_1311),
.C(n_1412),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1335),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1406),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1411),
.B(n_1387),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1325),
.A2(n_1402),
.B(n_1312),
.C(n_1330),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1325),
.A2(n_1359),
.B(n_1316),
.C(n_1327),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1292),
.B(n_1293),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1284),
.A2(n_1403),
.B1(n_1399),
.B2(n_1365),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1329),
.A2(n_1337),
.B(n_1342),
.Y(n_1442)
);

O2A1O1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1327),
.A2(n_1358),
.B(n_1333),
.C(n_1284),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1403),
.A2(n_1365),
.B1(n_1333),
.B2(n_1341),
.Y(n_1444)
);

NOR2xp67_ASAP7_75t_L g1445 ( 
.A(n_1373),
.B(n_1383),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1279),
.A2(n_1413),
.B(n_1404),
.C(n_1341),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1291),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1410),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1332),
.B(n_1306),
.Y(n_1449)
);

NOR2xp67_ASAP7_75t_L g1450 ( 
.A(n_1348),
.B(n_1326),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1306),
.B(n_1307),
.Y(n_1451)
);

AND2x4_ASAP7_75t_SL g1452 ( 
.A(n_1291),
.B(n_1408),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1307),
.B(n_1326),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1344),
.B(n_1372),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1357),
.A2(n_1302),
.B1(n_1347),
.B2(n_1344),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1291),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1302),
.A2(n_1347),
.B1(n_1409),
.B2(n_1416),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1355),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1290),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1295),
.B(n_1299),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1303),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1391),
.A2(n_1416),
.B1(n_1409),
.B2(n_1334),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1315),
.B(n_1321),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1386),
.B(n_1388),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1392),
.B(n_1395),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1367),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1396),
.B(n_1400),
.Y(n_1467)
);

OR2x6_ASAP7_75t_L g1468 ( 
.A(n_1356),
.B(n_1319),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1329),
.A2(n_1342),
.B(n_1337),
.Y(n_1469)
);

INVx5_ASAP7_75t_L g1470 ( 
.A(n_1408),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1281),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1364),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1308),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1391),
.A2(n_1367),
.B1(n_1339),
.B2(n_1361),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1283),
.B(n_1289),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1368),
.A2(n_1324),
.B(n_1366),
.Y(n_1476)
);

BUFx12f_ASAP7_75t_L g1477 ( 
.A(n_1360),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1279),
.A2(n_1404),
.B(n_1413),
.C(n_1361),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1283),
.B(n_1289),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1339),
.B(n_1356),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1317),
.B(n_1370),
.Y(n_1481)
);

BUFx8_ASAP7_75t_SL g1482 ( 
.A(n_1360),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1369),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1369),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1285),
.Y(n_1485)
);

AOI221x1_ASAP7_75t_SL g1486 ( 
.A1(n_1345),
.A2(n_1353),
.B1(n_1354),
.B2(n_1349),
.C(n_1318),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1296),
.A2(n_1408),
.B1(n_1346),
.B2(n_1353),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1350),
.B(n_1352),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1350),
.B(n_1352),
.Y(n_1489)
);

A2O1A1Ixp33_ASAP7_75t_SL g1490 ( 
.A1(n_1318),
.A2(n_1345),
.B(n_1354),
.C(n_1349),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1362),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1362),
.B(n_1336),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1286),
.B(n_1301),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1296),
.A2(n_1340),
.B1(n_1379),
.B2(n_1375),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1322),
.B(n_1363),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1375),
.A2(n_1331),
.B(n_1313),
.Y(n_1496)
);

A2O1A1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1363),
.A2(n_1322),
.B(n_1384),
.C(n_1390),
.Y(n_1497)
);

BUFx4f_ASAP7_75t_L g1498 ( 
.A(n_1314),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1294),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1294),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1374),
.B(n_1377),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1380),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1380),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1384),
.A2(n_1390),
.B(n_1393),
.C(n_1401),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1393),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1415),
.B(n_1385),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1280),
.B(n_1389),
.Y(n_1507)
);

BUFx12f_ASAP7_75t_L g1508 ( 
.A(n_1360),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1341),
.B(n_1288),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_SL g1510 ( 
.A1(n_1378),
.A2(n_1034),
.B1(n_880),
.B2(n_545),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1280),
.B(n_1389),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1492),
.B(n_1506),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1479),
.B(n_1475),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1421),
.B(n_1420),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1454),
.B(n_1459),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1458),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1491),
.B(n_1488),
.Y(n_1517)
);

BUFx4f_ASAP7_75t_SL g1518 ( 
.A(n_1477),
.Y(n_1518)
);

INVxp67_ASAP7_75t_SL g1519 ( 
.A(n_1437),
.Y(n_1519)
);

CKINVDCx8_ASAP7_75t_R g1520 ( 
.A(n_1419),
.Y(n_1520)
);

INVx5_ASAP7_75t_L g1521 ( 
.A(n_1468),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1493),
.B(n_1432),
.Y(n_1522)
);

NOR2x1_ASAP7_75t_SL g1523 ( 
.A(n_1468),
.B(n_1455),
.Y(n_1523)
);

AO21x2_ASAP7_75t_L g1524 ( 
.A1(n_1504),
.A2(n_1497),
.B(n_1496),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1461),
.B(n_1460),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1507),
.B(n_1511),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1423),
.B(n_1418),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1436),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1433),
.B(n_1424),
.C(n_1434),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1443),
.B(n_1431),
.Y(n_1530)
);

CKINVDCx8_ASAP7_75t_R g1531 ( 
.A(n_1448),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1509),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1495),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1465),
.B(n_1467),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1463),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1425),
.B(n_1472),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1489),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1417),
.B(n_1425),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1425),
.B(n_1476),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1483),
.A2(n_1484),
.B(n_1503),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1480),
.B(n_1468),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1422),
.B(n_1446),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1476),
.Y(n_1543)
);

AO21x2_ASAP7_75t_L g1544 ( 
.A1(n_1490),
.A2(n_1478),
.B(n_1434),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1431),
.B(n_1449),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1464),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1453),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1486),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1424),
.A2(n_1439),
.B(n_1438),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1436),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1500),
.Y(n_1551)
);

OR2x6_ASAP7_75t_L g1552 ( 
.A(n_1441),
.B(n_1494),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1451),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1502),
.Y(n_1554)
);

AO21x2_ASAP7_75t_L g1555 ( 
.A1(n_1505),
.A2(n_1501),
.B(n_1481),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1481),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1487),
.B(n_1444),
.Y(n_1557)
);

OR2x6_ASAP7_75t_L g1558 ( 
.A(n_1499),
.B(n_1509),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1498),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1462),
.B(n_1457),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1498),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1429),
.Y(n_1562)
);

INVx5_ASAP7_75t_SL g1563 ( 
.A(n_1466),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1538),
.B(n_1442),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1538),
.B(n_1442),
.Y(n_1565)
);

AND2x4_ASAP7_75t_SL g1566 ( 
.A(n_1542),
.B(n_1466),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1529),
.A2(n_1510),
.B1(n_1440),
.B2(n_1435),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1533),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1513),
.B(n_1537),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1543),
.B(n_1469),
.Y(n_1570)
);

INVxp67_ASAP7_75t_SL g1571 ( 
.A(n_1536),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1543),
.B(n_1469),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1537),
.B(n_1428),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1533),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1529),
.A2(n_1473),
.B1(n_1430),
.B2(n_1508),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1513),
.B(n_1450),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1555),
.B(n_1426),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1522),
.B(n_1485),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1516),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1540),
.Y(n_1580)
);

AO21x2_ASAP7_75t_L g1581 ( 
.A1(n_1544),
.A2(n_1426),
.B(n_1427),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1549),
.A2(n_1474),
.B1(n_1430),
.B2(n_1466),
.C(n_1471),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1530),
.A2(n_1466),
.B1(n_1482),
.B2(n_1445),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1519),
.B(n_1456),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1554),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1554),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1522),
.B(n_1456),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1540),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1585),
.Y(n_1589)
);

OAI33xp33_ASAP7_75t_L g1590 ( 
.A1(n_1567),
.A2(n_1548),
.A3(n_1556),
.B1(n_1514),
.B2(n_1545),
.B3(n_1526),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1587),
.B(n_1555),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1585),
.Y(n_1592)
);

OA222x2_ASAP7_75t_L g1593 ( 
.A1(n_1577),
.A2(n_1542),
.B1(n_1552),
.B2(n_1557),
.C1(n_1560),
.C2(n_1558),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1567),
.A2(n_1560),
.B1(n_1557),
.B2(n_1542),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1573),
.B(n_1527),
.Y(n_1595)
);

NAND4xp25_ASAP7_75t_L g1596 ( 
.A(n_1567),
.B(n_1556),
.C(n_1548),
.D(n_1515),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1574),
.Y(n_1597)
);

OAI211xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1575),
.A2(n_1562),
.B(n_1528),
.C(n_1550),
.Y(n_1598)
);

NAND4xp25_ASAP7_75t_SL g1599 ( 
.A(n_1575),
.B(n_1515),
.C(n_1561),
.D(n_1534),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1586),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1583),
.A2(n_1542),
.B1(n_1560),
.B2(n_1557),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1586),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1576),
.B(n_1535),
.Y(n_1603)
);

AO21x2_ASAP7_75t_L g1604 ( 
.A1(n_1580),
.A2(n_1544),
.B(n_1524),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1582),
.A2(n_1542),
.B(n_1557),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1582),
.A2(n_1557),
.B1(n_1560),
.B2(n_1552),
.Y(n_1606)
);

OAI21xp33_ASAP7_75t_L g1607 ( 
.A1(n_1576),
.A2(n_1552),
.B(n_1560),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1576),
.B(n_1535),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1573),
.B(n_1520),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1566),
.A2(n_1523),
.B1(n_1552),
.B2(n_1551),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1568),
.B(n_1512),
.Y(n_1611)
);

AOI222xp33_ASAP7_75t_L g1612 ( 
.A1(n_1583),
.A2(n_1518),
.B1(n_1523),
.B2(n_1546),
.C1(n_1551),
.C2(n_1525),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1566),
.A2(n_1552),
.B1(n_1541),
.B2(n_1532),
.Y(n_1613)
);

OAI211xp5_ASAP7_75t_L g1614 ( 
.A1(n_1577),
.A2(n_1546),
.B(n_1520),
.C(n_1531),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1566),
.A2(n_1512),
.B1(n_1541),
.B2(n_1561),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1579),
.Y(n_1616)
);

NAND2xp33_ASAP7_75t_SL g1617 ( 
.A(n_1584),
.B(n_1559),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1588),
.Y(n_1618)
);

NAND3xp33_ASAP7_75t_L g1619 ( 
.A(n_1577),
.B(n_1517),
.C(n_1553),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1566),
.A2(n_1541),
.B1(n_1532),
.B2(n_1512),
.Y(n_1620)
);

NOR3xp33_ASAP7_75t_L g1621 ( 
.A(n_1584),
.B(n_1577),
.C(n_1569),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1581),
.A2(n_1563),
.B1(n_1521),
.B2(n_1559),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1587),
.B(n_1531),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1588),
.Y(n_1624)
);

NOR3xp33_ASAP7_75t_L g1625 ( 
.A(n_1569),
.B(n_1447),
.C(n_1541),
.Y(n_1625)
);

NAND3xp33_ASAP7_75t_SL g1626 ( 
.A(n_1569),
.B(n_1539),
.C(n_1547),
.Y(n_1626)
);

OAI211xp5_ASAP7_75t_L g1627 ( 
.A1(n_1587),
.A2(n_1539),
.B(n_1547),
.C(n_1553),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1578),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1616),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1594),
.B(n_1578),
.C(n_1517),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1616),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1589),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1597),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1589),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1612),
.B(n_1521),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1611),
.B(n_1621),
.Y(n_1636)
);

INVxp67_ASAP7_75t_SL g1637 ( 
.A(n_1592),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1602),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1600),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1618),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1617),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1611),
.B(n_1564),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1602),
.Y(n_1643)
);

AND2x6_ASAP7_75t_L g1644 ( 
.A(n_1615),
.B(n_1563),
.Y(n_1644)
);

INVxp67_ASAP7_75t_SL g1645 ( 
.A(n_1618),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1597),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1628),
.B(n_1571),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1624),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1624),
.Y(n_1649)
);

NAND3xp33_ASAP7_75t_SL g1650 ( 
.A(n_1605),
.B(n_1578),
.C(n_1568),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1591),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1604),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1619),
.A2(n_1572),
.B(n_1570),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1593),
.B(n_1564),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1627),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1604),
.Y(n_1656)
);

NOR2x1p5_ASAP7_75t_L g1657 ( 
.A(n_1596),
.B(n_1571),
.Y(n_1657)
);

OA21x2_ASAP7_75t_L g1658 ( 
.A1(n_1607),
.A2(n_1572),
.B(n_1570),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1604),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1641),
.B(n_1482),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1629),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1646),
.B(n_1625),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1655),
.B(n_1595),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1654),
.B(n_1610),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1629),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1655),
.B(n_1628),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1655),
.B(n_1651),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1657),
.B(n_1603),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1657),
.B(n_1636),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1654),
.B(n_1564),
.Y(n_1670)
);

NAND2x1_ASAP7_75t_L g1671 ( 
.A(n_1653),
.B(n_1564),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1633),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1657),
.B(n_1636),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1654),
.B(n_1565),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1629),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1636),
.B(n_1565),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1641),
.B(n_1565),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1631),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1647),
.B(n_1608),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1639),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1631),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1633),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1653),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1647),
.B(n_1609),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1639),
.Y(n_1685)
);

NAND2xp33_ASAP7_75t_SL g1686 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1630),
.B(n_1623),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1630),
.B(n_1590),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1651),
.B(n_1626),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1642),
.B(n_1658),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1631),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1637),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1650),
.B(n_1534),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1646),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1642),
.B(n_1622),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1632),
.Y(n_1696)
);

NAND4xp25_ASAP7_75t_SL g1697 ( 
.A(n_1635),
.B(n_1614),
.C(n_1613),
.D(n_1620),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1632),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1633),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1651),
.B(n_1617),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1637),
.B(n_1555),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1686),
.A2(n_1601),
.B1(n_1598),
.B2(n_1650),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1694),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1695),
.B(n_1646),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1696),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1694),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1666),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1664),
.B(n_1512),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1688),
.B(n_1643),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1692),
.B(n_1632),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1682),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1696),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1698),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1695),
.B(n_1658),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1698),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1682),
.B(n_1634),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1664),
.B(n_1658),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1663),
.B(n_1684),
.Y(n_1718)
);

OAI21xp33_ASAP7_75t_L g1719 ( 
.A1(n_1697),
.A2(n_1599),
.B(n_1643),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1661),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1680),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1687),
.B(n_1658),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1672),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1672),
.B(n_1634),
.Y(n_1724)
);

INVxp33_ASAP7_75t_L g1725 ( 
.A(n_1660),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1670),
.B(n_1658),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1667),
.B(n_1634),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1667),
.B(n_1658),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1670),
.B(n_1653),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1661),
.Y(n_1730)
);

AND3x2_ASAP7_75t_L g1731 ( 
.A(n_1685),
.B(n_1638),
.C(n_1568),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1699),
.B(n_1638),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1674),
.B(n_1653),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1669),
.B(n_1638),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1665),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1699),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1665),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1721),
.B(n_1707),
.Y(n_1738)
);

NOR2x1_ASAP7_75t_L g1739 ( 
.A(n_1711),
.B(n_1709),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1704),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1727),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1719),
.A2(n_1673),
.B1(n_1644),
.B2(n_1668),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1704),
.B(n_1674),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1717),
.B(n_1662),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1731),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1711),
.B(n_1689),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1708),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1727),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1717),
.B(n_1662),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1703),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1703),
.B(n_1662),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1705),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1718),
.B(n_1679),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1725),
.B(n_1702),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1702),
.B(n_1693),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1705),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1712),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1723),
.B(n_1689),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1706),
.B(n_1676),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1712),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1722),
.A2(n_1644),
.B1(n_1662),
.B2(n_1677),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1706),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1714),
.A2(n_1644),
.B1(n_1677),
.B2(n_1676),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1750),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1740),
.B(n_1734),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1739),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1754),
.B(n_1738),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1750),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1746),
.B(n_1723),
.Y(n_1769)
);

OA22x2_ASAP7_75t_L g1770 ( 
.A1(n_1742),
.A2(n_1671),
.B1(n_1736),
.B2(n_1683),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1752),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1752),
.Y(n_1772)
);

AOI21xp33_ASAP7_75t_L g1773 ( 
.A1(n_1755),
.A2(n_1710),
.B(n_1736),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1747),
.A2(n_1743),
.B1(n_1745),
.B2(n_1744),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1756),
.Y(n_1775)
);

OAI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1745),
.A2(n_1671),
.B1(n_1728),
.B2(n_1700),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1756),
.Y(n_1777)
);

INVxp67_ASAP7_75t_SL g1778 ( 
.A(n_1762),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1743),
.A2(n_1744),
.B1(n_1749),
.B2(n_1751),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1749),
.B(n_1714),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1751),
.A2(n_1644),
.B1(n_1726),
.B2(n_1733),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1761),
.A2(n_1729),
.B1(n_1733),
.B2(n_1726),
.C(n_1700),
.Y(n_1782)
);

AOI21xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1746),
.A2(n_1710),
.B(n_1716),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1774),
.B(n_1778),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1766),
.B(n_1753),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1779),
.B(n_1759),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1768),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1769),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1764),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1767),
.B(n_1783),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1780),
.B(n_1741),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1770),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1773),
.B(n_1741),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1771),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1773),
.A2(n_1758),
.B1(n_1748),
.B2(n_1763),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1765),
.B(n_1758),
.C(n_1748),
.Y(n_1796)
);

OAI211xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1790),
.A2(n_1777),
.B(n_1772),
.C(n_1775),
.Y(n_1797)
);

OAI211xp5_ASAP7_75t_L g1798 ( 
.A1(n_1784),
.A2(n_1782),
.B(n_1781),
.C(n_1757),
.Y(n_1798)
);

NAND4xp25_ASAP7_75t_SL g1799 ( 
.A(n_1795),
.B(n_1793),
.C(n_1792),
.D(n_1788),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1795),
.A2(n_1770),
.B1(n_1776),
.B2(n_1729),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1791),
.Y(n_1801)
);

AOI322xp5_ASAP7_75t_L g1802 ( 
.A1(n_1785),
.A2(n_1690),
.A3(n_1683),
.B1(n_1716),
.B2(n_1760),
.C1(n_1757),
.C2(n_1724),
.Y(n_1802)
);

OAI31xp33_ASAP7_75t_L g1803 ( 
.A1(n_1796),
.A2(n_1716),
.A3(n_1760),
.B(n_1683),
.Y(n_1803)
);

A2O1A1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1792),
.A2(n_1716),
.B(n_1701),
.C(n_1690),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1786),
.A2(n_1644),
.B1(n_1724),
.B2(n_1713),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1787),
.A2(n_1653),
.B1(n_1732),
.B2(n_1735),
.Y(n_1806)
);

OAI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1789),
.A2(n_1732),
.B1(n_1735),
.B2(n_1737),
.C(n_1730),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1801),
.Y(n_1808)
);

AOI221x1_ASAP7_75t_SL g1809 ( 
.A1(n_1800),
.A2(n_1789),
.B1(n_1794),
.B2(n_1715),
.C(n_1713),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1799),
.A2(n_1724),
.B(n_1730),
.Y(n_1810)
);

NOR2x1p5_ASAP7_75t_L g1811 ( 
.A(n_1797),
.B(n_1715),
.Y(n_1811)
);

XNOR2xp5_ASAP7_75t_L g1812 ( 
.A(n_1798),
.B(n_1724),
.Y(n_1812)
);

AOI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1805),
.A2(n_1644),
.B1(n_1720),
.B2(n_1737),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1812),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1808),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1810),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1811),
.B(n_1803),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1809),
.B(n_1802),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1813),
.Y(n_1819)
);

AOI21xp33_ASAP7_75t_SL g1820 ( 
.A1(n_1816),
.A2(n_1807),
.B(n_1804),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1814),
.B(n_1806),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1817),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1815),
.Y(n_1823)
);

AO22x2_ASAP7_75t_L g1824 ( 
.A1(n_1818),
.A2(n_1720),
.B1(n_1691),
.B2(n_1675),
.Y(n_1824)
);

NOR2xp67_ASAP7_75t_L g1825 ( 
.A(n_1820),
.B(n_1819),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1823),
.B(n_1818),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1822),
.B(n_1821),
.Y(n_1827)
);

INVx5_ASAP7_75t_L g1828 ( 
.A(n_1826),
.Y(n_1828)
);

OAI321xp33_ASAP7_75t_L g1829 ( 
.A1(n_1828),
.A2(n_1827),
.A3(n_1825),
.B1(n_1824),
.B2(n_1701),
.C(n_1691),
.Y(n_1829)
);

NAND2x1p5_ASAP7_75t_L g1830 ( 
.A(n_1829),
.B(n_1828),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1829),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1831),
.A2(n_1681),
.B(n_1678),
.Y(n_1832)
);

OAI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1830),
.A2(n_1681),
.B(n_1678),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1833),
.A2(n_1675),
.B1(n_1656),
.B2(n_1659),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1832),
.A2(n_1653),
.B1(n_1656),
.B2(n_1470),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1834),
.A2(n_1656),
.B1(n_1659),
.B2(n_1652),
.Y(n_1836)
);

OAI21xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1836),
.A2(n_1835),
.B(n_1452),
.Y(n_1837)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1838 ( 
.A1(n_1837),
.A2(n_1645),
.B(n_1640),
.C(n_1649),
.D(n_1648),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1838),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1839),
.A2(n_1656),
.B1(n_1659),
.B2(n_1652),
.C(n_1640),
.Y(n_1840)
);

AOI211xp5_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_1652),
.B(n_1659),
.C(n_1447),
.Y(n_1841)
);


endmodule