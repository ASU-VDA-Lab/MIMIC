module real_jpeg_7094_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_1),
.A2(n_244),
.B1(n_245),
.B2(n_248),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_1),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_2),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_3),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_3),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_3),
.A2(n_75),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_4),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_4),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_5),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_5),
.A2(n_108),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_5),
.A2(n_108),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_5),
.A2(n_108),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_6),
.A2(n_59),
.B1(n_64),
.B2(n_66),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_6),
.A2(n_66),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_7),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_7),
.Y(n_242)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_9),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_9),
.Y(n_140)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_11),
.A2(n_43),
.B1(n_181),
.B2(n_182),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_11),
.B(n_291),
.C(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_11),
.B(n_91),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_11),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_11),
.B(n_238),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_11),
.B(n_26),
.Y(n_351)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_12),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_12),
.Y(n_137)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_12),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_12),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_13),
.A2(n_105),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_13),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_13),
.A2(n_112),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_13),
.A2(n_112),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_13),
.A2(n_64),
.B1(n_112),
.B2(n_303),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_14),
.A2(n_172),
.B1(n_175),
.B2(n_178),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_14),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_14),
.A2(n_178),
.B1(n_219),
.B2(n_222),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_14),
.A2(n_178),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_15),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_15),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_15),
.A2(n_113),
.B1(n_122),
.B2(n_130),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_15),
.A2(n_96),
.B1(n_122),
.B2(n_182),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_15),
.A2(n_122),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_16),
.Y(n_154)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_16),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_16),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_253),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_252),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_209),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_21),
.B(n_209),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_143),
.C(n_193),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_22),
.B(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_77),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_23),
.B(n_79),
.C(n_117),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_24),
.A2(n_48),
.B1(n_49),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_24),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.A3(n_33),
.B1(n_36),
.B2(n_42),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_30),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_30),
.Y(n_221)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_32),
.A2(n_120),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_41),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g202 ( 
.A1(n_42),
.A2(n_43),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_43),
.B(n_125),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_43),
.A2(n_50),
.B(n_300),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_SL g348 ( 
.A1(n_43),
.A2(n_349),
.B(n_350),
.Y(n_348)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_57),
.B1(n_67),
.B2(n_69),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_50),
.A2(n_185),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_50),
.A2(n_296),
.B(n_300),
.Y(n_295)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_51),
.A2(n_70),
.B1(n_184),
.B2(n_191),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_51),
.A2(n_58),
.B1(n_267),
.B2(n_271),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_51),
.B(n_302),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_51),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_53),
.Y(n_272)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_53),
.Y(n_315)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_53),
.Y(n_332)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_56),
.Y(n_190)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_56),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_61),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_63),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_67),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_67),
.A2(n_319),
.B(n_324),
.Y(n_318)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_71),
.Y(n_320)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_76),
.B(n_314),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_117),
.B2(n_118),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_103),
.B(n_110),
.Y(n_79)
);

AOI22x1_ASAP7_75t_L g215 ( 
.A1(n_80),
.A2(n_91),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_80),
.B(n_216),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_80),
.A2(n_110),
.B(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_81),
.A2(n_104),
.B1(n_116),
.B2(n_208),
.Y(n_207)
);

OR2x2_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_91),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B1(n_89),
.B2(n_90),
.Y(n_82)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_83),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

AO22x2_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_94),
.Y(n_361)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_96),
.Y(n_234)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_96),
.B(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_97),
.Y(n_237)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_97),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_99),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_115),
.Y(n_222)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_115),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_116),
.A2(n_208),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_123),
.B(n_134),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_119),
.A2(n_125),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_124),
.B(n_135),
.Y(n_206)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_132),
.Y(n_125)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_127),
.Y(n_349)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_137),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_138),
.A2(n_202),
.B(n_205),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_138),
.Y(n_224)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_143),
.A2(n_144),
.B1(n_193),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_183),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_145),
.B(n_183),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_162),
.B1(n_171),
.B2(n_179),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_146),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_146),
.A2(n_162),
.B1(n_307),
.B2(n_343),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_146),
.A2(n_285),
.B(n_343),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_147),
.A2(n_180),
.B1(n_233),
.B2(n_238),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_162),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_152),
.B1(n_155),
.B2(n_159),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVx5_ASAP7_75t_SL g360 ( 
.A(n_159),
.Y(n_360)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_162),
.A2(n_171),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_162),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_162),
.A2(n_195),
.B(n_307),
.Y(n_306)
);

AOI22x1_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_167),
.B2(n_168),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_165),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_166),
.Y(n_249)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_166),
.Y(n_323)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_167),
.Y(n_293)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_186),
.Y(n_268)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_187),
.Y(n_299)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_193),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.C(n_207),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_194),
.B(n_207),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_196),
.B(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_197),
.Y(n_344)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_200),
.A2(n_201),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_231),
.B1(n_250),
.B2(n_251),
.Y(n_211)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_223),
.B1(n_229),
.B2(n_230),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

INVx6_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_237),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_242),
.Y(n_356)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_277),
.B(n_382),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_274),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_256),
.B(n_274),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.C(n_263),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_257),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_258),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_263),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.C(n_273),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_264),
.B(n_373),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_266),
.B(n_273),
.Y(n_373)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_267),
.Y(n_354)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_376),
.B(n_381),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_365),
.B(n_375),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_337),
.B(n_364),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_310),
.B(n_336),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_294),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_294),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_283),
.A2(n_286),
.B1(n_287),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_304),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_305),
.C(n_309),
.Y(n_338)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_327),
.B(n_335),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_317),
.B(n_326),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_325),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_325),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_324),
.A2(n_354),
.B(n_355),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_333),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_333),
.Y(n_335)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_339),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_352),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_346),
.B2(n_347),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_342),
.B(n_346),
.C(n_352),
.Y(n_366)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AOI32xp33_ASAP7_75t_L g357 ( 
.A1(n_351),
.A2(n_358),
.A3(n_360),
.B1(n_361),
.B2(n_362),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_357),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_357),
.Y(n_371)
);

INVx3_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_SL g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_366),
.B(n_367),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_372),
.B2(n_374),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_371),
.C(n_374),
.Y(n_377)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_372),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_377),
.B(n_378),
.Y(n_381)
);


endmodule