module fake_ibex_729_n_4732 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_810, n_768, n_338, n_173, n_696, n_796, n_797, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_217, n_324, n_391, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_232, n_380, n_749, n_281, n_559, n_425, n_4732);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_810;
input n_768;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4732;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_4557;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_4688;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_4687;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_4632;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_4607;
wire n_3750;
wire n_3838;
wire n_957;
wire n_4514;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_4550;
wire n_4668;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_2640;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_4731;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4343;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4353;
wire n_4648;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4421;
wire n_4179;
wire n_4601;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_4360;
wire n_3519;
wire n_3653;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_4585;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_4378;
wire n_850;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_4654;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_4418;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4708;
wire n_4592;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_1307;
wire n_875;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4445;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_4652;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_4673;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_4690;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_1636;
wire n_939;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3896;
wire n_3753;
wire n_2192;
wire n_4423;
wire n_4584;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_4578;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_4403;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_4002;
wire n_3631;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_1081;
wire n_4437;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_4447;
wire n_4491;
wire n_4672;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_4569;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_4723;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_4510;
wire n_2846;
wire n_2685;
wire n_3197;
wire n_3699;
wire n_1955;
wire n_3668;
wire n_4312;
wire n_4567;
wire n_917;
wire n_4556;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_4014;
wire n_3766;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_4430;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_4724;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_4721;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_4650;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_4563;
wire n_3809;
wire n_979;
wire n_4503;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4517;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_4511;
wire n_1007;
wire n_2253;
wire n_4479;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_869;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_4513;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_4667;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_4610;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_4711;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_4671;
wire n_1326;
wire n_971;
wire n_4444;
wire n_1350;
wire n_3627;
wire n_906;
wire n_4499;
wire n_2957;
wire n_4676;
wire n_2586;
wire n_3958;
wire n_1764;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_4595;
wire n_2541;
wire n_4598;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_4553;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_4533;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_4714;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4518;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_4548;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_4535;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_4505;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_4577;
wire n_2292;
wire n_3573;
wire n_4604;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2625;
wire n_1742;
wire n_2350;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4522;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_4692;
wire n_4713;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_4615;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3963;
wire n_3887;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4126;
wire n_3583;
wire n_2019;
wire n_4103;
wire n_4710;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_4680;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_4649;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_4693;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_4653;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_4568;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4549;
wire n_4573;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_4623;
wire n_1041;
wire n_4700;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_4156;
wire n_4411;
wire n_1964;
wire n_4523;
wire n_3754;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_4712;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3733;
wire n_3626;
wire n_864;
wire n_1987;
wire n_4571;
wire n_959;
wire n_1106;
wire n_1312;
wire n_4655;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_4725;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_4570;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4681;
wire n_4122;
wire n_4542;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_4572;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1985;
wire n_1140;
wire n_4375;
wire n_4501;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_2573;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2423;
wire n_4230;
wire n_859;
wire n_3849;
wire n_1109;
wire n_965;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_4558;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4504;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_4527;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_4485;
wire n_4608;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_3364;
wire n_1236;
wire n_4384;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_4537;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4407;
wire n_4323;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1890;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_4646;
wire n_1990;
wire n_1179;
wire n_907;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_4540;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_3503;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_4362;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_4706;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_4525;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_4625;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_4554;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4674;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4679;
wire n_4596;
wire n_4415;
wire n_1345;
wire n_4215;
wire n_4456;
wire n_4587;
wire n_4315;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_3470;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_4500;
wire n_4559;
wire n_998;
wire n_1395;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_4641;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4660;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_4664;
wire n_3829;
wire n_4579;
wire n_1864;
wire n_4624;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_2398;
wire n_1836;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_4709;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_4552;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1539;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4640;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4561;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_4642;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_4683;
wire n_3557;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_4614;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_4694;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_4117;
wire n_3999;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3498;
wire n_2986;
wire n_3238;
wire n_4520;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_4717;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2654;
wire n_2463;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4566;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_4719;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_4647;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4636;
wire n_4195;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1185;
wire n_1683;
wire n_4256;
wire n_3575;
wire n_4454;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_4278;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_4609;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_4685;
wire n_2948;
wire n_916;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_4716;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_4276;
wire n_831;
wire n_4612;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_3284;
wire n_2524;
wire n_3835;
wire n_1437;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_3927;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_4185;
wire n_2422;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_961;
wire n_991;
wire n_2127;
wire n_3891;
wire n_1323;
wire n_3735;
wire n_1739;
wire n_4704;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_4536;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_4633;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_4593;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_4512;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4483;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4142;
wire n_4183;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_4621;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_4066;
wire n_3990;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_4619;
wire n_4645;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3696;
wire n_3113;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_4707;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1991;
wire n_1025;
wire n_1177;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_4695;
wire n_982;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_4638;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1348;
wire n_838;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_3356;
wire n_1191;
wire n_2004;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_3899;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_4149;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_4118;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_4101;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_4637;
wire n_1396;
wire n_2916;
wire n_1923;
wire n_1224;
wire n_3206;
wire n_4021;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_3736;
wire n_1538;
wire n_3773;
wire n_2528;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_4543;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_4643;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_4603;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_3746;
wire n_2758;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_826;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_4436;
wire n_4599;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_4697;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_4538;
wire n_3096;
wire n_3333;
wire n_4509;
wire n_839;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_4730;
wire n_1415;
wire n_1238;
wire n_4616;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2251;
wire n_2012;
wire n_2963;
wire n_3512;
wire n_4720;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_4586;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_4622;
wire n_3273;
wire n_4367;
wire n_950;
wire n_3139;
wire n_2700;
wire n_1222;
wire n_4282;
wire n_4715;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_4588;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_4143;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_4698;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_3604;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3649;
wire n_833;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_4529;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2576;
wire n_2348;
wire n_2675;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4162;
wire n_4408;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_4575;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_4341;
wire n_3846;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_4620;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_4666;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_885;
wire n_4722;
wire n_1530;
wire n_4200;
wire n_3215;
wire n_3413;
wire n_877;
wire n_4580;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_4565;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_4663;
wire n_2471;
wire n_4581;
wire n_1288;
wire n_4058;
wire n_4487;
wire n_4618;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4519;
wire n_4148;
wire n_897;
wire n_1622;
wire n_2757;
wire n_4611;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_4541;
wire n_4515;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_4530;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_4463;
wire n_4591;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_4670;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1809;
wire n_1206;
wire n_855;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_4265;
wire n_3062;
wire n_4524;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2864;
wire n_2406;
wire n_1632;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4628;
wire n_4017;
wire n_1547;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1542;
wire n_3497;
wire n_4696;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3561;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_3368;
wire n_956;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4597;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_4574;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1887;
wire n_1212;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2593;
wire n_2911;
wire n_1623;
wire n_861;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_4729;
wire n_1798;
wire n_4555;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_4562;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3863;
wire n_1363;
wire n_3403;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1366;
wire n_1518;
wire n_4350;
wire n_4380;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_2653;
wire n_3173;
wire n_4345;
wire n_4281;
wire n_2411;
wire n_4478;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_4464;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_4675;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_4605;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_4546;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1635;
wire n_1572;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_3163;
wire n_2929;
wire n_2701;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_4432;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1369;
wire n_1912;
wire n_1297;
wire n_3143;
wire n_3543;
wire n_1734;
wire n_3742;
wire n_3655;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_4516;
wire n_2913;
wire n_2491;
wire n_4686;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_4682;
wire n_4528;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_4502;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_4147;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_4705;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_4471;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_4547;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_4684;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1992;
wire n_1685;
wire n_1784;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_4493;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1488;
wire n_980;
wire n_849;
wire n_1193;
wire n_2928;
wire n_3225;
wire n_2227;
wire n_2652;
wire n_3067;
wire n_1074;
wire n_3380;
wire n_3596;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_4657;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4718;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_4634;
wire n_4644;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_4412;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_4560;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_4472;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_4639;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_4635;
wire n_4521;
wire n_1230;
wire n_4459;
wire n_1516;
wire n_1027;
wire n_4551;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2618;
wire n_2357;
wire n_2855;
wire n_4448;
wire n_3938;
wire n_4354;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4401;
wire n_4532;
wire n_4727;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_4701;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4627;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_4726;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3189;
wire n_3052;
wire n_4544;
wire n_4728;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_4275;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_4589;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4617;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_4689;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_4594;
wire n_2609;
wire n_4018;
wire n_2749;
wire n_888;
wire n_2378;
wire n_3658;
wire n_1325;
wire n_4613;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_4629;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_4539;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_4702;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_4486;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_3516;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3933;
wire n_2262;
wire n_3562;
wire n_4188;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_4506;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_3691;
wire n_4452;
wire n_2544;
wire n_856;
wire n_3193;
wire n_4534;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_4590;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_4602;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_4576;
wire n_2583;
wire n_3417;
wire n_1678;
wire n_1780;
wire n_1091;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_4606;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_4508;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_4425;
wire n_4213;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_3980;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_4703;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_984;
wire n_3040;
wire n_3494;
wire n_4691;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_3180;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_203),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_482),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_588),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_62),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_767),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_673),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_212),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_662),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_514),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_438),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_529),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_679),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_75),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_544),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_503),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_820),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_638),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_633),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_678),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_458),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_502),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_709),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_469),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_624),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_750),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_323),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_663),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_333),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_658),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_794),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_644),
.Y(n_855)
);

CKINVDCx14_ASAP7_75t_R g856 ( 
.A(n_804),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_654),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_13),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_60),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_175),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_22),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_35),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_749),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_673),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_0),
.Y(n_865)
);

BUFx10_ASAP7_75t_L g866 ( 
.A(n_496),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_250),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_31),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_108),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_565),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_632),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_548),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_530),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_332),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_680),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_9),
.Y(n_876)
);

BUFx2_ASAP7_75t_R g877 ( 
.A(n_101),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_323),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_135),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_687),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_258),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_635),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_17),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_543),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_329),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_69),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_815),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_196),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_187),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_271),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_124),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_111),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_576),
.Y(n_893)
);

BUFx8_ASAP7_75t_SL g894 ( 
.A(n_816),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_810),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_604),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_48),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_685),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_329),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_316),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_597),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_176),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_679),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_497),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_375),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_496),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_239),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_297),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_330),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_737),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_560),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_622),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_675),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_29),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_119),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_18),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_569),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_266),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_666),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_615),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_210),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_237),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_734),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_556),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_422),
.Y(n_925)
);

CKINVDCx14_ASAP7_75t_R g926 ( 
.A(n_718),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_397),
.Y(n_927)
);

BUFx10_ASAP7_75t_L g928 ( 
.A(n_788),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_132),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_161),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_10),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_42),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_798),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_246),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_96),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_216),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_711),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_240),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_572),
.Y(n_939)
);

CKINVDCx14_ASAP7_75t_R g940 ( 
.A(n_119),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_690),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_224),
.Y(n_942)
);

CKINVDCx16_ASAP7_75t_R g943 ( 
.A(n_247),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_766),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_456),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_818),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_655),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_668),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_128),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_284),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_699),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_223),
.Y(n_952)
);

CKINVDCx16_ASAP7_75t_R g953 ( 
.A(n_287),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_274),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_765),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_340),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_289),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_509),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_763),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_824),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_523),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_653),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_128),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_640),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_267),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_533),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_366),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_144),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_16),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_177),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_286),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_648),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_363),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_755),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_164),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_432),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_452),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_672),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_764),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_657),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_412),
.Y(n_981)
);

BUFx10_ASAP7_75t_L g982 ( 
.A(n_486),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_160),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_49),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_91),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_629),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_192),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_464),
.Y(n_988)
);

CKINVDCx16_ASAP7_75t_R g989 ( 
.A(n_731),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_22),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_643),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_681),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_172),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_813),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_660),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_563),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_295),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_363),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_573),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_55),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_528),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_451),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_175),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_774),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_647),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_494),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_27),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_7),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_293),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_268),
.Y(n_1010)
);

BUFx10_ASAP7_75t_L g1011 ( 
.A(n_325),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_299),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_590),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_665),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_771),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_304),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_313),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_307),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_647),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_473),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_272),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_639),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_635),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_777),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_404),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_152),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_561),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_465),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_293),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_55),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_17),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_142),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_319),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_46),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_76),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_563),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_167),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_101),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_99),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_591),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_686),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_452),
.Y(n_1042)
);

BUFx10_ASAP7_75t_L g1043 ( 
.A(n_726),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_728),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_250),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_173),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_154),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_404),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_572),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_585),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_412),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_389),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_20),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_667),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_462),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_623),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_677),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_44),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_801),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_569),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_738),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_49),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_821),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_304),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_652),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_468),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_411),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_62),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_93),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_212),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_124),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_700),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_57),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_488),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_650),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_585),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_5),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_637),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_532),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_659),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_419),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_633),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_292),
.Y(n_1083)
);

CKINVDCx16_ASAP7_75t_R g1084 ( 
.A(n_393),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_321),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_206),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_817),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_653),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_10),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_137),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_252),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_417),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_414),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_651),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_520),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_485),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_423),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_594),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_547),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_205),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_108),
.Y(n_1101)
);

CKINVDCx16_ASAP7_75t_R g1102 ( 
.A(n_584),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_504),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_678),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_501),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_565),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_456),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_272),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_661),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_189),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_50),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_131),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_758),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_97),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_797),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_670),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_174),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_461),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_113),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_360),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_390),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_195),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_315),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_790),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_632),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_671),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_155),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_341),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_230),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_822),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_194),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_332),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_645),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_169),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_221),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_642),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_628),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_273),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_413),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_208),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_4),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_702),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_566),
.Y(n_1143)
);

CKINVDCx14_ASAP7_75t_R g1144 ( 
.A(n_526),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_288),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_316),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_570),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_724),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_57),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_748),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_112),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_722),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_248),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_823),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_162),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_347),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_449),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_138),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_576),
.Y(n_1159)
);

CKINVDCx16_ASAP7_75t_R g1160 ( 
.A(n_392),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_140),
.Y(n_1161)
);

CKINVDCx16_ASAP7_75t_R g1162 ( 
.A(n_253),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_13),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_803),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_177),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_725),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_328),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_706),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_609),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_205),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_627),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_775),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_641),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_495),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_93),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_535),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_455),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_497),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_789),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_181),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_139),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_302),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_213),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_422),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_545),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_259),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_515),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_161),
.Y(n_1188)
);

BUFx10_ASAP7_75t_L g1189 ( 
.A(n_327),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_403),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_129),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_607),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_469),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_529),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_568),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_26),
.Y(n_1196)
);

BUFx10_ASAP7_75t_L g1197 ( 
.A(n_570),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_462),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_47),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_83),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_371),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_405),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_665),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_587),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_574),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_528),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_483),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_683),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_203),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_495),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_802),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_229),
.Y(n_1212)
);

BUFx10_ASAP7_75t_L g1213 ( 
.A(n_403),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_418),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_545),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_514),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_423),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_357),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_312),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_90),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_421),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_745),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_773),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_697),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_254),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_660),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_814),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_646),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_430),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_620),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_550),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_407),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_300),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_61),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_94),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_393),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_453),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_656),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_167),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_657),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_793),
.Y(n_1241)
);

BUFx5_ASAP7_75t_L g1242 ( 
.A(n_509),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_433),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_380),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_209),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_266),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_714),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_594),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_631),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_688),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_539),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_623),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_712),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_303),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_217),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_436),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_631),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_193),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_257),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_106),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_636),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_99),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_90),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_735),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_634),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_676),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_245),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_446),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_591),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_141),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_310),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_50),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_134),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_781),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_491),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_649),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_302),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_135),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_477),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_105),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_279),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_759),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_259),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_174),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_146),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_753),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_140),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_490),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_58),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_52),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_536),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_102),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_282),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_146),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_599),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_674),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_717),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_805),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_46),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_592),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_716),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_136),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_110),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_517),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_23),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_76),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_386),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_378),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_157),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_424),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_664),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_9),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_184),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_705),
.Y(n_1314)
);

CKINVDCx16_ASAP7_75t_R g1315 ( 
.A(n_638),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_286),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_21),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_588),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_534),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_682),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_60),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_136),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_145),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_819),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_327),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_164),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_508),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_669),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_684),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_100),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_198),
.Y(n_1332)
);

BUFx5_ASAP7_75t_L g1333 ( 
.A(n_144),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_196),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_352),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_986),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_986),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_940),
.Y(n_1338)
);

INVxp67_ASAP7_75t_SL g1339 ( 
.A(n_837),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1192),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1192),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_874),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1242),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1232),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_894),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1232),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1242),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_928),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_833),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_833),
.Y(n_1350)
);

INVxp33_ASAP7_75t_SL g1351 ( 
.A(n_902),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1242),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_894),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1004),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_969),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_876),
.Y(n_1356)
);

INVxp33_ASAP7_75t_SL g1357 ( 
.A(n_1098),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1025),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_940),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_876),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_904),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1142),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1298),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_989),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1154),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1144),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_928),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1144),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_904),
.Y(n_1369)
);

INVxp33_ASAP7_75t_SL g1370 ( 
.A(n_1187),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1100),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_975),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1242),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1152),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1242),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_975),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_943),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1069),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1293),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_953),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1084),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1102),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1069),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_1160),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1162),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1183),
.Y(n_1386)
);

INVxp33_ASAP7_75t_L g1387 ( 
.A(n_1185),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1152),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1075),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1075),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1164),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1209),
.Y(n_1392)
);

INVxp67_ASAP7_75t_SL g1393 ( 
.A(n_1209),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1164),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1260),
.Y(n_1395)
);

CKINVDCx14_ASAP7_75t_R g1396 ( 
.A(n_856),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1315),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1260),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1267),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1267),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_827),
.Y(n_1401)
);

INVxp33_ASAP7_75t_SL g1402 ( 
.A(n_1195),
.Y(n_1402)
);

INVxp33_ASAP7_75t_L g1403 ( 
.A(n_834),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_827),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1171),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_838),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_838),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_847),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1222),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_847),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_899),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1222),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_899),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_914),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_914),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_972),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_972),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_856),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_999),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_999),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1017),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1171),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1176),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1017),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_926),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1048),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1048),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1188),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_926),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1057),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1057),
.Y(n_1431)
);

INVxp67_ASAP7_75t_SL g1432 ( 
.A(n_1099),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_825),
.Y(n_1433)
);

INVxp67_ASAP7_75t_SL g1434 ( 
.A(n_1099),
.Y(n_1434)
);

INVxp33_ASAP7_75t_L g1435 ( 
.A(n_836),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_1105),
.Y(n_1436)
);

INVxp33_ASAP7_75t_SL g1437 ( 
.A(n_826),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1105),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1108),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1335),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1108),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1173),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_866),
.Y(n_1443)
);

INVxp67_ASAP7_75t_SL g1444 ( 
.A(n_1186),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1173),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_830),
.Y(n_1446)
);

BUFx5_ASAP7_75t_L g1447 ( 
.A(n_846),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1242),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_835),
.Y(n_1449)
);

CKINVDCx16_ASAP7_75t_R g1450 ( 
.A(n_866),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_841),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_928),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1186),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_842),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1207),
.Y(n_1455)
);

CKINVDCx16_ASAP7_75t_R g1456 ( 
.A(n_866),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1207),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_1180),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1284),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1043),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1284),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_982),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_843),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_845),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1180),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_848),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1294),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1294),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1242),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_852),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1043),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1296),
.Y(n_1472)
);

INVxp67_ASAP7_75t_SL g1473 ( 
.A(n_1296),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1299),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1181),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_855),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_858),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1336),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1337),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1432),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1340),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1432),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1436),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1405),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1436),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1443),
.B(n_978),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1441),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1422),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1338),
.B(n_1007),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1365),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1387),
.B(n_982),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1365),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1441),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1443),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1365),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1473),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1346),
.B(n_1070),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1462),
.B(n_1121),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1341),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1473),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1344),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1462),
.B(n_1138),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1365),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1343),
.Y(n_1504)
);

INVx6_ASAP7_75t_L g1505 ( 
.A(n_1450),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1442),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1393),
.B(n_1320),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1348),
.B(n_1322),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1367),
.B(n_1327),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1452),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1349),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1355),
.Y(n_1512)
);

INVxp33_ASAP7_75t_L g1513 ( 
.A(n_1463),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1460),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1471),
.B(n_1024),
.Y(n_1515)
);

INVx4_ASAP7_75t_L g1516 ( 
.A(n_1448),
.Y(n_1516)
);

CKINVDCx11_ASAP7_75t_R g1517 ( 
.A(n_1445),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1350),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1342),
.B(n_1328),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1347),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1352),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1356),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1345),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1373),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1342),
.B(n_982),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1358),
.B(n_1371),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1360),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1361),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1375),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1369),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1458),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1372),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1469),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1376),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1339),
.B(n_1299),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1437),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1378),
.A2(n_1247),
.B(n_1087),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1383),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1358),
.B(n_1371),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1389),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1420),
.B(n_1332),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1390),
.Y(n_1542)
);

BUFx8_ASAP7_75t_L g1543 ( 
.A(n_1456),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1434),
.B(n_1444),
.Y(n_1544)
);

CKINVDCx16_ASAP7_75t_R g1545 ( 
.A(n_1359),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_1418),
.B(n_1043),
.Y(n_1546)
);

BUFx6f_ASAP7_75t_L g1547 ( 
.A(n_1401),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1339),
.B(n_859),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1379),
.B(n_1011),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1379),
.B(n_1302),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1396),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1404),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1392),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1395),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1403),
.B(n_861),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1423),
.B(n_1302),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1398),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1433),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1399),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1400),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1406),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1407),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_SL g1563 ( 
.A(n_1425),
.B(n_946),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1435),
.B(n_862),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1428),
.B(n_1011),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1408),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1410),
.Y(n_1567)
);

AND2x6_ASAP7_75t_L g1568 ( 
.A(n_1411),
.B(n_1024),
.Y(n_1568)
);

OAI22x1_ASAP7_75t_L g1569 ( 
.A1(n_1374),
.A2(n_877),
.B1(n_1215),
.B2(n_1181),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1413),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1414),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1415),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1402),
.B(n_1366),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1416),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1417),
.Y(n_1575)
);

BUFx8_ASAP7_75t_L g1576 ( 
.A(n_1447),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1419),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1421),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1424),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1426),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1368),
.B(n_1011),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1427),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1430),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1431),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1438),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1439),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1453),
.Y(n_1587)
);

NOR2xp67_ASAP7_75t_L g1588 ( 
.A(n_1455),
.B(n_863),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1457),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1440),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1429),
.B(n_1317),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1459),
.B(n_1311),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1446),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1461),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1467),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1468),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1472),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1474),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1447),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1353),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1447),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1465),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1447),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1475),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1447),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1354),
.Y(n_1606)
);

BUFx8_ASAP7_75t_L g1607 ( 
.A(n_1447),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1351),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1357),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1449),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1370),
.B(n_1318),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1451),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1454),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1464),
.B(n_1311),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1466),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1470),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1476),
.B(n_1120),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1477),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1364),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1388),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1362),
.Y(n_1621)
);

INVx6_ASAP7_75t_L g1622 ( 
.A(n_1377),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1391),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1394),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1380),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1409),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1363),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1412),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1381),
.A2(n_868),
.B1(n_870),
.B2(n_864),
.Y(n_1629)
);

AND2x2_ASAP7_75t_SL g1630 ( 
.A(n_1397),
.B(n_1321),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1382),
.B(n_1120),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1384),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1385),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1386),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1432),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1338),
.B(n_1325),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1345),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1336),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1443),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1432),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1345),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1348),
.B(n_937),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1432),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1348),
.B(n_941),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1336),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1443),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1387),
.B(n_1120),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1336),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1405),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1336),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1336),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1338),
.B(n_873),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1432),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_R g1654 ( 
.A(n_1396),
.B(n_829),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1432),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1338),
.B(n_884),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1338),
.B(n_849),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1443),
.B(n_1321),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1365),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1443),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1432),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1348),
.B(n_951),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1336),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1338),
.B(n_1312),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1338),
.B(n_1313),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1432),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1463),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1348),
.B(n_979),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1443),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1443),
.B(n_1329),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1338),
.B(n_1316),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1432),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1338),
.B(n_1319),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1348),
.B(n_1059),
.Y(n_1674)
);

CKINVDCx11_ASAP7_75t_R g1675 ( 
.A(n_1405),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1432),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1443),
.B(n_1329),
.Y(n_1677)
);

CKINVDCx16_ASAP7_75t_R g1678 ( 
.A(n_1450),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1343),
.A2(n_1247),
.B(n_1087),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1338),
.B(n_885),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1348),
.B(n_1061),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1336),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1405),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1443),
.B(n_1334),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1463),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1336),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1336),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1338),
.B(n_886),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1336),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1443),
.Y(n_1690)
);

NAND2xp33_ASAP7_75t_R g1691 ( 
.A(n_1345),
.B(n_888),
.Y(n_1691)
);

OA21x2_ASAP7_75t_L g1692 ( 
.A1(n_1343),
.A2(n_1113),
.B(n_1072),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1387),
.B(n_1128),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1345),
.Y(n_1694)
);

XNOR2xp5_ASAP7_75t_L g1695 ( 
.A(n_1377),
.B(n_1215),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1345),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1443),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_1405),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1512),
.Y(n_1699)
);

INVxp33_ASAP7_75t_L g1700 ( 
.A(n_1513),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1539),
.A2(n_1526),
.B1(n_1548),
.B2(n_1482),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1480),
.A2(n_844),
.B1(n_850),
.B2(n_839),
.Y(n_1702)
);

NOR2x1p5_ASAP7_75t_L g1703 ( 
.A(n_1633),
.B(n_889),
.Y(n_1703)
);

INVx3_ASAP7_75t_L g1704 ( 
.A(n_1547),
.Y(n_1704)
);

INVx8_ASAP7_75t_L g1705 ( 
.A(n_1612),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1576),
.B(n_840),
.Y(n_1706)
);

NAND2xp33_ASAP7_75t_SL g1707 ( 
.A(n_1654),
.B(n_1225),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1547),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1679),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1547),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1537),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1537),
.Y(n_1712)
);

NAND2xp33_ASAP7_75t_L g1713 ( 
.A(n_1568),
.B(n_854),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1576),
.B(n_887),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1483),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1485),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1543),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1552),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1544),
.B(n_895),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1552),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1552),
.Y(n_1721)
);

BUFx10_ASAP7_75t_L g1722 ( 
.A(n_1505),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1607),
.B(n_910),
.Y(n_1723)
);

INVx2_ASAP7_75t_SL g1724 ( 
.A(n_1505),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1487),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1493),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1496),
.Y(n_1727)
);

INVx4_ASAP7_75t_L g1728 ( 
.A(n_1615),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1500),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1635),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1640),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1574),
.Y(n_1732)
);

INVx4_ASAP7_75t_L g1733 ( 
.A(n_1494),
.Y(n_1733)
);

BUFx4f_ASAP7_75t_L g1734 ( 
.A(n_1610),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1574),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1639),
.B(n_960),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1491),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1607),
.B(n_933),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1574),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1643),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1577),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_SL g1742 ( 
.A(n_1630),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1577),
.Y(n_1743)
);

BUFx8_ASAP7_75t_SL g1744 ( 
.A(n_1484),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1577),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1653),
.A2(n_853),
.B1(n_860),
.B2(n_851),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1655),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1585),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1536),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1585),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1488),
.A2(n_1225),
.B1(n_831),
.B2(n_879),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1661),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1519),
.B(n_891),
.C(n_890),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1543),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1585),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1516),
.B(n_1535),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1561),
.Y(n_1757)
);

AND2x6_ASAP7_75t_L g1758 ( 
.A(n_1610),
.B(n_923),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1647),
.B(n_1128),
.Y(n_1759)
);

OAI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1678),
.A2(n_881),
.B1(n_897),
.B2(n_867),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_SL g1761 ( 
.A(n_1558),
.B(n_950),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_1693),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1566),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1535),
.B(n_944),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1666),
.B(n_1672),
.Y(n_1765)
);

BUFx3_ASAP7_75t_L g1766 ( 
.A(n_1612),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1571),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1676),
.Y(n_1768)
);

AND2x6_ASAP7_75t_L g1769 ( 
.A(n_1610),
.B(n_923),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1575),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1658),
.Y(n_1771)
);

INVx2_ASAP7_75t_SL g1772 ( 
.A(n_1549),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1586),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_SL g1774 ( 
.A1(n_1525),
.A2(n_1085),
.B1(n_1094),
.B2(n_1027),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1555),
.B(n_896),
.C(n_892),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1565),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1598),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1578),
.Y(n_1778)
);

CKINVDCx16_ASAP7_75t_R g1779 ( 
.A(n_1545),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1550),
.B(n_955),
.Y(n_1780)
);

BUFx6f_ASAP7_75t_L g1781 ( 
.A(n_1692),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1541),
.B(n_974),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1562),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1658),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1692),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1567),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1507),
.B(n_994),
.Y(n_1787)
);

CKINVDCx6p67_ASAP7_75t_R g1788 ( 
.A(n_1517),
.Y(n_1788)
);

OR2x6_ASAP7_75t_L g1789 ( 
.A(n_1622),
.B(n_1334),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1550),
.B(n_1015),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1570),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1564),
.B(n_1044),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1660),
.B(n_1063),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1667),
.B(n_857),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1521),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1572),
.Y(n_1796)
);

BUFx6f_ASAP7_75t_L g1797 ( 
.A(n_1521),
.Y(n_1797)
);

CKINVDCx20_ASAP7_75t_R g1798 ( 
.A(n_1675),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1579),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1497),
.B(n_1115),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1669),
.B(n_1124),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1506),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1510),
.B(n_1130),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1690),
.B(n_1150),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1580),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1670),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1670),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1582),
.Y(n_1808)
);

BUFx10_ASAP7_75t_L g1809 ( 
.A(n_1573),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1583),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1584),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1587),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1685),
.B(n_1128),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1677),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1591),
.B(n_1616),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1697),
.B(n_1636),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1589),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1594),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1595),
.Y(n_1819)
);

NAND2xp33_ASAP7_75t_SL g1820 ( 
.A(n_1613),
.B(n_903),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1646),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1677),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1596),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1597),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1684),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1684),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1554),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1522),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_L g1829 ( 
.A(n_1611),
.B(n_909),
.C(n_908),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1530),
.Y(n_1830)
);

NAND3xp33_ASAP7_75t_L g1831 ( 
.A(n_1652),
.B(n_915),
.C(n_913),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_R g1832 ( 
.A(n_1523),
.B(n_1310),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1559),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1532),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1557),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1521),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1657),
.B(n_1166),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1524),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1524),
.Y(n_1839)
);

NAND2xp33_ASAP7_75t_SL g1840 ( 
.A(n_1613),
.B(n_1307),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1524),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1478),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1479),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1481),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1499),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1618),
.B(n_1211),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1486),
.B(n_1227),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1527),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1638),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1645),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1648),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1656),
.B(n_1241),
.Y(n_1852)
);

NAND2xp33_ASAP7_75t_L g1853 ( 
.A(n_1568),
.B(n_1253),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1592),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1650),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_L g1856 ( 
.A(n_1664),
.B(n_921),
.C(n_919),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1651),
.Y(n_1857)
);

INVxp33_ASAP7_75t_L g1858 ( 
.A(n_1620),
.Y(n_1858)
);

BUFx4f_ASAP7_75t_L g1859 ( 
.A(n_1613),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1592),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1590),
.Y(n_1861)
);

OAI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1608),
.A2(n_945),
.B1(n_952),
.B2(n_916),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1665),
.B(n_1264),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1663),
.Y(n_1864)
);

BUFx3_ASAP7_75t_L g1865 ( 
.A(n_1551),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1486),
.B(n_1274),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1671),
.B(n_1282),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1682),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1556),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1540),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1581),
.B(n_1286),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1686),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1498),
.B(n_1301),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1617),
.B(n_1314),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1673),
.B(n_1680),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1531),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1502),
.B(n_1333),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1687),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1689),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1511),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1688),
.B(n_1148),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1518),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1528),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1533),
.Y(n_1884)
);

BUFx8_ASAP7_75t_SL g1885 ( 
.A(n_1602),
.Y(n_1885)
);

BUFx6f_ASAP7_75t_L g1886 ( 
.A(n_1553),
.Y(n_1886)
);

CKINVDCx16_ASAP7_75t_R g1887 ( 
.A(n_1604),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1533),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1534),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1538),
.Y(n_1890)
);

INVx4_ASAP7_75t_L g1891 ( 
.A(n_1568),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1542),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1508),
.B(n_1509),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1560),
.Y(n_1894)
);

BUFx6f_ASAP7_75t_L g1895 ( 
.A(n_1490),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1501),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1614),
.B(n_1168),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_SL g1898 ( 
.A(n_1632),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1504),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1588),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1520),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1529),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1515),
.B(n_1333),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1489),
.B(n_1172),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1601),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1599),
.Y(n_1906)
);

INVx3_ASAP7_75t_L g1907 ( 
.A(n_1514),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1614),
.A2(n_1556),
.B1(n_1609),
.B2(n_1642),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1546),
.B(n_1563),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1644),
.B(n_1333),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1603),
.Y(n_1911)
);

BUFx4f_ASAP7_75t_L g1912 ( 
.A(n_1551),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1662),
.B(n_1179),
.Y(n_1913)
);

BUFx10_ASAP7_75t_L g1914 ( 
.A(n_1600),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1668),
.B(n_1333),
.Y(n_1915)
);

CKINVDCx6p67_ASAP7_75t_R g1916 ( 
.A(n_1569),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1674),
.B(n_1223),
.Y(n_1917)
);

NOR3xp33_ASAP7_75t_L g1918 ( 
.A(n_1625),
.B(n_882),
.C(n_865),
.Y(n_1918)
);

AO22x2_ASAP7_75t_L g1919 ( 
.A1(n_1634),
.A2(n_1631),
.B1(n_1624),
.B2(n_1626),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1619),
.B(n_922),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1605),
.Y(n_1921)
);

NAND3xp33_ASAP7_75t_L g1922 ( 
.A(n_1681),
.B(n_1629),
.C(n_1623),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1593),
.B(n_828),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1621),
.B(n_1333),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_L g1925 ( 
.A(n_1490),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_1490),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1606),
.B(n_1695),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1492),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1637),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1621),
.A2(n_871),
.B1(n_872),
.B2(n_869),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1492),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1492),
.Y(n_1932)
);

INVx2_ASAP7_75t_SL g1933 ( 
.A(n_1622),
.Y(n_1933)
);

NAND3xp33_ASAP7_75t_L g1934 ( 
.A(n_1691),
.B(n_925),
.C(n_924),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_SL g1935 ( 
.A1(n_1628),
.A2(n_1331),
.B1(n_1037),
.B2(n_983),
.Y(n_1935)
);

INVx1_ASAP7_75t_SL g1936 ( 
.A(n_1649),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1495),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1621),
.B(n_828),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1627),
.B(n_828),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1641),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1628),
.B(n_927),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1495),
.Y(n_1942)
);

BUFx4f_ASAP7_75t_L g1943 ( 
.A(n_1627),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1627),
.B(n_828),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1495),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1683),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1694),
.B(n_930),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1503),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1503),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1696),
.B(n_929),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1698),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1503),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1659),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1659),
.Y(n_1954)
);

BUFx8_ASAP7_75t_SL g1955 ( 
.A(n_1659),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1547),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1505),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1547),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1576),
.B(n_832),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1679),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1576),
.B(n_832),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1512),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1480),
.Y(n_1963)
);

NAND3xp33_ASAP7_75t_L g1964 ( 
.A(n_1519),
.B(n_934),
.C(n_932),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1494),
.B(n_936),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1547),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1543),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1480),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_SL g1969 ( 
.A(n_1536),
.B(n_961),
.Y(n_1969)
);

AOI22xp33_ASAP7_75t_SL g1970 ( 
.A1(n_1512),
.A2(n_1228),
.B1(n_1082),
.B2(n_1005),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1547),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1547),
.Y(n_1972)
);

AOI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1526),
.A2(n_956),
.B1(n_958),
.B2(n_948),
.Y(n_1973)
);

INVx3_ASAP7_75t_L g1974 ( 
.A(n_1547),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1547),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1512),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1547),
.Y(n_1977)
);

INVx3_ASAP7_75t_L g1978 ( 
.A(n_1547),
.Y(n_1978)
);

OR2x6_ASAP7_75t_L g1979 ( 
.A(n_1505),
.B(n_1323),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1547),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1480),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1547),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1547),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1505),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1576),
.B(n_832),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1480),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1544),
.B(n_1333),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1480),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1547),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1480),
.Y(n_1990)
);

AOI21x1_ASAP7_75t_L g1991 ( 
.A1(n_1599),
.A2(n_1304),
.B(n_1300),
.Y(n_1991)
);

BUFx10_ASAP7_75t_L g1992 ( 
.A(n_1505),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1480),
.Y(n_1993)
);

INVx2_ASAP7_75t_SL g1994 ( 
.A(n_1512),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1679),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1679),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1547),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1994),
.B(n_963),
.Y(n_1998)
);

AOI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1772),
.A2(n_1875),
.B1(n_1701),
.B2(n_1716),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1765),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1715),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1725),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1699),
.A2(n_967),
.B1(n_970),
.B2(n_964),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_L g2004 ( 
.A(n_1722),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1726),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1976),
.B(n_1163),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1892),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1727),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1892),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1729),
.B(n_973),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_1728),
.B(n_875),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1892),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1728),
.B(n_1962),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1730),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1731),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1740),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1747),
.B(n_976),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1700),
.B(n_988),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1752),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1768),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1963),
.Y(n_2021)
);

INVxp33_ASAP7_75t_L g2022 ( 
.A(n_1832),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1858),
.B(n_1065),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1737),
.B(n_878),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1968),
.Y(n_2025)
);

BUFx3_ASAP7_75t_L g2026 ( 
.A(n_1754),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1981),
.B(n_977),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1986),
.Y(n_2028)
);

INVx2_ASAP7_75t_SL g2029 ( 
.A(n_1722),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1749),
.B(n_1163),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1861),
.B(n_1163),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1762),
.B(n_1907),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1992),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1988),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1990),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1993),
.B(n_980),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1992),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1907),
.B(n_880),
.Y(n_2038)
);

BUFx2_ASAP7_75t_L g2039 ( 
.A(n_1979),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1821),
.B(n_883),
.Y(n_2040)
);

NAND3x1_ASAP7_75t_L g2041 ( 
.A(n_1788),
.B(n_1109),
.C(n_1096),
.Y(n_2041)
);

INVx1_ASAP7_75t_SL g2042 ( 
.A(n_1865),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1705),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1896),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1778),
.B(n_981),
.Y(n_2045)
);

BUFx6f_ASAP7_75t_L g2046 ( 
.A(n_1705),
.Y(n_2046)
);

INVx3_ASAP7_75t_L g2047 ( 
.A(n_1957),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1880),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1776),
.B(n_1122),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1778),
.B(n_1882),
.Y(n_2050)
);

INVxp67_ASAP7_75t_L g2051 ( 
.A(n_1969),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1883),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1889),
.Y(n_2053)
);

BUFx3_ASAP7_75t_L g2054 ( 
.A(n_1984),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1813),
.B(n_1141),
.Y(n_2055)
);

INVxp67_ASAP7_75t_SL g2056 ( 
.A(n_1781),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1848),
.B(n_1870),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1890),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1771),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1783),
.Y(n_2060)
);

BUFx6f_ASAP7_75t_L g2061 ( 
.A(n_1848),
.Y(n_2061)
);

INVx4_ASAP7_75t_L g2062 ( 
.A(n_1979),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1759),
.B(n_1246),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_L g2064 ( 
.A(n_1922),
.B(n_1252),
.Y(n_2064)
);

BUFx4f_ASAP7_75t_L g2065 ( 
.A(n_1916),
.Y(n_2065)
);

OR2x2_ASAP7_75t_SL g2066 ( 
.A(n_1887),
.B(n_1262),
.Y(n_2066)
);

AO21x2_ASAP7_75t_L g2067 ( 
.A1(n_1711),
.A2(n_898),
.B(n_893),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1784),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1815),
.B(n_900),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1794),
.B(n_1189),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1806),
.Y(n_2071)
);

INVx5_ASAP7_75t_L g2072 ( 
.A(n_1955),
.Y(n_2072)
);

CKINVDCx8_ASAP7_75t_R g2073 ( 
.A(n_1717),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1881),
.B(n_990),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_1950),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_1869),
.B(n_1271),
.Y(n_2076)
);

AND2x4_ASAP7_75t_L g2077 ( 
.A(n_1830),
.B(n_901),
.Y(n_2077)
);

INVx2_ASAP7_75t_SL g2078 ( 
.A(n_1912),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1807),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_1848),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_1912),
.Y(n_2081)
);

AO22x2_ASAP7_75t_L g2082 ( 
.A1(n_1936),
.A2(n_1014),
.B1(n_1088),
.B2(n_985),
.Y(n_2082)
);

AO22x2_ASAP7_75t_L g2083 ( 
.A1(n_1946),
.A2(n_1205),
.B1(n_1214),
.B2(n_1107),
.Y(n_2083)
);

INVx3_ASAP7_75t_L g2084 ( 
.A(n_1870),
.Y(n_2084)
);

INVxp67_ASAP7_75t_SL g2085 ( 
.A(n_1781),
.Y(n_2085)
);

INVx1_ASAP7_75t_SL g2086 ( 
.A(n_1789),
.Y(n_2086)
);

AO21x2_ASAP7_75t_L g2087 ( 
.A1(n_1711),
.A2(n_906),
.B(n_905),
.Y(n_2087)
);

BUFx3_ASAP7_75t_L g2088 ( 
.A(n_1967),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1870),
.Y(n_2089)
);

INVx3_ASAP7_75t_L g2090 ( 
.A(n_1886),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1814),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_1862),
.B(n_1235),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_1789),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_1904),
.A2(n_907),
.B1(n_917),
.B2(n_911),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1822),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1825),
.Y(n_2096)
);

INVx4_ASAP7_75t_L g2097 ( 
.A(n_1886),
.Y(n_2097)
);

INVx1_ASAP7_75t_SL g2098 ( 
.A(n_1744),
.Y(n_2098)
);

OR2x6_ASAP7_75t_L g2099 ( 
.A(n_1724),
.B(n_1751),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_1830),
.B(n_918),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1786),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1826),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1894),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1854),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1854),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1791),
.B(n_993),
.Y(n_2106)
);

INVx3_ASAP7_75t_L g2107 ( 
.A(n_1886),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1796),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1860),
.Y(n_2109)
);

AND2x4_ASAP7_75t_L g2110 ( 
.A(n_1835),
.B(n_920),
.Y(n_2110)
);

NAND2x1p5_ASAP7_75t_L g2111 ( 
.A(n_1734),
.B(n_1249),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1860),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_SL g2113 ( 
.A1(n_1761),
.A2(n_1197),
.B1(n_1213),
.B2(n_1189),
.Y(n_2113)
);

BUFx3_ASAP7_75t_L g2114 ( 
.A(n_1766),
.Y(n_2114)
);

AOI22xp5_ASAP7_75t_L g2115 ( 
.A1(n_1908),
.A2(n_996),
.B1(n_997),
.B2(n_995),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1799),
.Y(n_2116)
);

AND2x4_ASAP7_75t_L g2117 ( 
.A(n_1835),
.B(n_931),
.Y(n_2117)
);

INVx4_ASAP7_75t_SL g2118 ( 
.A(n_1758),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1805),
.Y(n_2119)
);

BUFx2_ASAP7_75t_L g2120 ( 
.A(n_1707),
.Y(n_2120)
);

BUFx3_ASAP7_75t_L g2121 ( 
.A(n_1798),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1808),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1810),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_1811),
.A2(n_938),
.B1(n_939),
.B2(n_935),
.Y(n_2124)
);

OAI221xp5_ASAP7_75t_L g2125 ( 
.A1(n_1973),
.A2(n_1326),
.B1(n_1280),
.B2(n_1278),
.C(n_1001),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1812),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1817),
.Y(n_2127)
);

INVx4_ASAP7_75t_L g2128 ( 
.A(n_1734),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1818),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_L g2130 ( 
.A(n_1874),
.B(n_998),
.Y(n_2130)
);

AND2x6_ASAP7_75t_L g2131 ( 
.A(n_1712),
.B(n_1781),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_1859),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1819),
.Y(n_2133)
);

INVx2_ASAP7_75t_SL g2134 ( 
.A(n_1859),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_1885),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1891),
.B(n_1000),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1823),
.B(n_1003),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1824),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1827),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1827),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1842),
.B(n_1006),
.Y(n_2141)
);

OAI21xp33_ASAP7_75t_L g2142 ( 
.A1(n_1719),
.A2(n_1290),
.B(n_1289),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_L g2143 ( 
.A(n_1785),
.Y(n_2143)
);

BUFx2_ASAP7_75t_L g2144 ( 
.A(n_1929),
.Y(n_2144)
);

BUFx4f_ASAP7_75t_L g2145 ( 
.A(n_1933),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_1733),
.B(n_942),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1906),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1774),
.B(n_1189),
.Y(n_2148)
);

INVx3_ASAP7_75t_L g2149 ( 
.A(n_1914),
.Y(n_2149)
);

AOI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_1756),
.A2(n_1919),
.B1(n_1920),
.B2(n_1897),
.Y(n_2150)
);

NOR2xp33_ASAP7_75t_L g2151 ( 
.A(n_1733),
.B(n_1008),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1906),
.Y(n_2152)
);

NAND3xp33_ASAP7_75t_L g2153 ( 
.A(n_1918),
.B(n_1013),
.C(n_1009),
.Y(n_2153)
);

A2O1A1Ixp33_ASAP7_75t_L g2154 ( 
.A1(n_1712),
.A2(n_949),
.B(n_954),
.C(n_947),
.Y(n_2154)
);

NOR2xp33_ASAP7_75t_L g2155 ( 
.A(n_1871),
.B(n_1018),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1844),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1891),
.B(n_1019),
.Y(n_2157)
);

CKINVDCx8_ASAP7_75t_R g2158 ( 
.A(n_1779),
.Y(n_2158)
);

BUFx6f_ASAP7_75t_L g2159 ( 
.A(n_1785),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1970),
.B(n_1197),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1850),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1809),
.B(n_1197),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_1831),
.B(n_957),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_1940),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_1847),
.B(n_1020),
.Y(n_2165)
);

NAND3xp33_ASAP7_75t_L g2166 ( 
.A(n_1947),
.B(n_1022),
.C(n_1021),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1851),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1864),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1872),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_1856),
.B(n_962),
.Y(n_2170)
);

INVxp67_ASAP7_75t_L g2171 ( 
.A(n_1965),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1879),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1800),
.B(n_1026),
.Y(n_2173)
);

BUFx2_ASAP7_75t_L g2174 ( 
.A(n_1758),
.Y(n_2174)
);

AOI22xp33_ASAP7_75t_L g2175 ( 
.A1(n_1764),
.A2(n_966),
.B1(n_968),
.B2(n_965),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1921),
.Y(n_2176)
);

AND2x4_ASAP7_75t_L g2177 ( 
.A(n_1706),
.B(n_971),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1843),
.Y(n_2178)
);

INVx3_ASAP7_75t_L g2179 ( 
.A(n_1914),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_SL g2180 ( 
.A1(n_1935),
.A2(n_1030),
.B1(n_1031),
.B2(n_1028),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1921),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1845),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1849),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_1943),
.Y(n_2184)
);

BUFx6f_ASAP7_75t_L g2185 ( 
.A(n_1785),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1901),
.Y(n_2186)
);

OAI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_1760),
.A2(n_1927),
.B1(n_1951),
.B2(n_1943),
.Y(n_2187)
);

INVx4_ASAP7_75t_L g2188 ( 
.A(n_1758),
.Y(n_2188)
);

BUFx4f_ASAP7_75t_L g2189 ( 
.A(n_1758),
.Y(n_2189)
);

BUFx4f_ASAP7_75t_L g2190 ( 
.A(n_1769),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_1809),
.B(n_1213),
.Y(n_2191)
);

INVx4_ASAP7_75t_L g2192 ( 
.A(n_1769),
.Y(n_2192)
);

AND2x4_ASAP7_75t_L g2193 ( 
.A(n_1714),
.B(n_984),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_1723),
.B(n_987),
.Y(n_2194)
);

INVx4_ASAP7_75t_L g2195 ( 
.A(n_1769),
.Y(n_2195)
);

NAND3xp33_ASAP7_75t_L g2196 ( 
.A(n_1753),
.B(n_1034),
.C(n_1032),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1855),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_1787),
.B(n_1036),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_L g2199 ( 
.A(n_1816),
.B(n_1038),
.Y(n_2199)
);

AND2x6_ASAP7_75t_L g2200 ( 
.A(n_1909),
.B(n_1828),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_L g2201 ( 
.A(n_1795),
.Y(n_2201)
);

AND2x4_ASAP7_75t_L g2202 ( 
.A(n_1738),
.B(n_991),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1782),
.B(n_1039),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1852),
.B(n_1040),
.Y(n_2204)
);

INVx4_ASAP7_75t_SL g2205 ( 
.A(n_1769),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1857),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_L g2207 ( 
.A(n_1829),
.B(n_1780),
.Y(n_2207)
);

AOI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_1790),
.A2(n_1002),
.B1(n_1010),
.B2(n_992),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1863),
.B(n_1041),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1867),
.B(n_1046),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1901),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1868),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1878),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_1919),
.B(n_1213),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_1964),
.B(n_1047),
.Y(n_2215)
);

BUFx3_ASAP7_75t_L g2216 ( 
.A(n_1802),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_1742),
.A2(n_1736),
.B1(n_1941),
.B2(n_1893),
.Y(n_2217)
);

INVx4_ASAP7_75t_SL g2218 ( 
.A(n_1742),
.Y(n_2218)
);

HB1xp67_ASAP7_75t_L g2219 ( 
.A(n_1876),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_1834),
.B(n_1016),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_L g2221 ( 
.A1(n_1833),
.A2(n_1902),
.B1(n_1775),
.B2(n_1763),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1902),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1757),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1767),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_1820),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_1770),
.Y(n_2226)
);

INVxp67_ASAP7_75t_L g2227 ( 
.A(n_1793),
.Y(n_2227)
);

AO22x2_ASAP7_75t_L g2228 ( 
.A1(n_1959),
.A2(n_1023),
.B1(n_1033),
.B2(n_1029),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1702),
.B(n_1049),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1746),
.B(n_1050),
.Y(n_2230)
);

AOI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_1773),
.A2(n_1042),
.B1(n_1045),
.B2(n_1035),
.Y(n_2231)
);

BUFx2_ASAP7_75t_L g2232 ( 
.A(n_1840),
.Y(n_2232)
);

BUFx2_ASAP7_75t_L g2233 ( 
.A(n_1777),
.Y(n_2233)
);

OAI22xp33_ASAP7_75t_L g2234 ( 
.A1(n_1873),
.A2(n_1303),
.B1(n_1305),
.B2(n_1292),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_1703),
.B(n_1051),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_1803),
.B(n_1846),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_1930),
.B(n_1866),
.Y(n_2237)
);

AND2x4_ASAP7_75t_L g2238 ( 
.A(n_1923),
.B(n_1054),
.Y(n_2238)
);

HB1xp67_ASAP7_75t_L g2239 ( 
.A(n_1987),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1792),
.B(n_1052),
.Y(n_2240)
);

BUFx2_ASAP7_75t_L g2241 ( 
.A(n_1899),
.Y(n_2241)
);

AO22x2_ASAP7_75t_L g2242 ( 
.A1(n_1961),
.A2(n_1985),
.B1(n_1960),
.B2(n_1709),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1924),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_1801),
.B(n_1053),
.Y(n_2244)
);

INVx3_ASAP7_75t_L g2245 ( 
.A(n_1898),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1877),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1704),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1900),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_1934),
.B(n_1055),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_1795),
.Y(n_2250)
);

INVxp67_ASAP7_75t_L g2251 ( 
.A(n_1804),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1910),
.Y(n_2252)
);

AO22x2_ASAP7_75t_L g2253 ( 
.A1(n_1709),
.A2(n_1058),
.B1(n_1062),
.B2(n_1060),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1915),
.Y(n_2254)
);

BUFx3_ASAP7_75t_L g2255 ( 
.A(n_1952),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_1837),
.B(n_1913),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1704),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_1708),
.B(n_1056),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_1917),
.B(n_1064),
.Y(n_2259)
);

HB1xp67_ASAP7_75t_L g2260 ( 
.A(n_1898),
.Y(n_2260)
);

BUFx6f_ASAP7_75t_L g2261 ( 
.A(n_1795),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1713),
.B(n_1066),
.Y(n_2262)
);

INVx1_ASAP7_75t_SL g2263 ( 
.A(n_1903),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1991),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1960),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_1708),
.B(n_1067),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1995),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1995),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1996),
.Y(n_2269)
);

CKINVDCx20_ASAP7_75t_R g2270 ( 
.A(n_1938),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1996),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_1853),
.B(n_1068),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1939),
.Y(n_2273)
);

BUFx6f_ASAP7_75t_L g2274 ( 
.A(n_1797),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_1944),
.B(n_1743),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1743),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_1905),
.B(n_1071),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1974),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1974),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_1978),
.B(n_1074),
.Y(n_2280)
);

INVx4_ASAP7_75t_L g2281 ( 
.A(n_1797),
.Y(n_2281)
);

BUFx3_ASAP7_75t_L g2282 ( 
.A(n_1978),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1982),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_1982),
.B(n_1076),
.Y(n_2284)
);

AO22x2_ASAP7_75t_L g2285 ( 
.A1(n_1710),
.A2(n_1073),
.B1(n_1106),
.B2(n_1080),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_1797),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_1838),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1718),
.Y(n_2288)
);

OAI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_1911),
.A2(n_1111),
.B1(n_1117),
.B2(n_1110),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_1720),
.B(n_1077),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1997),
.B(n_1078),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1721),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_1838),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1732),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_1735),
.B(n_1079),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1739),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_1741),
.B(n_1081),
.Y(n_2297)
);

OAI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_1989),
.A2(n_1283),
.B1(n_1285),
.B2(n_1281),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1745),
.Y(n_2299)
);

BUFx3_ASAP7_75t_L g2300 ( 
.A(n_1748),
.Y(n_2300)
);

OAI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_1750),
.A2(n_1119),
.B1(n_1123),
.B2(n_1118),
.Y(n_2301)
);

BUFx3_ASAP7_75t_L g2302 ( 
.A(n_1755),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1956),
.Y(n_2303)
);

BUFx4f_ASAP7_75t_L g2304 ( 
.A(n_1958),
.Y(n_2304)
);

BUFx3_ASAP7_75t_L g2305 ( 
.A(n_1966),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1971),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1972),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1975),
.Y(n_2308)
);

INVx4_ASAP7_75t_L g2309 ( 
.A(n_1838),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1977),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_1980),
.B(n_1083),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_1983),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_1836),
.Y(n_2313)
);

BUFx3_ASAP7_75t_L g2314 ( 
.A(n_1884),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_1888),
.B(n_1086),
.Y(n_2315)
);

NAND2x1p5_ASAP7_75t_L g2316 ( 
.A(n_1895),
.B(n_1129),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1839),
.Y(n_2317)
);

BUFx2_ASAP7_75t_L g2318 ( 
.A(n_1841),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1937),
.Y(n_2319)
);

BUFx3_ASAP7_75t_L g2320 ( 
.A(n_1931),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_1895),
.B(n_1089),
.Y(n_2321)
);

INVxp67_ASAP7_75t_L g2322 ( 
.A(n_1895),
.Y(n_2322)
);

INVx5_ASAP7_75t_L g2323 ( 
.A(n_1925),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_1931),
.B(n_1132),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1937),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1948),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_L g2327 ( 
.A(n_1948),
.B(n_1090),
.Y(n_2327)
);

NAND3x1_ASAP7_75t_L g2328 ( 
.A(n_1953),
.B(n_1140),
.C(n_1135),
.Y(n_2328)
);

BUFx6f_ASAP7_75t_L g2329 ( 
.A(n_1925),
.Y(n_2329)
);

NAND3x1_ASAP7_75t_L g2330 ( 
.A(n_1953),
.B(n_1156),
.C(n_1145),
.Y(n_2330)
);

BUFx10_ASAP7_75t_L g2331 ( 
.A(n_1925),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_1926),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1954),
.B(n_1091),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1928),
.Y(n_2334)
);

OAI22xp33_ASAP7_75t_L g2335 ( 
.A1(n_1926),
.A2(n_1279),
.B1(n_1287),
.B2(n_1277),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_1932),
.B(n_1092),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_1942),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1945),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_1926),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_1949),
.B(n_1093),
.Y(n_2340)
);

AND2x6_ASAP7_75t_L g2341 ( 
.A(n_1754),
.B(n_959),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_1701),
.B(n_1095),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1765),
.Y(n_2343)
);

INVx5_ASAP7_75t_L g2344 ( 
.A(n_1955),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_1892),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_1892),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2000),
.B(n_1097),
.Y(n_2347)
);

BUFx2_ASAP7_75t_L g2348 ( 
.A(n_2039),
.Y(n_2348)
);

AOI22xp33_ASAP7_75t_L g2349 ( 
.A1(n_2064),
.A2(n_1103),
.B1(n_1104),
.B2(n_1101),
.Y(n_2349)
);

NOR2x2_ASAP7_75t_L g2350 ( 
.A(n_2099),
.B(n_1112),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2075),
.A2(n_1116),
.B1(n_1125),
.B2(n_1114),
.Y(n_2351)
);

INVx2_ASAP7_75t_SL g2352 ( 
.A(n_2004),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2343),
.B(n_1126),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2147),
.Y(n_2354)
);

BUFx4f_ASAP7_75t_L g2355 ( 
.A(n_2004),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_2046),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2152),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2070),
.B(n_1127),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2014),
.Y(n_2359)
);

AOI22xp33_ASAP7_75t_SL g2360 ( 
.A1(n_2082),
.A2(n_1133),
.B1(n_1137),
.B2(n_1134),
.Y(n_2360)
);

NOR3xp33_ASAP7_75t_SL g2361 ( 
.A(n_2135),
.B(n_1143),
.C(n_1139),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2044),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1999),
.B(n_1146),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_2329),
.Y(n_2364)
);

INVx2_ASAP7_75t_SL g2365 ( 
.A(n_2033),
.Y(n_2365)
);

INVx2_ASAP7_75t_SL g2366 ( 
.A(n_2033),
.Y(n_2366)
);

OAI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2176),
.A2(n_1149),
.B1(n_1151),
.B2(n_1147),
.Y(n_2367)
);

INVx1_ASAP7_75t_SL g2368 ( 
.A(n_2042),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2001),
.B(n_1153),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2048),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_2039),
.B(n_1155),
.Y(n_2371)
);

INVxp67_ASAP7_75t_SL g2372 ( 
.A(n_2239),
.Y(n_2372)
);

INVx4_ASAP7_75t_L g2373 ( 
.A(n_2046),
.Y(n_2373)
);

NOR2xp67_ASAP7_75t_L g2374 ( 
.A(n_2062),
.B(n_0),
.Y(n_2374)
);

INVx3_ASAP7_75t_L g2375 ( 
.A(n_2061),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2229),
.B(n_1157),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2002),
.B(n_2005),
.Y(n_2377)
);

AND2x4_ASAP7_75t_L g2378 ( 
.A(n_2062),
.B(n_1159),
.Y(n_2378)
);

BUFx8_ASAP7_75t_L g2379 ( 
.A(n_2121),
.Y(n_2379)
);

AOI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_2023),
.A2(n_1165),
.B1(n_1169),
.B2(n_1158),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2019),
.Y(n_2381)
);

AND2x2_ASAP7_75t_SL g2382 ( 
.A(n_2065),
.B(n_832),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2008),
.B(n_1170),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2015),
.B(n_1174),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2016),
.B(n_1175),
.Y(n_2385)
);

INVx2_ASAP7_75t_SL g2386 ( 
.A(n_2043),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2230),
.B(n_1177),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2031),
.B(n_1182),
.Y(n_2388)
);

BUFx12f_ASAP7_75t_SL g2389 ( 
.A(n_2099),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2021),
.B(n_1184),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2028),
.B(n_1190),
.Y(n_2391)
);

BUFx6f_ASAP7_75t_L g2392 ( 
.A(n_2329),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2052),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_2073),
.Y(n_2394)
);

NOR2x2_ASAP7_75t_L g2395 ( 
.A(n_2158),
.B(n_1191),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_SL g2396 ( 
.A(n_2335),
.B(n_1194),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2034),
.B(n_2035),
.Y(n_2397)
);

NOR3xp33_ASAP7_75t_SL g2398 ( 
.A(n_2187),
.B(n_1198),
.C(n_1196),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2053),
.Y(n_2399)
);

CKINVDCx11_ASAP7_75t_R g2400 ( 
.A(n_2098),
.Y(n_2400)
);

OAI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2181),
.A2(n_1200),
.B1(n_1201),
.B2(n_1199),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2058),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2020),
.B(n_1202),
.Y(n_2403)
);

INVx3_ASAP7_75t_SL g2404 ( 
.A(n_2072),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2025),
.Y(n_2405)
);

AOI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2063),
.A2(n_1206),
.B1(n_1210),
.B2(n_1203),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_SL g2407 ( 
.A(n_2144),
.B(n_1216),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_2236),
.B(n_1178),
.Y(n_2408)
);

AOI22xp33_ASAP7_75t_L g2409 ( 
.A1(n_2148),
.A2(n_1220),
.B1(n_1226),
.B2(n_1218),
.Y(n_2409)
);

AND2x4_ASAP7_75t_L g2410 ( 
.A(n_2236),
.B(n_1193),
.Y(n_2410)
);

NOR3xp33_ASAP7_75t_SL g2411 ( 
.A(n_2125),
.B(n_1236),
.C(n_1231),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2265),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2237),
.B(n_1239),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_L g2414 ( 
.A(n_2055),
.B(n_1240),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2086),
.B(n_1243),
.Y(n_2415)
);

AND2x4_ASAP7_75t_L g2416 ( 
.A(n_2078),
.B(n_1204),
.Y(n_2416)
);

INVx4_ASAP7_75t_L g2417 ( 
.A(n_2072),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2103),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_2049),
.B(n_2093),
.Y(n_2419)
);

NOR3xp33_ASAP7_75t_SL g2420 ( 
.A(n_2180),
.B(n_2153),
.C(n_2018),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2150),
.B(n_1248),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_2088),
.Y(n_2422)
);

NOR3xp33_ASAP7_75t_SL g2423 ( 
.A(n_1998),
.B(n_2166),
.C(n_2234),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2006),
.B(n_1250),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2069),
.B(n_2256),
.Y(n_2425)
);

AOI22xp33_ASAP7_75t_L g2426 ( 
.A1(n_2160),
.A2(n_1257),
.B1(n_1261),
.B2(n_1255),
.Y(n_2426)
);

INVxp67_ASAP7_75t_SL g2427 ( 
.A(n_2144),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2116),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2061),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2267),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2119),
.Y(n_2431)
);

AND2x2_ASAP7_75t_SL g2432 ( 
.A(n_2189),
.B(n_912),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2268),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2069),
.B(n_1263),
.Y(n_2434)
);

OR2x6_ASAP7_75t_L g2435 ( 
.A(n_2041),
.B(n_2081),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2123),
.Y(n_2436)
);

INVx2_ASAP7_75t_SL g2437 ( 
.A(n_2026),
.Y(n_2437)
);

AOI22xp33_ASAP7_75t_L g2438 ( 
.A1(n_2214),
.A2(n_1268),
.B1(n_1270),
.B2(n_1265),
.Y(n_2438)
);

AOI22xp33_ASAP7_75t_L g2439 ( 
.A1(n_2092),
.A2(n_1276),
.B1(n_1308),
.B2(n_1273),
.Y(n_2439)
);

NOR2x2_ASAP7_75t_L g2440 ( 
.A(n_2066),
.B(n_1),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2126),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2059),
.B(n_1208),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2138),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_2216),
.Y(n_2444)
);

AOI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_2269),
.A2(n_1224),
.B(n_959),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_R g2446 ( 
.A(n_2149),
.B(n_2),
.Y(n_2446)
);

NOR2xp33_ASAP7_75t_L g2447 ( 
.A(n_2076),
.B(n_1259),
.Y(n_2447)
);

AOI22xp33_ASAP7_75t_L g2448 ( 
.A1(n_2024),
.A2(n_1333),
.B1(n_1217),
.B2(n_1219),
.Y(n_2448)
);

HB1xp67_ASAP7_75t_L g2449 ( 
.A(n_2164),
.Y(n_2449)
);

AOI22xp33_ASAP7_75t_L g2450 ( 
.A1(n_2024),
.A2(n_1221),
.B1(n_1229),
.B2(n_1212),
.Y(n_2450)
);

INVxp67_ASAP7_75t_L g2451 ( 
.A(n_2285),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2030),
.B(n_1291),
.Y(n_2452)
);

NAND2x1p5_ASAP7_75t_L g2453 ( 
.A(n_2179),
.B(n_912),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2068),
.B(n_1295),
.Y(n_2454)
);

BUFx6f_ASAP7_75t_L g2455 ( 
.A(n_2201),
.Y(n_2455)
);

BUFx12f_ASAP7_75t_L g2456 ( 
.A(n_2072),
.Y(n_2456)
);

BUFx4f_ASAP7_75t_L g2457 ( 
.A(n_2341),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2071),
.B(n_1306),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2271),
.Y(n_2459)
);

AOI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2003),
.A2(n_1233),
.B1(n_1234),
.B2(n_1230),
.Y(n_2460)
);

BUFx6f_ASAP7_75t_L g2461 ( 
.A(n_2201),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2171),
.B(n_1330),
.Y(n_2462)
);

O2A1O1Ixp33_ASAP7_75t_L g2463 ( 
.A1(n_2154),
.A2(n_1237),
.B(n_1244),
.C(n_1238),
.Y(n_2463)
);

BUFx4f_ASAP7_75t_SL g2464 ( 
.A(n_2054),
.Y(n_2464)
);

HB1xp67_ASAP7_75t_L g2465 ( 
.A(n_2029),
.Y(n_2465)
);

BUFx2_ASAP7_75t_L g2466 ( 
.A(n_2285),
.Y(n_2466)
);

BUFx6f_ASAP7_75t_L g2467 ( 
.A(n_2250),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2060),
.Y(n_2468)
);

INVx4_ASAP7_75t_L g2469 ( 
.A(n_2344),
.Y(n_2469)
);

NAND2xp33_ASAP7_75t_SL g2470 ( 
.A(n_2188),
.B(n_912),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2101),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2079),
.B(n_1245),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2108),
.Y(n_2473)
);

AOI22xp5_ASAP7_75t_L g2474 ( 
.A1(n_2051),
.A2(n_1256),
.B1(n_1258),
.B2(n_1251),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_L g2475 ( 
.A(n_2120),
.B(n_1266),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2091),
.B(n_1269),
.Y(n_2476)
);

A2O1A1Ixp33_ASAP7_75t_L g2477 ( 
.A1(n_2252),
.A2(n_1275),
.B(n_1309),
.C(n_1288),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2095),
.B(n_1324),
.Y(n_2478)
);

BUFx3_ASAP7_75t_L g2479 ( 
.A(n_2114),
.Y(n_2479)
);

NOR2xp33_ASAP7_75t_L g2480 ( 
.A(n_2120),
.B(n_2),
.Y(n_2480)
);

NAND2x2_ASAP7_75t_L g2481 ( 
.A(n_2218),
.B(n_1224),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2122),
.Y(n_2482)
);

BUFx6f_ASAP7_75t_L g2483 ( 
.A(n_2250),
.Y(n_2483)
);

AOI22xp33_ASAP7_75t_L g2484 ( 
.A1(n_2163),
.A2(n_2170),
.B1(n_2040),
.B2(n_2233),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2127),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2080),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2096),
.B(n_912),
.Y(n_2487)
);

BUFx6f_ASAP7_75t_L g2488 ( 
.A(n_2261),
.Y(n_2488)
);

BUFx3_ASAP7_75t_L g2489 ( 
.A(n_2344),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2102),
.B(n_1012),
.Y(n_2490)
);

AND2x2_ASAP7_75t_SL g2491 ( 
.A(n_2190),
.B(n_1012),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2129),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2133),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_R g2494 ( 
.A(n_2037),
.B(n_3),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_R g2495 ( 
.A(n_2245),
.B(n_3),
.Y(n_2495)
);

BUFx3_ASAP7_75t_L g2496 ( 
.A(n_2344),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2156),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_2219),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2233),
.B(n_1012),
.Y(n_2499)
);

INVx4_ASAP7_75t_L g2500 ( 
.A(n_2080),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2161),
.Y(n_2501)
);

AND2x4_ASAP7_75t_L g2502 ( 
.A(n_2218),
.B(n_1297),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2167),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2094),
.B(n_2168),
.Y(n_2504)
);

O2A1O1Ixp33_ASAP7_75t_L g2505 ( 
.A1(n_2342),
.A2(n_1297),
.B(n_1131),
.C(n_1136),
.Y(n_2505)
);

NOR2xp33_ASAP7_75t_L g2506 ( 
.A(n_2227),
.B(n_4),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2186),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2211),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2222),
.Y(n_2509)
);

INVx3_ASAP7_75t_L g2510 ( 
.A(n_2089),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2169),
.Y(n_2511)
);

BUFx12f_ASAP7_75t_L g2512 ( 
.A(n_2341),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2139),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2140),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_2089),
.B(n_2298),
.Y(n_2515)
);

HB1xp67_ASAP7_75t_L g2516 ( 
.A(n_2241),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2172),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2226),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2178),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2207),
.B(n_1012),
.Y(n_2520)
);

INVx3_ASAP7_75t_L g2521 ( 
.A(n_2188),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2182),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2200),
.B(n_1131),
.Y(n_2523)
);

AND2x6_ASAP7_75t_SL g2524 ( 
.A(n_2235),
.B(n_5),
.Y(n_2524)
);

BUFx6f_ASAP7_75t_L g2525 ( 
.A(n_2261),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2274),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_2241),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_SL g2528 ( 
.A(n_2113),
.B(n_1131),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2162),
.B(n_2191),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2183),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_L g2531 ( 
.A(n_2251),
.B(n_6),
.Y(n_2531)
);

INVxp67_ASAP7_75t_L g2532 ( 
.A(n_2228),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2200),
.B(n_1131),
.Y(n_2533)
);

OR2x2_ASAP7_75t_L g2534 ( 
.A(n_2115),
.B(n_6),
.Y(n_2534)
);

INVxp67_ASAP7_75t_L g2535 ( 
.A(n_2228),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2197),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2206),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2128),
.B(n_1136),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_2260),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2217),
.B(n_7),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2212),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_SL g2542 ( 
.A(n_2128),
.B(n_1136),
.Y(n_2542)
);

HB1xp67_ASAP7_75t_L g2543 ( 
.A(n_2255),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2111),
.B(n_8),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2177),
.B(n_1136),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_2151),
.B(n_1161),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2213),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_SL g2548 ( 
.A(n_2192),
.B(n_1161),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2223),
.Y(n_2549)
);

AND2x4_ASAP7_75t_L g2550 ( 
.A(n_2177),
.B(n_1161),
.Y(n_2550)
);

BUFx6f_ASAP7_75t_L g2551 ( 
.A(n_2274),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2224),
.Y(n_2552)
);

NOR2xp33_ASAP7_75t_L g2553 ( 
.A(n_2022),
.B(n_8),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2263),
.B(n_1161),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2077),
.Y(n_2555)
);

AOI22xp33_ASAP7_75t_SL g2556 ( 
.A1(n_2082),
.A2(n_1167),
.B1(n_1272),
.B2(n_1254),
.Y(n_2556)
);

BUFx6f_ASAP7_75t_L g2557 ( 
.A(n_2286),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_2199),
.A2(n_1167),
.B1(n_1272),
.B2(n_1254),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2083),
.B(n_1167),
.Y(n_2559)
);

INVx2_ASAP7_75t_SL g2560 ( 
.A(n_2145),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2200),
.B(n_2010),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2104),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2083),
.B(n_2011),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2011),
.B(n_1167),
.Y(n_2564)
);

O2A1O1Ixp5_ASAP7_75t_L g2565 ( 
.A1(n_2057),
.A2(n_1154),
.B(n_1272),
.C(n_1254),
.Y(n_2565)
);

AOI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2193),
.A2(n_1254),
.B1(n_1272),
.B2(n_1154),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2077),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2100),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2105),
.Y(n_2569)
);

BUFx6f_ASAP7_75t_L g2570 ( 
.A(n_2286),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2100),
.Y(n_2571)
);

INVx5_ASAP7_75t_L g2572 ( 
.A(n_2192),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2110),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_SL g2574 ( 
.A(n_2032),
.B(n_1154),
.Y(n_2574)
);

AOI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_2193),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_2575)
);

INVx5_ASAP7_75t_L g2576 ( 
.A(n_2195),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2050),
.Y(n_2577)
);

AND2x4_ASAP7_75t_L g2578 ( 
.A(n_2194),
.B(n_2202),
.Y(n_2578)
);

HB1xp67_ASAP7_75t_L g2579 ( 
.A(n_2280),
.Y(n_2579)
);

AND2x6_ASAP7_75t_L g2580 ( 
.A(n_2143),
.B(n_11),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2017),
.B(n_12),
.Y(n_2581)
);

AND2x4_ASAP7_75t_L g2582 ( 
.A(n_2194),
.B(n_14),
.Y(n_2582)
);

INVx2_ASAP7_75t_SL g2583 ( 
.A(n_2047),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2246),
.Y(n_2584)
);

BUFx6f_ASAP7_75t_L g2585 ( 
.A(n_2287),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2067),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2027),
.B(n_15),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2036),
.B(n_15),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2087),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2109),
.Y(n_2590)
);

BUFx3_ASAP7_75t_L g2591 ( 
.A(n_2341),
.Y(n_2591)
);

INVx2_ASAP7_75t_SL g2592 ( 
.A(n_2032),
.Y(n_2592)
);

INVxp67_ASAP7_75t_L g2593 ( 
.A(n_2253),
.Y(n_2593)
);

OR2x2_ASAP7_75t_L g2594 ( 
.A(n_2074),
.B(n_16),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_2013),
.B(n_18),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2220),
.B(n_2163),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_2165),
.B(n_19),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2220),
.B(n_19),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2254),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2170),
.B(n_20),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2175),
.B(n_21),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_SL g2602 ( 
.A(n_2323),
.B(n_2195),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2208),
.B(n_23),
.Y(n_2603)
);

AND2x4_ASAP7_75t_L g2604 ( 
.A(n_2202),
.B(n_24),
.Y(n_2604)
);

AOI22xp33_ASAP7_75t_L g2605 ( 
.A1(n_2040),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_2130),
.B(n_25),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_SL g2607 ( 
.A(n_2323),
.B(n_2287),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2253),
.B(n_27),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2293),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2110),
.B(n_28),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2243),
.Y(n_2611)
);

O2A1O1Ixp33_ASAP7_75t_L g2612 ( 
.A1(n_2289),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2117),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2117),
.B(n_30),
.Y(n_2614)
);

OAI22xp5_ASAP7_75t_SL g2615 ( 
.A1(n_2270),
.A2(n_2155),
.B1(n_2232),
.B2(n_2225),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2112),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_2323),
.B(n_31),
.Y(n_2617)
);

INVx4_ASAP7_75t_L g2618 ( 
.A(n_2118),
.Y(n_2618)
);

AND2x4_ASAP7_75t_L g2619 ( 
.A(n_2248),
.B(n_32),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2324),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_2293),
.B(n_32),
.Y(n_2621)
);

AOI22xp33_ASAP7_75t_L g2622 ( 
.A1(n_2038),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2038),
.Y(n_2623)
);

INVx3_ASAP7_75t_L g2624 ( 
.A(n_2097),
.Y(n_2624)
);

BUFx2_ASAP7_75t_L g2625 ( 
.A(n_2284),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2240),
.B(n_33),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2146),
.B(n_34),
.Y(n_2627)
);

INVx1_ASAP7_75t_SL g2628 ( 
.A(n_2146),
.Y(n_2628)
);

AND3x1_ASAP7_75t_L g2629 ( 
.A(n_2184),
.B(n_36),
.C(n_37),
.Y(n_2629)
);

AND2x6_ASAP7_75t_L g2630 ( 
.A(n_2143),
.B(n_36),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_L g2631 ( 
.A(n_2198),
.B(n_37),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2331),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2173),
.B(n_38),
.Y(n_2633)
);

INVx3_ASAP7_75t_L g2634 ( 
.A(n_2331),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_2225),
.Y(n_2635)
);

AND2x4_ASAP7_75t_L g2636 ( 
.A(n_2118),
.B(n_38),
.Y(n_2636)
);

BUFx6f_ASAP7_75t_L g2637 ( 
.A(n_2159),
.Y(n_2637)
);

INVxp67_ASAP7_75t_L g2638 ( 
.A(n_2045),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2124),
.B(n_39),
.Y(n_2639)
);

AOI21xp5_ASAP7_75t_L g2640 ( 
.A1(n_2264),
.A2(n_691),
.B(n_689),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2324),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2336),
.Y(n_2642)
);

AOI22xp33_ASAP7_75t_L g2643 ( 
.A1(n_2259),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_2643)
);

BUFx6f_ASAP7_75t_L g2644 ( 
.A(n_2159),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2311),
.Y(n_2645)
);

OAI22xp5_ASAP7_75t_L g2646 ( 
.A1(n_2221),
.A2(n_2304),
.B1(n_2316),
.B2(n_2141),
.Y(n_2646)
);

NAND3xp33_ASAP7_75t_SL g2647 ( 
.A(n_2204),
.B(n_40),
.C(n_41),
.Y(n_2647)
);

AOI22xp5_ASAP7_75t_L g2648 ( 
.A1(n_2244),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2106),
.A2(n_47),
.B1(n_43),
.B2(n_45),
.Y(n_2649)
);

NOR2x2_ASAP7_75t_L g2650 ( 
.A(n_2205),
.B(n_45),
.Y(n_2650)
);

INVx1_ASAP7_75t_SL g2651 ( 
.A(n_2315),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2137),
.Y(n_2652)
);

AOI21xp33_ASAP7_75t_L g2653 ( 
.A1(n_2272),
.A2(n_48),
.B(n_51),
.Y(n_2653)
);

AND2x2_ASAP7_75t_SL g2654 ( 
.A(n_2174),
.B(n_2232),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2290),
.B(n_51),
.Y(n_2655)
);

AND2x2_ASAP7_75t_L g2656 ( 
.A(n_2295),
.B(n_52),
.Y(n_2656)
);

BUFx2_ASAP7_75t_L g2657 ( 
.A(n_2328),
.Y(n_2657)
);

AND2x4_ASAP7_75t_L g2658 ( 
.A(n_2205),
.B(n_53),
.Y(n_2658)
);

HB1xp67_ASAP7_75t_L g2659 ( 
.A(n_2297),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2231),
.B(n_53),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2301),
.Y(n_2661)
);

INVx4_ASAP7_75t_L g2662 ( 
.A(n_2131),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2238),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2209),
.B(n_54),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_2132),
.B(n_54),
.Y(n_2665)
);

AND2x4_ASAP7_75t_L g2666 ( 
.A(n_2136),
.B(n_56),
.Y(n_2666)
);

AND2x4_ASAP7_75t_L g2667 ( 
.A(n_2157),
.B(n_56),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2238),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2291),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2210),
.B(n_58),
.Y(n_2670)
);

INVx3_ASAP7_75t_L g2671 ( 
.A(n_2084),
.Y(n_2671)
);

AND3x1_ASAP7_75t_L g2672 ( 
.A(n_2134),
.B(n_59),
.C(n_61),
.Y(n_2672)
);

INVx2_ASAP7_75t_SL g2673 ( 
.A(n_2090),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2319),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2142),
.B(n_59),
.Y(n_2675)
);

AND2x4_ASAP7_75t_L g2676 ( 
.A(n_2203),
.B(n_63),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2333),
.Y(n_2677)
);

NOR2x1_ASAP7_75t_R g2678 ( 
.A(n_2174),
.B(n_63),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_SL g2679 ( 
.A(n_2185),
.B(n_64),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2249),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2277),
.B(n_64),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2215),
.B(n_65),
.Y(n_2682)
);

AOI22xp33_ASAP7_75t_L g2683 ( 
.A1(n_2196),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2330),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2262),
.B(n_66),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2326),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2327),
.B(n_67),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2258),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2325),
.Y(n_2689)
);

OR2x2_ASAP7_75t_SL g2690 ( 
.A(n_2185),
.B(n_68),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2266),
.B(n_2107),
.Y(n_2691)
);

INVx4_ASAP7_75t_L g2692 ( 
.A(n_2131),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2340),
.Y(n_2693)
);

BUFx3_ASAP7_75t_L g2694 ( 
.A(n_2282),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2288),
.Y(n_2695)
);

HB1xp67_ASAP7_75t_L g2696 ( 
.A(n_2242),
.Y(n_2696)
);

BUFx6f_ASAP7_75t_L g2697 ( 
.A(n_2131),
.Y(n_2697)
);

BUFx6f_ASAP7_75t_L g2698 ( 
.A(n_2281),
.Y(n_2698)
);

NAND2xp33_ASAP7_75t_SL g2699 ( 
.A(n_2281),
.B(n_68),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2299),
.Y(n_2700)
);

A2O1A1Ixp33_ASAP7_75t_L g2701 ( 
.A1(n_2273),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_2701)
);

OR2x2_ASAP7_75t_L g2702 ( 
.A(n_2321),
.B(n_2314),
.Y(n_2702)
);

BUFx3_ASAP7_75t_L g2703 ( 
.A(n_2320),
.Y(n_2703)
);

BUFx8_ASAP7_75t_L g2704 ( 
.A(n_2275),
.Y(n_2704)
);

AOI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_2056),
.A2(n_693),
.B(n_692),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2242),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2318),
.B(n_2309),
.Y(n_2707)
);

OR2x6_ASAP7_75t_L g2708 ( 
.A(n_2309),
.B(n_70),
.Y(n_2708)
);

INVx4_ASAP7_75t_L g2709 ( 
.A(n_2275),
.Y(n_2709)
);

INVx2_ASAP7_75t_SL g2710 ( 
.A(n_2276),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2292),
.Y(n_2711)
);

INVx3_ASAP7_75t_L g2712 ( 
.A(n_2300),
.Y(n_2712)
);

INVx2_ASAP7_75t_SL g2713 ( 
.A(n_2279),
.Y(n_2713)
);

AOI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2085),
.A2(n_695),
.B(n_694),
.Y(n_2714)
);

HB1xp67_ASAP7_75t_L g2715 ( 
.A(n_2322),
.Y(n_2715)
);

NOR2x2_ASAP7_75t_L g2716 ( 
.A(n_2247),
.B(n_71),
.Y(n_2716)
);

AOI21xp5_ASAP7_75t_L g2717 ( 
.A1(n_2007),
.A2(n_698),
.B(n_696),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2312),
.Y(n_2718)
);

NOR2xp33_ASAP7_75t_SL g2719 ( 
.A(n_2009),
.B(n_72),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2294),
.Y(n_2720)
);

NAND3xp33_ASAP7_75t_SL g2721 ( 
.A(n_2283),
.B(n_72),
.C(n_73),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2296),
.Y(n_2722)
);

AND2x6_ASAP7_75t_L g2723 ( 
.A(n_2012),
.B(n_73),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2303),
.Y(n_2724)
);

INVx1_ASAP7_75t_SL g2725 ( 
.A(n_2318),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2306),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2345),
.B(n_74),
.Y(n_2727)
);

AND2x6_ASAP7_75t_SL g2728 ( 
.A(n_2307),
.B(n_74),
.Y(n_2728)
);

BUFx2_ASAP7_75t_L g2729 ( 
.A(n_2346),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_SL g2730 ( 
.A(n_2257),
.B(n_75),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2308),
.Y(n_2731)
);

AND2x4_ASAP7_75t_L g2732 ( 
.A(n_2278),
.B(n_77),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2310),
.B(n_77),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_SL g2734 ( 
.A(n_2302),
.B(n_78),
.Y(n_2734)
);

INVx5_ASAP7_75t_L g2735 ( 
.A(n_2305),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2317),
.B(n_78),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2313),
.Y(n_2737)
);

OAI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2334),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2337),
.B(n_79),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2338),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2332),
.B(n_80),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_SL g2742 ( 
.A(n_2339),
.B(n_81),
.Y(n_2742)
);

AOI22xp33_ASAP7_75t_L g2743 ( 
.A1(n_2064),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2000),
.B(n_82),
.Y(n_2744)
);

BUFx3_ASAP7_75t_L g2745 ( 
.A(n_2046),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2000),
.Y(n_2746)
);

BUFx2_ASAP7_75t_L g2747 ( 
.A(n_2039),
.Y(n_2747)
);

BUFx6f_ASAP7_75t_L g2748 ( 
.A(n_2329),
.Y(n_2748)
);

BUFx3_ASAP7_75t_L g2749 ( 
.A(n_2046),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2147),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2075),
.B(n_84),
.Y(n_2751)
);

INVx3_ASAP7_75t_L g2752 ( 
.A(n_2061),
.Y(n_2752)
);

AOI21xp5_ASAP7_75t_L g2753 ( 
.A1(n_2265),
.A2(n_703),
.B(n_701),
.Y(n_2753)
);

NAND2x1p5_ASAP7_75t_L g2754 ( 
.A(n_2046),
.B(n_86),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2000),
.B(n_85),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2014),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2329),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2000),
.B(n_85),
.Y(n_2758)
);

AOI22xp33_ASAP7_75t_L g2759 ( 
.A1(n_2064),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2014),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2000),
.Y(n_2761)
);

BUFx3_ASAP7_75t_L g2762 ( 
.A(n_2046),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2000),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2000),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2000),
.B(n_87),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2000),
.Y(n_2766)
);

INVx2_ASAP7_75t_SL g2767 ( 
.A(n_2004),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2014),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_2135),
.Y(n_2769)
);

OR2x2_ASAP7_75t_L g2770 ( 
.A(n_2075),
.B(n_88),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2000),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2000),
.B(n_89),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2000),
.B(n_89),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2000),
.Y(n_2774)
);

NAND3xp33_ASAP7_75t_L g2775 ( 
.A(n_2171),
.B(n_91),
.C(n_92),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2000),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_2039),
.B(n_92),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2000),
.B(n_94),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2014),
.Y(n_2779)
);

AOI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2265),
.A2(n_707),
.B(n_704),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2000),
.Y(n_2781)
);

BUFx6f_ASAP7_75t_L g2782 ( 
.A(n_2329),
.Y(n_2782)
);

AND2x4_ASAP7_75t_L g2783 ( 
.A(n_2000),
.B(n_95),
.Y(n_2783)
);

XNOR2xp5_ASAP7_75t_L g2784 ( 
.A(n_2041),
.B(n_95),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_2064),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_2785)
);

INVx3_ASAP7_75t_L g2786 ( 
.A(n_2061),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_L g2787 ( 
.A(n_2075),
.B(n_98),
.Y(n_2787)
);

INVx3_ASAP7_75t_L g2788 ( 
.A(n_2061),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2075),
.B(n_100),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2000),
.Y(n_2790)
);

OR2x6_ASAP7_75t_L g2791 ( 
.A(n_2062),
.B(n_102),
.Y(n_2791)
);

BUFx3_ASAP7_75t_L g2792 ( 
.A(n_2046),
.Y(n_2792)
);

HB1xp67_ASAP7_75t_L g2793 ( 
.A(n_2042),
.Y(n_2793)
);

OR2x2_ASAP7_75t_L g2794 ( 
.A(n_2075),
.B(n_103),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_SL g2795 ( 
.A(n_2039),
.B(n_103),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2000),
.Y(n_2796)
);

INVx4_ASAP7_75t_L g2797 ( 
.A(n_2046),
.Y(n_2797)
);

INVx1_ASAP7_75t_SL g2798 ( 
.A(n_2042),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2000),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2000),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2000),
.Y(n_2801)
);

CKINVDCx5p33_ASAP7_75t_R g2802 ( 
.A(n_2135),
.Y(n_2802)
);

AND2x6_ASAP7_75t_SL g2803 ( 
.A(n_2099),
.B(n_104),
.Y(n_2803)
);

BUFx4f_ASAP7_75t_L g2804 ( 
.A(n_2004),
.Y(n_2804)
);

AND2x4_ASAP7_75t_L g2805 ( 
.A(n_2000),
.B(n_104),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2000),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2000),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2000),
.B(n_105),
.Y(n_2808)
);

AND3x1_ASAP7_75t_SL g2809 ( 
.A(n_2125),
.B(n_106),
.C(n_107),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2000),
.Y(n_2810)
);

BUFx3_ASAP7_75t_L g2811 ( 
.A(n_2046),
.Y(n_2811)
);

NAND2x1p5_ASAP7_75t_L g2812 ( 
.A(n_2046),
.B(n_109),
.Y(n_2812)
);

INVx2_ASAP7_75t_SL g2813 ( 
.A(n_2004),
.Y(n_2813)
);

BUFx2_ASAP7_75t_L g2814 ( 
.A(n_2039),
.Y(n_2814)
);

AOI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2064),
.A2(n_110),
.B1(n_107),
.B2(n_109),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2000),
.B(n_111),
.Y(n_2816)
);

INVxp67_ASAP7_75t_L g2817 ( 
.A(n_2039),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2000),
.B(n_112),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2000),
.Y(n_2819)
);

AOI22xp33_ASAP7_75t_L g2820 ( 
.A1(n_2064),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2000),
.Y(n_2821)
);

INVxp67_ASAP7_75t_SL g2822 ( 
.A(n_2000),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2039),
.B(n_114),
.Y(n_2823)
);

O2A1O1Ixp33_ASAP7_75t_L g2824 ( 
.A1(n_2154),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_2824)
);

NAND3xp33_ASAP7_75t_SL g2825 ( 
.A(n_2075),
.B(n_116),
.C(n_117),
.Y(n_2825)
);

NOR3xp33_ASAP7_75t_L g2826 ( 
.A(n_2187),
.B(n_118),
.C(n_120),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2000),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_SL g2828 ( 
.A(n_2039),
.B(n_118),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2000),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2147),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2014),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_R g2832 ( 
.A(n_2135),
.B(n_120),
.Y(n_2832)
);

BUFx8_ASAP7_75t_L g2833 ( 
.A(n_2121),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2000),
.B(n_121),
.Y(n_2834)
);

AOI22xp33_ASAP7_75t_L g2835 ( 
.A1(n_2064),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_2835)
);

INVx2_ASAP7_75t_SL g2836 ( 
.A(n_2004),
.Y(n_2836)
);

NOR3xp33_ASAP7_75t_SL g2837 ( 
.A(n_2135),
.B(n_122),
.C(n_123),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2147),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2014),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2014),
.Y(n_2840)
);

NOR2xp33_ASAP7_75t_L g2841 ( 
.A(n_2075),
.B(n_125),
.Y(n_2841)
);

NOR2x1_ASAP7_75t_L g2842 ( 
.A(n_2791),
.B(n_125),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2584),
.Y(n_2843)
);

BUFx6f_ASAP7_75t_L g2844 ( 
.A(n_2637),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_L g2845 ( 
.A(n_2578),
.B(n_126),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2746),
.Y(n_2846)
);

BUFx3_ASAP7_75t_L g2847 ( 
.A(n_2355),
.Y(n_2847)
);

BUFx2_ASAP7_75t_L g2848 ( 
.A(n_2372),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2584),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2761),
.Y(n_2850)
);

CKINVDCx6p67_ASAP7_75t_R g2851 ( 
.A(n_2404),
.Y(n_2851)
);

AND2x2_ASAP7_75t_L g2852 ( 
.A(n_2578),
.B(n_2822),
.Y(n_2852)
);

NOR2xp33_ASAP7_75t_L g2853 ( 
.A(n_2425),
.B(n_126),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2763),
.Y(n_2854)
);

BUFx3_ASAP7_75t_L g2855 ( 
.A(n_2355),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2764),
.B(n_127),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2766),
.B(n_127),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2771),
.Y(n_2858)
);

INVx4_ASAP7_75t_L g2859 ( 
.A(n_2804),
.Y(n_2859)
);

INVx3_ASAP7_75t_L g2860 ( 
.A(n_2618),
.Y(n_2860)
);

O2A1O1Ixp33_ASAP7_75t_L g2861 ( 
.A1(n_2593),
.A2(n_131),
.B(n_129),
.C(n_130),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2774),
.B(n_2776),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2781),
.B(n_130),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2790),
.Y(n_2864)
);

CKINVDCx16_ASAP7_75t_R g2865 ( 
.A(n_2446),
.Y(n_2865)
);

BUFx3_ASAP7_75t_L g2866 ( 
.A(n_2804),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2796),
.B(n_132),
.Y(n_2867)
);

AND2x4_ASAP7_75t_L g2868 ( 
.A(n_2799),
.B(n_133),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2800),
.B(n_133),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2801),
.B(n_134),
.Y(n_2870)
);

INVx4_ASAP7_75t_SL g2871 ( 
.A(n_2580),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2806),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_SL g2873 ( 
.A(n_2432),
.B(n_137),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2807),
.Y(n_2874)
);

BUFx3_ASAP7_75t_L g2875 ( 
.A(n_2464),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2810),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2819),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2821),
.B(n_138),
.Y(n_2878)
);

AOI22xp5_ASAP7_75t_L g2879 ( 
.A1(n_2466),
.A2(n_142),
.B1(n_139),
.B2(n_141),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2827),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2376),
.B(n_143),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_L g2882 ( 
.A(n_2529),
.B(n_143),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_R g2883 ( 
.A(n_2394),
.B(n_145),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2829),
.B(n_147),
.Y(n_2884)
);

OR2x6_ASAP7_75t_L g2885 ( 
.A(n_2791),
.B(n_147),
.Y(n_2885)
);

A2O1A1Ixp33_ASAP7_75t_L g2886 ( 
.A1(n_2826),
.A2(n_150),
.B(n_148),
.C(n_149),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2599),
.B(n_148),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2599),
.B(n_149),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2387),
.B(n_150),
.Y(n_2889)
);

HB1xp67_ASAP7_75t_L g2890 ( 
.A(n_2368),
.Y(n_2890)
);

AND3x1_ASAP7_75t_SL g2891 ( 
.A(n_2395),
.B(n_153),
.C(n_152),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2484),
.B(n_151),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_SL g2893 ( 
.A(n_2491),
.B(n_2382),
.Y(n_2893)
);

INVx3_ASAP7_75t_L g2894 ( 
.A(n_2618),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2504),
.B(n_151),
.Y(n_2895)
);

CKINVDCx5p33_ASAP7_75t_R g2896 ( 
.A(n_2400),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2563),
.B(n_153),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2611),
.B(n_154),
.Y(n_2898)
);

AOI221x1_ASAP7_75t_L g2899 ( 
.A1(n_2699),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.C(n_158),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2362),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2611),
.B(n_156),
.Y(n_2901)
);

O2A1O1Ixp5_ASAP7_75t_L g2902 ( 
.A1(n_2470),
.A2(n_710),
.B(n_713),
.C(n_708),
.Y(n_2902)
);

INVx4_ASAP7_75t_L g2903 ( 
.A(n_2457),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2596),
.B(n_2652),
.Y(n_2904)
);

CKINVDCx5p33_ASAP7_75t_R g2905 ( 
.A(n_2769),
.Y(n_2905)
);

BUFx3_ASAP7_75t_L g2906 ( 
.A(n_2356),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2628),
.B(n_158),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2642),
.B(n_2645),
.Y(n_2908)
);

INVx2_ASAP7_75t_SL g2909 ( 
.A(n_2745),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2370),
.B(n_159),
.Y(n_2910)
);

BUFx3_ASAP7_75t_L g2911 ( 
.A(n_2749),
.Y(n_2911)
);

INVx4_ASAP7_75t_L g2912 ( 
.A(n_2457),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2412),
.Y(n_2913)
);

AND3x2_ASAP7_75t_SL g2914 ( 
.A(n_2440),
.B(n_159),
.C(n_160),
.Y(n_2914)
);

INVx3_ASAP7_75t_L g2915 ( 
.A(n_2572),
.Y(n_2915)
);

NOR2x1p5_ASAP7_75t_L g2916 ( 
.A(n_2512),
.B(n_162),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2393),
.B(n_163),
.Y(n_2917)
);

INVx3_ASAP7_75t_L g2918 ( 
.A(n_2572),
.Y(n_2918)
);

INVx2_ASAP7_75t_SL g2919 ( 
.A(n_2762),
.Y(n_2919)
);

BUFx6f_ASAP7_75t_L g2920 ( 
.A(n_2637),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_2798),
.B(n_163),
.Y(n_2921)
);

BUFx8_ASAP7_75t_L g2922 ( 
.A(n_2456),
.Y(n_2922)
);

INVx4_ASAP7_75t_L g2923 ( 
.A(n_2708),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2399),
.Y(n_2924)
);

INVx4_ASAP7_75t_L g2925 ( 
.A(n_2708),
.Y(n_2925)
);

BUFx8_ASAP7_75t_L g2926 ( 
.A(n_2489),
.Y(n_2926)
);

NOR3xp33_ASAP7_75t_L g2927 ( 
.A(n_2360),
.B(n_165),
.C(n_166),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2402),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2430),
.Y(n_2929)
);

BUFx3_ASAP7_75t_L g2930 ( 
.A(n_2792),
.Y(n_2930)
);

AND2x4_ASAP7_75t_L g2931 ( 
.A(n_2577),
.B(n_165),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2497),
.Y(n_2932)
);

CKINVDCx20_ASAP7_75t_R g2933 ( 
.A(n_2379),
.Y(n_2933)
);

HB1xp67_ASAP7_75t_L g2934 ( 
.A(n_2793),
.Y(n_2934)
);

BUFx2_ASAP7_75t_L g2935 ( 
.A(n_2498),
.Y(n_2935)
);

AOI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_2419),
.A2(n_169),
.B1(n_166),
.B2(n_168),
.Y(n_2936)
);

AND2x4_ASAP7_75t_L g2937 ( 
.A(n_2577),
.B(n_168),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2433),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2459),
.Y(n_2939)
);

BUFx8_ASAP7_75t_L g2940 ( 
.A(n_2496),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2359),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2377),
.B(n_170),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2397),
.B(n_170),
.Y(n_2943)
);

BUFx2_ASAP7_75t_L g2944 ( 
.A(n_2427),
.Y(n_2944)
);

NAND3xp33_ASAP7_75t_L g2945 ( 
.A(n_2556),
.B(n_171),
.C(n_172),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2651),
.B(n_171),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2659),
.B(n_2501),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2503),
.B(n_173),
.Y(n_2948)
);

INVx3_ASAP7_75t_L g2949 ( 
.A(n_2572),
.Y(n_2949)
);

HB1xp67_ASAP7_75t_L g2950 ( 
.A(n_2516),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2511),
.B(n_176),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2517),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_L g2953 ( 
.A(n_2817),
.B(n_178),
.Y(n_2953)
);

NOR2xp33_ASAP7_75t_SL g2954 ( 
.A(n_2389),
.B(n_178),
.Y(n_2954)
);

HB1xp67_ASAP7_75t_L g2955 ( 
.A(n_2527),
.Y(n_2955)
);

AOI22x1_ASAP7_75t_L g2956 ( 
.A1(n_2453),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2418),
.Y(n_2957)
);

AND2x4_ASAP7_75t_L g2958 ( 
.A(n_2677),
.B(n_2669),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2428),
.Y(n_2959)
);

AND2x4_ASAP7_75t_L g2960 ( 
.A(n_2709),
.B(n_2373),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2431),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2436),
.Y(n_2962)
);

BUFx2_ASAP7_75t_L g2963 ( 
.A(n_2444),
.Y(n_2963)
);

CKINVDCx5p33_ASAP7_75t_R g2964 ( 
.A(n_2802),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2637),
.Y(n_2965)
);

CKINVDCx5p33_ASAP7_75t_R g2966 ( 
.A(n_2379),
.Y(n_2966)
);

AOI22xp33_ASAP7_75t_L g2967 ( 
.A1(n_2532),
.A2(n_182),
.B1(n_179),
.B2(n_180),
.Y(n_2967)
);

CKINVDCx14_ASAP7_75t_R g2968 ( 
.A(n_2832),
.Y(n_2968)
);

BUFx12f_ASAP7_75t_L g2969 ( 
.A(n_2833),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2441),
.Y(n_2970)
);

BUFx2_ASAP7_75t_L g2971 ( 
.A(n_2811),
.Y(n_2971)
);

BUFx6f_ASAP7_75t_L g2972 ( 
.A(n_2644),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2579),
.B(n_182),
.Y(n_2973)
);

AND2x4_ASAP7_75t_L g2974 ( 
.A(n_2709),
.B(n_183),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_SL g2975 ( 
.A(n_2654),
.B(n_183),
.Y(n_2975)
);

NOR2xp33_ASAP7_75t_L g2976 ( 
.A(n_2638),
.B(n_184),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2443),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_SL g2978 ( 
.A(n_2783),
.B(n_185),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_2644),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2381),
.Y(n_2980)
);

AND2x2_ASAP7_75t_L g2981 ( 
.A(n_2582),
.B(n_185),
.Y(n_2981)
);

CKINVDCx11_ASAP7_75t_R g2982 ( 
.A(n_2417),
.Y(n_2982)
);

CKINVDCx11_ASAP7_75t_R g2983 ( 
.A(n_2417),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2519),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2661),
.B(n_186),
.Y(n_2985)
);

AND2x4_ASAP7_75t_L g2986 ( 
.A(n_2373),
.B(n_186),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2452),
.B(n_187),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2522),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2405),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2756),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2518),
.B(n_188),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_SL g2992 ( 
.A(n_2783),
.B(n_188),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2760),
.Y(n_2993)
);

CKINVDCx5p33_ASAP7_75t_R g2994 ( 
.A(n_2833),
.Y(n_2994)
);

BUFx12f_ASAP7_75t_L g2995 ( 
.A(n_2422),
.Y(n_2995)
);

NOR2xp33_ASAP7_75t_R g2996 ( 
.A(n_2539),
.B(n_2591),
.Y(n_2996)
);

OAI21xp5_ASAP7_75t_L g2997 ( 
.A1(n_2347),
.A2(n_189),
.B(n_190),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2477),
.B(n_190),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2768),
.Y(n_2999)
);

BUFx6f_ASAP7_75t_L g3000 ( 
.A(n_2644),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2779),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2625),
.B(n_191),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2663),
.B(n_2668),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2530),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2364),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2831),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2358),
.B(n_2462),
.Y(n_3007)
);

CKINVDCx5p33_ASAP7_75t_R g3008 ( 
.A(n_2494),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2506),
.B(n_191),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2839),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2840),
.Y(n_3011)
);

INVx2_ASAP7_75t_SL g3012 ( 
.A(n_2797),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2541),
.Y(n_3013)
);

INVx6_ASAP7_75t_L g3014 ( 
.A(n_2797),
.Y(n_3014)
);

HB1xp67_ASAP7_75t_L g3015 ( 
.A(n_2543),
.Y(n_3015)
);

BUFx3_ASAP7_75t_L g3016 ( 
.A(n_2479),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2547),
.Y(n_3017)
);

BUFx4f_ASAP7_75t_SL g3018 ( 
.A(n_2469),
.Y(n_3018)
);

INVx3_ASAP7_75t_L g3019 ( 
.A(n_2576),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2513),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2531),
.B(n_192),
.Y(n_3021)
);

BUFx12f_ASAP7_75t_L g3022 ( 
.A(n_2469),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_SL g3023 ( 
.A(n_2805),
.B(n_193),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2514),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2536),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2537),
.Y(n_3026)
);

OR2x2_ASAP7_75t_L g3027 ( 
.A(n_2770),
.B(n_194),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2582),
.B(n_195),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2604),
.B(n_197),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2413),
.B(n_197),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2398),
.B(n_198),
.Y(n_3031)
);

OAI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2451),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2549),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2552),
.Y(n_3034)
);

AND2x2_ASAP7_75t_L g3035 ( 
.A(n_2604),
.B(n_199),
.Y(n_3035)
);

INVx2_ASAP7_75t_SL g3036 ( 
.A(n_2352),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2535),
.B(n_200),
.Y(n_3037)
);

BUFx3_ASAP7_75t_L g3038 ( 
.A(n_2365),
.Y(n_3038)
);

AND2x6_ASAP7_75t_L g3039 ( 
.A(n_2805),
.B(n_201),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2473),
.Y(n_3040)
);

BUFx5_ASAP7_75t_L g3041 ( 
.A(n_2580),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2450),
.B(n_202),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2447),
.B(n_202),
.Y(n_3043)
);

BUFx6f_ASAP7_75t_L g3044 ( 
.A(n_2364),
.Y(n_3044)
);

BUFx4f_ASAP7_75t_L g3045 ( 
.A(n_2580),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2507),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2508),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2388),
.B(n_204),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2492),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2493),
.Y(n_3050)
);

INVxp67_ASAP7_75t_SL g3051 ( 
.A(n_2619),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2619),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2751),
.B(n_204),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2744),
.Y(n_3054)
);

AND2x4_ASAP7_75t_L g3055 ( 
.A(n_2576),
.B(n_206),
.Y(n_3055)
);

AOI22xp33_ASAP7_75t_L g3056 ( 
.A1(n_2559),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2755),
.Y(n_3057)
);

NAND2xp33_ASAP7_75t_L g3058 ( 
.A(n_2580),
.B(n_207),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2509),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2424),
.B(n_210),
.Y(n_3060)
);

BUFx2_ASAP7_75t_L g3061 ( 
.A(n_2348),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_2789),
.B(n_211),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2758),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2765),
.Y(n_3064)
);

BUFx6f_ASAP7_75t_L g3065 ( 
.A(n_2364),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_2411),
.B(n_211),
.Y(n_3066)
);

A2O1A1Ixp33_ASAP7_75t_L g3067 ( 
.A1(n_2606),
.A2(n_215),
.B(n_213),
.C(n_214),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2623),
.B(n_214),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2354),
.Y(n_3069)
);

BUFx6f_ASAP7_75t_L g3070 ( 
.A(n_2392),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2620),
.B(n_2641),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_SL g3072 ( 
.A(n_2635),
.B(n_215),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2555),
.B(n_2567),
.Y(n_3073)
);

OAI22xp5_ASAP7_75t_L g3074 ( 
.A1(n_2690),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_3074)
);

AOI22xp5_ASAP7_75t_L g3075 ( 
.A1(n_2414),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2657),
.B(n_219),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2568),
.B(n_220),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2416),
.B(n_221),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2772),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2571),
.B(n_222),
.Y(n_3080)
);

HB1xp67_ASAP7_75t_L g3081 ( 
.A(n_2725),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2354),
.Y(n_3082)
);

OR2x2_ASAP7_75t_L g3083 ( 
.A(n_2794),
.B(n_222),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2773),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2416),
.B(n_2747),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2573),
.B(n_223),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2778),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2808),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2816),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2613),
.B(n_224),
.Y(n_3090)
);

AOI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_2540),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2818),
.Y(n_3092)
);

AND2x2_ASAP7_75t_L g3093 ( 
.A(n_2814),
.B(n_225),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2834),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2357),
.Y(n_3095)
);

CKINVDCx20_ASAP7_75t_R g3096 ( 
.A(n_2495),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2460),
.B(n_226),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2711),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2357),
.Y(n_3099)
);

NOR2x1_ASAP7_75t_L g3100 ( 
.A(n_2435),
.B(n_227),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2750),
.Y(n_3101)
);

NAND2xp33_ASAP7_75t_L g3102 ( 
.A(n_2630),
.B(n_228),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2720),
.Y(n_3103)
);

AND2x2_ASAP7_75t_L g3104 ( 
.A(n_2545),
.B(n_2550),
.Y(n_3104)
);

AND2x6_ASAP7_75t_L g3105 ( 
.A(n_2697),
.B(n_228),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2750),
.Y(n_3106)
);

INVx3_ASAP7_75t_L g3107 ( 
.A(n_2576),
.Y(n_3107)
);

INVx4_ASAP7_75t_L g3108 ( 
.A(n_2630),
.Y(n_3108)
);

AOI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_2684),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2545),
.B(n_231),
.Y(n_3110)
);

OR2x2_ASAP7_75t_L g3111 ( 
.A(n_2434),
.B(n_232),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2722),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_SL g3113 ( 
.A(n_2735),
.B(n_2615),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2550),
.B(n_232),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2724),
.Y(n_3115)
);

AOI22xp5_ASAP7_75t_L g3116 ( 
.A1(n_2597),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2830),
.Y(n_3117)
);

INVx1_ASAP7_75t_SL g3118 ( 
.A(n_2465),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2608),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2732),
.Y(n_3120)
);

BUFx6f_ASAP7_75t_L g3121 ( 
.A(n_2392),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_2787),
.B(n_233),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2732),
.Y(n_3123)
);

HB1xp67_ASAP7_75t_L g3124 ( 
.A(n_2449),
.Y(n_3124)
);

BUFx6f_ASAP7_75t_L g3125 ( 
.A(n_2392),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2830),
.B(n_234),
.Y(n_3126)
);

AOI221xp5_ASAP7_75t_L g3127 ( 
.A1(n_2463),
.A2(n_237),
.B1(n_239),
.B2(n_236),
.C(n_238),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2838),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2838),
.Y(n_3129)
);

INVx3_ASAP7_75t_L g3130 ( 
.A(n_2698),
.Y(n_3130)
);

NOR2xp33_ASAP7_75t_R g3131 ( 
.A(n_2560),
.B(n_235),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2468),
.Y(n_3132)
);

BUFx6f_ASAP7_75t_L g3133 ( 
.A(n_2455),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_SL g3134 ( 
.A(n_2735),
.B(n_236),
.Y(n_3134)
);

INVx3_ASAP7_75t_L g3135 ( 
.A(n_2698),
.Y(n_3135)
);

BUFx3_ASAP7_75t_L g3136 ( 
.A(n_2366),
.Y(n_3136)
);

BUFx6f_ASAP7_75t_L g3137 ( 
.A(n_2455),
.Y(n_3137)
);

INVx3_ASAP7_75t_L g3138 ( 
.A(n_2698),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2408),
.B(n_238),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2471),
.Y(n_3140)
);

OR2x2_ASAP7_75t_SL g3141 ( 
.A(n_2544),
.B(n_240),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2482),
.Y(n_3142)
);

NOR2xp33_ASAP7_75t_L g3143 ( 
.A(n_2371),
.B(n_241),
.Y(n_3143)
);

HB1xp67_ASAP7_75t_L g3144 ( 
.A(n_2767),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_SL g3145 ( 
.A(n_2735),
.B(n_241),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2841),
.B(n_242),
.Y(n_3146)
);

OAI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_2594),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_3147)
);

AND2x4_ASAP7_75t_L g3148 ( 
.A(n_2662),
.B(n_243),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2485),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2487),
.Y(n_3150)
);

AOI22x1_ASAP7_75t_L g3151 ( 
.A1(n_2705),
.A2(n_719),
.B1(n_720),
.B2(n_715),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2490),
.Y(n_3152)
);

OR2x2_ASAP7_75t_L g3153 ( 
.A(n_2813),
.B(n_244),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2408),
.B(n_245),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2410),
.B(n_246),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2674),
.Y(n_3156)
);

INVx2_ASAP7_75t_SL g3157 ( 
.A(n_2836),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2686),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2564),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_SL g3160 ( 
.A(n_2719),
.B(n_247),
.Y(n_3160)
);

AND2x4_ASAP7_75t_L g3161 ( 
.A(n_2662),
.B(n_248),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2689),
.Y(n_3162)
);

BUFx2_ASAP7_75t_L g3163 ( 
.A(n_2630),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2410),
.B(n_249),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2726),
.Y(n_3165)
);

NOR2x1_ASAP7_75t_R g3166 ( 
.A(n_2636),
.B(n_249),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2731),
.Y(n_3167)
);

INVxp67_ASAP7_75t_L g3168 ( 
.A(n_2678),
.Y(n_3168)
);

BUFx2_ASAP7_75t_L g3169 ( 
.A(n_2630),
.Y(n_3169)
);

BUFx12f_ASAP7_75t_L g3170 ( 
.A(n_2803),
.Y(n_3170)
);

AND2x4_ASAP7_75t_SL g3171 ( 
.A(n_2435),
.B(n_251),
.Y(n_3171)
);

CKINVDCx5p33_ASAP7_75t_R g3172 ( 
.A(n_2524),
.Y(n_3172)
);

NOR2xp33_ASAP7_75t_L g3173 ( 
.A(n_2363),
.B(n_251),
.Y(n_3173)
);

BUFx6f_ASAP7_75t_L g3174 ( 
.A(n_2455),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2740),
.Y(n_3175)
);

OAI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_2655),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2733),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2475),
.B(n_255),
.Y(n_3178)
);

BUFx12f_ASAP7_75t_L g3179 ( 
.A(n_2437),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_SL g3180 ( 
.A(n_2672),
.B(n_255),
.Y(n_3180)
);

BUFx12f_ASAP7_75t_L g3181 ( 
.A(n_2386),
.Y(n_3181)
);

HB1xp67_ASAP7_75t_L g3182 ( 
.A(n_2715),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_SL g3183 ( 
.A(n_2374),
.B(n_256),
.Y(n_3183)
);

AND2x2_ASAP7_75t_L g3184 ( 
.A(n_2439),
.B(n_256),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2695),
.Y(n_3185)
);

AOI22xp5_ASAP7_75t_L g3186 ( 
.A1(n_2676),
.A2(n_260),
.B1(n_257),
.B2(n_258),
.Y(n_3186)
);

BUFx2_ASAP7_75t_L g3187 ( 
.A(n_2704),
.Y(n_3187)
);

BUFx2_ASAP7_75t_L g3188 ( 
.A(n_2704),
.Y(n_3188)
);

INVx1_ASAP7_75t_SL g3189 ( 
.A(n_2716),
.Y(n_3189)
);

INVxp67_ASAP7_75t_L g3190 ( 
.A(n_2676),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_2420),
.B(n_260),
.Y(n_3191)
);

BUFx3_ASAP7_75t_L g3192 ( 
.A(n_2694),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_2700),
.Y(n_3193)
);

INVx5_ASAP7_75t_L g3194 ( 
.A(n_2461),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2736),
.Y(n_3195)
);

INVx2_ASAP7_75t_SL g3196 ( 
.A(n_2703),
.Y(n_3196)
);

INVx3_ASAP7_75t_L g3197 ( 
.A(n_2692),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2353),
.B(n_2656),
.Y(n_3198)
);

BUFx2_ASAP7_75t_L g3199 ( 
.A(n_2500),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2739),
.Y(n_3200)
);

AND2x4_ASAP7_75t_L g3201 ( 
.A(n_2692),
.B(n_261),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2627),
.Y(n_3202)
);

OAI21xp33_ASAP7_75t_L g3203 ( 
.A1(n_2681),
.A2(n_261),
.B(n_262),
.Y(n_3203)
);

INVx3_ASAP7_75t_L g3204 ( 
.A(n_2500),
.Y(n_3204)
);

NAND2x1_ASAP7_75t_L g3205 ( 
.A(n_2461),
.B(n_721),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2718),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2534),
.Y(n_3207)
);

NOR2xp33_ASAP7_75t_SL g3208 ( 
.A(n_2548),
.B(n_262),
.Y(n_3208)
);

OAI22xp5_ASAP7_75t_L g3209 ( 
.A1(n_2605),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_3209)
);

INVx2_ASAP7_75t_L g3210 ( 
.A(n_2737),
.Y(n_3210)
);

CKINVDCx5p33_ASAP7_75t_R g3211 ( 
.A(n_2728),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2423),
.B(n_263),
.Y(n_3212)
);

INVx3_ASAP7_75t_L g3213 ( 
.A(n_2697),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_SL g3214 ( 
.A(n_2646),
.B(n_264),
.Y(n_3214)
);

BUFx3_ASAP7_75t_L g3215 ( 
.A(n_2583),
.Y(n_3215)
);

BUFx2_ASAP7_75t_L g3216 ( 
.A(n_2723),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_2349),
.B(n_265),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2592),
.B(n_267),
.Y(n_3218)
);

AND2x6_ASAP7_75t_L g3219 ( 
.A(n_2697),
.B(n_268),
.Y(n_3219)
);

CKINVDCx5p33_ASAP7_75t_R g3220 ( 
.A(n_2361),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2598),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2562),
.Y(n_3222)
);

BUFx2_ASAP7_75t_L g3223 ( 
.A(n_2723),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2421),
.B(n_269),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2600),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_2569),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2442),
.B(n_269),
.Y(n_3227)
);

AND2x4_ASAP7_75t_L g3228 ( 
.A(n_2688),
.B(n_270),
.Y(n_3228)
);

BUFx6f_ASAP7_75t_L g3229 ( 
.A(n_2461),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2590),
.Y(n_3230)
);

CKINVDCx5p33_ASAP7_75t_R g3231 ( 
.A(n_2784),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_2454),
.B(n_270),
.Y(n_3232)
);

CKINVDCx5p33_ASAP7_75t_R g3233 ( 
.A(n_2837),
.Y(n_3233)
);

AOI22xp33_ASAP7_75t_L g3234 ( 
.A1(n_2666),
.A2(n_274),
.B1(n_271),
.B2(n_273),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_2458),
.B(n_275),
.Y(n_3235)
);

INVx3_ASAP7_75t_L g3236 ( 
.A(n_2632),
.Y(n_3236)
);

AND2x4_ASAP7_75t_L g3237 ( 
.A(n_2616),
.B(n_275),
.Y(n_3237)
);

BUFx6f_ASAP7_75t_L g3238 ( 
.A(n_2467),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_SL g3239 ( 
.A(n_2467),
.B(n_276),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2586),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_SL g3241 ( 
.A(n_2467),
.B(n_276),
.Y(n_3241)
);

CKINVDCx20_ASAP7_75t_R g3242 ( 
.A(n_2351),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_SL g3243 ( 
.A(n_2483),
.B(n_277),
.Y(n_3243)
);

INVx2_ASAP7_75t_SL g3244 ( 
.A(n_2702),
.Y(n_3244)
);

BUFx3_ASAP7_75t_L g3245 ( 
.A(n_2632),
.Y(n_3245)
);

AND2x4_ASAP7_75t_L g3246 ( 
.A(n_2693),
.B(n_277),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2586),
.Y(n_3247)
);

INVx1_ASAP7_75t_SL g3248 ( 
.A(n_2650),
.Y(n_3248)
);

AND2x4_ASAP7_75t_L g3249 ( 
.A(n_2707),
.B(n_2561),
.Y(n_3249)
);

BUFx2_ASAP7_75t_SL g3250 ( 
.A(n_2636),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2472),
.B(n_278),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2610),
.Y(n_3252)
);

NOR2x1_ASAP7_75t_L g3253 ( 
.A(n_2658),
.B(n_278),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2476),
.B(n_279),
.Y(n_3254)
);

AND2x4_ASAP7_75t_L g3255 ( 
.A(n_2634),
.B(n_280),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_2378),
.B(n_280),
.Y(n_3256)
);

CKINVDCx20_ASAP7_75t_R g3257 ( 
.A(n_2680),
.Y(n_3257)
);

BUFx3_ASAP7_75t_L g3258 ( 
.A(n_2634),
.Y(n_3258)
);

INVx3_ASAP7_75t_L g3259 ( 
.A(n_2483),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_2614),
.Y(n_3260)
);

INVx1_ASAP7_75t_SL g3261 ( 
.A(n_2378),
.Y(n_3261)
);

NOR2xp67_ASAP7_75t_L g3262 ( 
.A(n_2658),
.B(n_281),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_2478),
.B(n_281),
.Y(n_3263)
);

AND2x2_ASAP7_75t_L g3264 ( 
.A(n_2438),
.B(n_282),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2589),
.Y(n_3265)
);

BUFx6f_ASAP7_75t_L g3266 ( 
.A(n_2483),
.Y(n_3266)
);

BUFx3_ASAP7_75t_L g3267 ( 
.A(n_2624),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2575),
.Y(n_3268)
);

INVxp67_ASAP7_75t_L g3269 ( 
.A(n_2415),
.Y(n_3269)
);

AND2x4_ASAP7_75t_L g3270 ( 
.A(n_2521),
.B(n_283),
.Y(n_3270)
);

INVx3_ASAP7_75t_L g3271 ( 
.A(n_2859),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_3207),
.B(n_2474),
.Y(n_3272)
);

CKINVDCx5p33_ASAP7_75t_R g3273 ( 
.A(n_2969),
.Y(n_3273)
);

INVx4_ASAP7_75t_L g3274 ( 
.A(n_2875),
.Y(n_3274)
);

AND2x4_ASAP7_75t_L g3275 ( 
.A(n_2923),
.B(n_2502),
.Y(n_3275)
);

O2A1O1Ixp33_ASAP7_75t_L g3276 ( 
.A1(n_3007),
.A2(n_2777),
.B(n_2823),
.C(n_2795),
.Y(n_3276)
);

INVx2_ASAP7_75t_SL g3277 ( 
.A(n_2922),
.Y(n_3277)
);

INVx3_ASAP7_75t_L g3278 ( 
.A(n_2859),
.Y(n_3278)
);

INVx3_ASAP7_75t_L g3279 ( 
.A(n_2847),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2846),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2850),
.Y(n_3281)
);

BUFx12f_ASAP7_75t_L g3282 ( 
.A(n_2922),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_3069),
.Y(n_3283)
);

BUFx2_ASAP7_75t_L g3284 ( 
.A(n_3108),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_3082),
.Y(n_3285)
);

OAI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_3189),
.A2(n_2648),
.B1(n_2825),
.B2(n_2481),
.Y(n_3286)
);

AND2x2_ASAP7_75t_L g3287 ( 
.A(n_2958),
.B(n_2666),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2854),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2872),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2958),
.B(n_2908),
.Y(n_3290)
);

AOI21xp5_ASAP7_75t_L g3291 ( 
.A1(n_3058),
.A2(n_3102),
.B(n_3208),
.Y(n_3291)
);

INVxp67_ASAP7_75t_L g3292 ( 
.A(n_2848),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_2852),
.B(n_2667),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_3051),
.A2(n_2589),
.B(n_2554),
.Y(n_3294)
);

INVx3_ASAP7_75t_L g3295 ( 
.A(n_2855),
.Y(n_3295)
);

BUFx3_ASAP7_75t_L g3296 ( 
.A(n_3022),
.Y(n_3296)
);

AOI22xp5_ASAP7_75t_L g3297 ( 
.A1(n_3039),
.A2(n_2809),
.B1(n_2480),
.B2(n_2667),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_2904),
.B(n_2426),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_2981),
.B(n_2367),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2874),
.Y(n_3300)
);

NAND3xp33_ASAP7_75t_L g3301 ( 
.A(n_2927),
.B(n_2775),
.C(n_2629),
.Y(n_3301)
);

CKINVDCx20_ASAP7_75t_R g3302 ( 
.A(n_2933),
.Y(n_3302)
);

OAI22xp33_ASAP7_75t_L g3303 ( 
.A1(n_2885),
.A2(n_2754),
.B1(n_2812),
.B2(n_2653),
.Y(n_3303)
);

NOR2x1_ASAP7_75t_L g3304 ( 
.A(n_2885),
.B(n_2502),
.Y(n_3304)
);

HB1xp67_ASAP7_75t_L g3305 ( 
.A(n_2944),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_2876),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3095),
.Y(n_3307)
);

AND2x4_ASAP7_75t_L g3308 ( 
.A(n_2923),
.B(n_2624),
.Y(n_3308)
);

BUFx3_ASAP7_75t_L g3309 ( 
.A(n_3181),
.Y(n_3309)
);

BUFx3_ASAP7_75t_L g3310 ( 
.A(n_2926),
.Y(n_3310)
);

AOI22xp33_ASAP7_75t_L g3311 ( 
.A1(n_3039),
.A2(n_2647),
.B1(n_2631),
.B2(n_2721),
.Y(n_3311)
);

HB1xp67_ASAP7_75t_L g3312 ( 
.A(n_3081),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2877),
.Y(n_3313)
);

NAND2x1_ASAP7_75t_L g3314 ( 
.A(n_3108),
.B(n_2723),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2858),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3268),
.B(n_2409),
.Y(n_3316)
);

AND2x2_ASAP7_75t_L g3317 ( 
.A(n_3028),
.B(n_2401),
.Y(n_3317)
);

CKINVDCx11_ASAP7_75t_R g3318 ( 
.A(n_2995),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_3099),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3101),
.Y(n_3320)
);

AND2x4_ASAP7_75t_L g3321 ( 
.A(n_2925),
.B(n_2407),
.Y(n_3321)
);

A2O1A1Ixp33_ASAP7_75t_L g3322 ( 
.A1(n_3045),
.A2(n_2612),
.B(n_2824),
.C(n_2595),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2843),
.B(n_2601),
.Y(n_3323)
);

AOI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_3039),
.A2(n_2828),
.B1(n_2553),
.B2(n_2639),
.Y(n_3324)
);

A2O1A1Ixp33_ASAP7_75t_L g3325 ( 
.A1(n_3045),
.A2(n_3262),
.B(n_2997),
.C(n_2937),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_3029),
.B(n_2403),
.Y(n_3326)
);

BUFx2_ASAP7_75t_L g3327 ( 
.A(n_3041),
.Y(n_3327)
);

BUFx4f_ASAP7_75t_SL g3328 ( 
.A(n_2851),
.Y(n_3328)
);

INVx5_ASAP7_75t_L g3329 ( 
.A(n_3105),
.Y(n_3329)
);

BUFx3_ASAP7_75t_L g3330 ( 
.A(n_2926),
.Y(n_3330)
);

BUFx6f_ASAP7_75t_L g3331 ( 
.A(n_2982),
.Y(n_3331)
);

OAI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_2954),
.A2(n_2738),
.B1(n_2660),
.B2(n_2649),
.Y(n_3332)
);

CKINVDCx16_ASAP7_75t_R g3333 ( 
.A(n_2865),
.Y(n_3333)
);

INVx2_ASAP7_75t_SL g3334 ( 
.A(n_3018),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3106),
.Y(n_3335)
);

BUFx6f_ASAP7_75t_L g3336 ( 
.A(n_2983),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_2864),
.Y(n_3337)
);

BUFx12f_ASAP7_75t_L g3338 ( 
.A(n_2966),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_3117),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_2849),
.B(n_2603),
.Y(n_3340)
);

AOI22xp33_ASAP7_75t_L g3341 ( 
.A1(n_3039),
.A2(n_2528),
.B1(n_2633),
.B2(n_2626),
.Y(n_3341)
);

OAI21x1_ASAP7_75t_L g3342 ( 
.A1(n_3240),
.A2(n_2565),
.B(n_2714),
.Y(n_3342)
);

BUFx6f_ASAP7_75t_L g3343 ( 
.A(n_3194),
.Y(n_3343)
);

INVx2_ASAP7_75t_SL g3344 ( 
.A(n_3014),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3035),
.B(n_2369),
.Y(n_3345)
);

NAND2x1p5_ASAP7_75t_L g3346 ( 
.A(n_2866),
.B(n_2488),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_2880),
.Y(n_3347)
);

BUFx6f_ASAP7_75t_L g3348 ( 
.A(n_3194),
.Y(n_3348)
);

BUFx8_ASAP7_75t_L g3349 ( 
.A(n_3187),
.Y(n_3349)
);

BUFx2_ASAP7_75t_SL g3350 ( 
.A(n_3041),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2862),
.B(n_2448),
.Y(n_3351)
);

OAI221xp5_ASAP7_75t_L g3352 ( 
.A1(n_3190),
.A2(n_2406),
.B1(n_2759),
.B2(n_2785),
.C(n_2743),
.Y(n_3352)
);

INVx2_ASAP7_75t_SL g3353 ( 
.A(n_3014),
.Y(n_3353)
);

OAI22xp5_ASAP7_75t_L g3354 ( 
.A1(n_2931),
.A2(n_2643),
.B1(n_2622),
.B2(n_2815),
.Y(n_3354)
);

O2A1O1Ixp5_ASAP7_75t_L g3355 ( 
.A1(n_2893),
.A2(n_2734),
.B(n_2679),
.C(n_2617),
.Y(n_3355)
);

BUFx2_ASAP7_75t_L g3356 ( 
.A(n_3041),
.Y(n_3356)
);

AOI22xp33_ASAP7_75t_L g3357 ( 
.A1(n_2925),
.A2(n_3119),
.B1(n_2931),
.B2(n_2937),
.Y(n_3357)
);

BUFx6f_ASAP7_75t_L g3358 ( 
.A(n_3194),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3129),
.Y(n_3359)
);

OR2x6_ASAP7_75t_L g3360 ( 
.A(n_3250),
.B(n_2665),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2900),
.B(n_2383),
.Y(n_3361)
);

NOR2xp67_ASAP7_75t_L g3362 ( 
.A(n_3168),
.B(n_2696),
.Y(n_3362)
);

OR2x6_ASAP7_75t_L g3363 ( 
.A(n_3188),
.B(n_2350),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2924),
.Y(n_3364)
);

OR2x6_ASAP7_75t_L g3365 ( 
.A(n_2903),
.B(n_2673),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_2928),
.Y(n_3366)
);

OAI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_3141),
.A2(n_2820),
.B1(n_2835),
.B2(n_2687),
.Y(n_3367)
);

NOR2xp67_ASAP7_75t_SL g3368 ( 
.A(n_3163),
.B(n_2488),
.Y(n_3368)
);

BUFx2_ASAP7_75t_SL g3369 ( 
.A(n_3041),
.Y(n_3369)
);

AO22x1_ASAP7_75t_L g3370 ( 
.A1(n_2842),
.A2(n_3100),
.B1(n_3219),
.B2(n_3105),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_3269),
.B(n_2380),
.Y(n_3371)
);

BUFx3_ASAP7_75t_L g3372 ( 
.A(n_2940),
.Y(n_3372)
);

BUFx2_ASAP7_75t_L g3373 ( 
.A(n_3041),
.Y(n_3373)
);

AOI21xp5_ASAP7_75t_L g3374 ( 
.A1(n_3150),
.A2(n_2520),
.B(n_2523),
.Y(n_3374)
);

OAI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_3248),
.A2(n_2581),
.B1(n_2588),
.B2(n_2587),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_2932),
.Y(n_3376)
);

INVx3_ASAP7_75t_L g3377 ( 
.A(n_3179),
.Y(n_3377)
);

BUFx3_ASAP7_75t_L g3378 ( 
.A(n_2940),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_2913),
.Y(n_3379)
);

INVx5_ASAP7_75t_L g3380 ( 
.A(n_3105),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2952),
.Y(n_3381)
);

OAI22xp5_ASAP7_75t_L g3382 ( 
.A1(n_3169),
.A2(n_2566),
.B1(n_2670),
.B2(n_2664),
.Y(n_3382)
);

CKINVDCx5p33_ASAP7_75t_R g3383 ( 
.A(n_2994),
.Y(n_3383)
);

AND2x4_ASAP7_75t_L g3384 ( 
.A(n_2871),
.B(n_2712),
.Y(n_3384)
);

CKINVDCx5p33_ASAP7_75t_R g3385 ( 
.A(n_2896),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_2947),
.B(n_2384),
.Y(n_3386)
);

NOR2xp67_ASAP7_75t_L g3387 ( 
.A(n_3008),
.B(n_2682),
.Y(n_3387)
);

CKINVDCx5p33_ASAP7_75t_R g3388 ( 
.A(n_2905),
.Y(n_3388)
);

INVx2_ASAP7_75t_SL g3389 ( 
.A(n_2906),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_2957),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_2929),
.Y(n_3391)
);

INVx4_ASAP7_75t_L g3392 ( 
.A(n_2964),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_2938),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3261),
.B(n_2385),
.Y(n_3394)
);

AO21x2_ASAP7_75t_L g3395 ( 
.A1(n_3214),
.A2(n_2706),
.B(n_2533),
.Y(n_3395)
);

BUFx2_ASAP7_75t_L g3396 ( 
.A(n_2871),
.Y(n_3396)
);

BUFx2_ASAP7_75t_L g3397 ( 
.A(n_3216),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_2959),
.Y(n_3398)
);

O2A1O1Ixp33_ASAP7_75t_L g3399 ( 
.A1(n_3180),
.A2(n_2701),
.B(n_2396),
.C(n_2685),
.Y(n_3399)
);

HB1xp67_ASAP7_75t_L g3400 ( 
.A(n_3182),
.Y(n_3400)
);

BUFx6f_ASAP7_75t_L g3401 ( 
.A(n_3016),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_2961),
.B(n_2390),
.Y(n_3402)
);

AND2x4_ASAP7_75t_L g3403 ( 
.A(n_2935),
.B(n_2712),
.Y(n_3403)
);

INVx4_ASAP7_75t_L g3404 ( 
.A(n_2911),
.Y(n_3404)
);

CKINVDCx6p67_ASAP7_75t_R g3405 ( 
.A(n_3096),
.Y(n_3405)
);

BUFx3_ASAP7_75t_L g3406 ( 
.A(n_3192),
.Y(n_3406)
);

O2A1O1Ixp33_ASAP7_75t_SL g3407 ( 
.A1(n_2873),
.A2(n_2602),
.B(n_2515),
.C(n_2621),
.Y(n_3407)
);

AOI22xp33_ASAP7_75t_L g3408 ( 
.A1(n_3173),
.A2(n_2723),
.B1(n_2730),
.B2(n_2675),
.Y(n_3408)
);

INVx2_ASAP7_75t_SL g3409 ( 
.A(n_2930),
.Y(n_3409)
);

BUFx6f_ASAP7_75t_L g3410 ( 
.A(n_2844),
.Y(n_3410)
);

BUFx8_ASAP7_75t_L g3411 ( 
.A(n_3170),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_2939),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_2962),
.B(n_2391),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_3152),
.A2(n_3057),
.B(n_3054),
.Y(n_3414)
);

INVx3_ASAP7_75t_L g3415 ( 
.A(n_2960),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2970),
.Y(n_3416)
);

O2A1O1Ixp33_ASAP7_75t_SL g3417 ( 
.A1(n_3160),
.A2(n_2574),
.B(n_2607),
.C(n_2542),
.Y(n_3417)
);

AOI21xp33_ASAP7_75t_L g3418 ( 
.A1(n_3030),
.A2(n_2505),
.B(n_3043),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_2977),
.Y(n_3419)
);

AOI22xp5_ASAP7_75t_L g3420 ( 
.A1(n_3242),
.A2(n_2683),
.B1(n_2742),
.B2(n_2713),
.Y(n_3420)
);

AOI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_2845),
.A2(n_2710),
.B1(n_2546),
.B2(n_2691),
.Y(n_3421)
);

INVx1_ASAP7_75t_SL g3422 ( 
.A(n_2971),
.Y(n_3422)
);

BUFx3_ASAP7_75t_L g3423 ( 
.A(n_3038),
.Y(n_3423)
);

AOI22xp33_ASAP7_75t_L g3424 ( 
.A1(n_2978),
.A2(n_2499),
.B1(n_2538),
.B2(n_2445),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_2984),
.Y(n_3425)
);

A2O1A1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_3253),
.A2(n_2558),
.B(n_2640),
.C(n_2753),
.Y(n_3426)
);

AOI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_3063),
.A2(n_2525),
.B(n_2488),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_2988),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3004),
.B(n_2671),
.Y(n_3429)
);

BUFx2_ASAP7_75t_L g3430 ( 
.A(n_3223),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3020),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3013),
.B(n_2671),
.Y(n_3432)
);

AOI21x1_ASAP7_75t_L g3433 ( 
.A1(n_3247),
.A2(n_2741),
.B(n_2780),
.Y(n_3433)
);

AND2x4_ASAP7_75t_SL g3434 ( 
.A(n_2960),
.B(n_2375),
.Y(n_3434)
);

HB1xp67_ASAP7_75t_L g3435 ( 
.A(n_2890),
.Y(n_3435)
);

INVx5_ASAP7_75t_L g3436 ( 
.A(n_3105),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3017),
.Y(n_3437)
);

BUFx3_ASAP7_75t_L g3438 ( 
.A(n_3136),
.Y(n_3438)
);

BUFx2_ASAP7_75t_L g3439 ( 
.A(n_3265),
.Y(n_3439)
);

INVx4_ASAP7_75t_L g3440 ( 
.A(n_2963),
.Y(n_3440)
);

CKINVDCx6p67_ASAP7_75t_R g3441 ( 
.A(n_3257),
.Y(n_3441)
);

BUFx2_ASAP7_75t_L g3442 ( 
.A(n_2844),
.Y(n_3442)
);

AOI22xp5_ASAP7_75t_L g3443 ( 
.A1(n_2853),
.A2(n_2521),
.B1(n_2727),
.B2(n_2729),
.Y(n_3443)
);

BUFx6f_ASAP7_75t_L g3444 ( 
.A(n_2844),
.Y(n_3444)
);

AND2x6_ASAP7_75t_L g3445 ( 
.A(n_3270),
.B(n_2525),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3024),
.Y(n_3446)
);

AND2x2_ASAP7_75t_L g3447 ( 
.A(n_3078),
.B(n_283),
.Y(n_3447)
);

BUFx6f_ASAP7_75t_L g3448 ( 
.A(n_2920),
.Y(n_3448)
);

NOR2xp33_ASAP7_75t_L g3449 ( 
.A(n_3166),
.B(n_2375),
.Y(n_3449)
);

INVx3_ASAP7_75t_L g3450 ( 
.A(n_3215),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3156),
.Y(n_3451)
);

BUFx3_ASAP7_75t_L g3452 ( 
.A(n_3196),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3098),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_2868),
.A2(n_2486),
.B1(n_2510),
.B2(n_2429),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_L g3455 ( 
.A1(n_2992),
.A2(n_2486),
.B1(n_2510),
.B2(n_2429),
.Y(n_3455)
);

BUFx2_ASAP7_75t_L g3456 ( 
.A(n_2920),
.Y(n_3456)
);

AND2x2_ASAP7_75t_SL g3457 ( 
.A(n_3171),
.B(n_2525),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3103),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3167),
.Y(n_3459)
);

INVx3_ASAP7_75t_L g3460 ( 
.A(n_3267),
.Y(n_3460)
);

AND2x2_ASAP7_75t_L g3461 ( 
.A(n_3256),
.B(n_284),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_L g3462 ( 
.A1(n_3023),
.A2(n_2752),
.B1(n_2788),
.B2(n_2786),
.Y(n_3462)
);

CKINVDCx5p33_ASAP7_75t_R g3463 ( 
.A(n_2968),
.Y(n_3463)
);

INVx3_ASAP7_75t_L g3464 ( 
.A(n_3245),
.Y(n_3464)
);

INVx4_ASAP7_75t_L g3465 ( 
.A(n_3055),
.Y(n_3465)
);

AND2x4_ASAP7_75t_L g3466 ( 
.A(n_3012),
.B(n_2752),
.Y(n_3466)
);

INVx3_ASAP7_75t_L g3467 ( 
.A(n_3258),
.Y(n_3467)
);

BUFx6f_ASAP7_75t_L g3468 ( 
.A(n_2920),
.Y(n_3468)
);

AOI222xp33_ASAP7_75t_L g3469 ( 
.A1(n_2916),
.A2(n_2788),
.B1(n_2786),
.B2(n_288),
.C1(n_290),
.C2(n_285),
.Y(n_3469)
);

HB1xp67_ASAP7_75t_L g3470 ( 
.A(n_2950),
.Y(n_3470)
);

BUFx6f_ASAP7_75t_L g3471 ( 
.A(n_2965),
.Y(n_3471)
);

AOI22xp33_ASAP7_75t_L g3472 ( 
.A1(n_2975),
.A2(n_2717),
.B1(n_2551),
.B2(n_2557),
.Y(n_3472)
);

BUFx4f_ASAP7_75t_L g3473 ( 
.A(n_3219),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3085),
.B(n_285),
.Y(n_3474)
);

BUFx3_ASAP7_75t_L g3475 ( 
.A(n_2909),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3112),
.B(n_287),
.Y(n_3476)
);

BUFx12f_ASAP7_75t_L g3477 ( 
.A(n_3172),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3115),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3025),
.Y(n_3479)
);

AOI21xp5_ASAP7_75t_L g3480 ( 
.A1(n_3064),
.A2(n_2551),
.B(n_2526),
.Y(n_3480)
);

BUFx10_ASAP7_75t_L g3481 ( 
.A(n_2986),
.Y(n_3481)
);

AND2x4_ASAP7_75t_L g3482 ( 
.A(n_2919),
.B(n_2526),
.Y(n_3482)
);

INVx3_ASAP7_75t_L g3483 ( 
.A(n_2903),
.Y(n_3483)
);

NOR2xp33_ASAP7_75t_L g3484 ( 
.A(n_3233),
.B(n_289),
.Y(n_3484)
);

AND2x4_ASAP7_75t_L g3485 ( 
.A(n_2912),
.B(n_2526),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3079),
.A2(n_2557),
.B(n_2551),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3026),
.Y(n_3487)
);

AO32x1_ASAP7_75t_L g3488 ( 
.A1(n_3074),
.A2(n_2585),
.A3(n_2609),
.B1(n_2570),
.B2(n_2557),
.Y(n_3488)
);

AND2x4_ASAP7_75t_L g3489 ( 
.A(n_2912),
.B(n_2570),
.Y(n_3489)
);

INVx3_ASAP7_75t_L g3490 ( 
.A(n_2860),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3128),
.B(n_290),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_L g3492 ( 
.A(n_3118),
.B(n_291),
.Y(n_3492)
);

NOR2xp67_ASAP7_75t_L g3493 ( 
.A(n_3220),
.B(n_291),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3225),
.B(n_292),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3033),
.Y(n_3495)
);

AOI22xp33_ASAP7_75t_L g3496 ( 
.A1(n_3184),
.A2(n_2585),
.B1(n_2609),
.B2(n_2570),
.Y(n_3496)
);

BUFx2_ASAP7_75t_L g3497 ( 
.A(n_2965),
.Y(n_3497)
);

NAND2x2_ASAP7_75t_L g3498 ( 
.A(n_2914),
.B(n_294),
.Y(n_3498)
);

AND2x6_ASAP7_75t_L g3499 ( 
.A(n_3270),
.B(n_2585),
.Y(n_3499)
);

BUFx2_ASAP7_75t_L g3500 ( 
.A(n_2965),
.Y(n_3500)
);

NOR2xp67_ASAP7_75t_SL g3501 ( 
.A(n_2945),
.B(n_2609),
.Y(n_3501)
);

AOI21xp5_ASAP7_75t_L g3502 ( 
.A1(n_3084),
.A2(n_2757),
.B(n_2748),
.Y(n_3502)
);

INVx3_ASAP7_75t_L g3503 ( 
.A(n_2860),
.Y(n_3503)
);

AND2x2_ASAP7_75t_L g3504 ( 
.A(n_2881),
.B(n_294),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_SL g3505 ( 
.A(n_3148),
.B(n_2782),
.Y(n_3505)
);

INVx2_ASAP7_75t_SL g3506 ( 
.A(n_2996),
.Y(n_3506)
);

BUFx3_ASAP7_75t_L g3507 ( 
.A(n_3199),
.Y(n_3507)
);

INVx2_ASAP7_75t_L g3508 ( 
.A(n_3034),
.Y(n_3508)
);

CKINVDCx5p33_ASAP7_75t_R g3509 ( 
.A(n_3131),
.Y(n_3509)
);

OA22x2_ASAP7_75t_L g3510 ( 
.A1(n_3211),
.A2(n_3113),
.B1(n_3186),
.B2(n_3231),
.Y(n_3510)
);

INVx2_ASAP7_75t_SL g3511 ( 
.A(n_2986),
.Y(n_3511)
);

AOI221xp5_ASAP7_75t_L g3512 ( 
.A1(n_3198),
.A2(n_2782),
.B1(n_2757),
.B2(n_2748),
.C(n_297),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3165),
.Y(n_3513)
);

AOI22xp33_ASAP7_75t_L g3514 ( 
.A1(n_3264),
.A2(n_2757),
.B1(n_2782),
.B2(n_2748),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3175),
.Y(n_3515)
);

AOI22xp5_ASAP7_75t_L g3516 ( 
.A1(n_2976),
.A2(n_298),
.B1(n_295),
.B2(n_296),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3040),
.Y(n_3517)
);

INVx3_ASAP7_75t_L g3518 ( 
.A(n_2894),
.Y(n_3518)
);

BUFx6f_ASAP7_75t_L g3519 ( 
.A(n_3266),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3158),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3049),
.Y(n_3521)
);

HB1xp67_ASAP7_75t_L g3522 ( 
.A(n_2955),
.Y(n_3522)
);

CKINVDCx5p33_ASAP7_75t_R g3523 ( 
.A(n_2883),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3050),
.Y(n_3524)
);

INVx3_ASAP7_75t_L g3525 ( 
.A(n_2894),
.Y(n_3525)
);

OR2x6_ASAP7_75t_L g3526 ( 
.A(n_3148),
.B(n_296),
.Y(n_3526)
);

INVxp67_ASAP7_75t_L g3527 ( 
.A(n_2934),
.Y(n_3527)
);

OAI22xp5_ASAP7_75t_L g3528 ( 
.A1(n_2868),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_3528)
);

NAND3xp33_ASAP7_75t_L g3529 ( 
.A(n_2899),
.B(n_301),
.C(n_303),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3244),
.B(n_301),
.Y(n_3530)
);

O2A1O1Ixp33_ASAP7_75t_SL g3531 ( 
.A1(n_3067),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_3531)
);

HB1xp67_ASAP7_75t_L g3532 ( 
.A(n_3015),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_2941),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3222),
.Y(n_3534)
);

AOI22xp5_ASAP7_75t_L g3535 ( 
.A1(n_2882),
.A2(n_308),
.B1(n_305),
.B2(n_306),
.Y(n_3535)
);

BUFx6f_ASAP7_75t_L g3536 ( 
.A(n_3266),
.Y(n_3536)
);

OAI22xp5_ASAP7_75t_L g3537 ( 
.A1(n_3234),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_3221),
.B(n_309),
.Y(n_3538)
);

BUFx6f_ASAP7_75t_L g3539 ( 
.A(n_3266),
.Y(n_3539)
);

BUFx2_ASAP7_75t_L g3540 ( 
.A(n_2972),
.Y(n_3540)
);

INVx1_ASAP7_75t_SL g3541 ( 
.A(n_3061),
.Y(n_3541)
);

OAI22x1_ASAP7_75t_L g3542 ( 
.A1(n_3255),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_2980),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_2889),
.B(n_311),
.Y(n_3544)
);

OR2x6_ASAP7_75t_L g3545 ( 
.A(n_3161),
.B(n_314),
.Y(n_3545)
);

OR2x2_ASAP7_75t_L g3546 ( 
.A(n_3027),
.B(n_314),
.Y(n_3546)
);

OR2x2_ASAP7_75t_L g3547 ( 
.A(n_3083),
.B(n_3226),
.Y(n_3547)
);

INVxp67_ASAP7_75t_SL g3548 ( 
.A(n_3237),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3230),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3202),
.B(n_315),
.Y(n_3550)
);

OAI21xp33_ASAP7_75t_L g3551 ( 
.A1(n_3212),
.A2(n_317),
.B(n_318),
.Y(n_3551)
);

INVx4_ASAP7_75t_L g3552 ( 
.A(n_3055),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3037),
.Y(n_3553)
);

INVx4_ASAP7_75t_L g3554 ( 
.A(n_3219),
.Y(n_3554)
);

INVxp67_ASAP7_75t_SL g3555 ( 
.A(n_3237),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_2989),
.Y(n_3556)
);

BUFx6f_ASAP7_75t_L g3557 ( 
.A(n_2972),
.Y(n_3557)
);

OAI22xp33_ASAP7_75t_L g3558 ( 
.A1(n_3091),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3132),
.Y(n_3559)
);

INVx2_ASAP7_75t_SL g3560 ( 
.A(n_3255),
.Y(n_3560)
);

INVx5_ASAP7_75t_L g3561 ( 
.A(n_3219),
.Y(n_3561)
);

BUFx3_ASAP7_75t_L g3562 ( 
.A(n_3036),
.Y(n_3562)
);

INVx1_ASAP7_75t_SL g3563 ( 
.A(n_3124),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3140),
.Y(n_3564)
);

OR2x6_ASAP7_75t_L g3565 ( 
.A(n_3161),
.B(n_3201),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_2897),
.B(n_320),
.Y(n_3566)
);

BUFx8_ASAP7_75t_SL g3567 ( 
.A(n_3191),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3252),
.B(n_3260),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3142),
.Y(n_3569)
);

AND2x4_ASAP7_75t_L g3570 ( 
.A(n_3157),
.B(n_320),
.Y(n_3570)
);

BUFx2_ASAP7_75t_L g3571 ( 
.A(n_2972),
.Y(n_3571)
);

INVx4_ASAP7_75t_L g3572 ( 
.A(n_2915),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3149),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_2990),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_2993),
.Y(n_3575)
);

NOR2xp33_ASAP7_75t_SL g3576 ( 
.A(n_2956),
.B(n_321),
.Y(n_3576)
);

BUFx6f_ASAP7_75t_L g3577 ( 
.A(n_2979),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3087),
.B(n_322),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_2999),
.Y(n_3579)
);

INVx5_ASAP7_75t_L g3580 ( 
.A(n_2979),
.Y(n_3580)
);

BUFx6f_ASAP7_75t_L g3581 ( 
.A(n_2979),
.Y(n_3581)
);

BUFx2_ASAP7_75t_L g3582 ( 
.A(n_3000),
.Y(n_3582)
);

AND2x4_ASAP7_75t_L g3583 ( 
.A(n_3249),
.B(n_322),
.Y(n_3583)
);

BUFx3_ASAP7_75t_L g3584 ( 
.A(n_3144),
.Y(n_3584)
);

BUFx3_ASAP7_75t_L g3585 ( 
.A(n_3130),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_3001),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3006),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3010),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3011),
.Y(n_3589)
);

BUFx6f_ASAP7_75t_L g3590 ( 
.A(n_3000),
.Y(n_3590)
);

OAI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_3224),
.A2(n_2886),
.B(n_3009),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_2991),
.Y(n_3592)
);

BUFx6f_ASAP7_75t_L g3593 ( 
.A(n_3000),
.Y(n_3593)
);

BUFx2_ASAP7_75t_L g3594 ( 
.A(n_3005),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3046),
.Y(n_3595)
);

INVx3_ASAP7_75t_L g3596 ( 
.A(n_2915),
.Y(n_3596)
);

AND2x4_ASAP7_75t_L g3597 ( 
.A(n_2974),
.B(n_324),
.Y(n_3597)
);

BUFx3_ASAP7_75t_L g3598 ( 
.A(n_3130),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3088),
.A2(n_727),
.B(n_723),
.Y(n_3599)
);

CKINVDCx5p33_ASAP7_75t_R g3600 ( 
.A(n_3066),
.Y(n_3600)
);

NAND3xp33_ASAP7_75t_SL g3601 ( 
.A(n_3031),
.B(n_324),
.C(n_325),
.Y(n_3601)
);

NOR2xp33_ASAP7_75t_L g3602 ( 
.A(n_3052),
.B(n_326),
.Y(n_3602)
);

AOI222xp33_ASAP7_75t_L g3603 ( 
.A1(n_3089),
.A2(n_330),
.B1(n_333),
.B2(n_326),
.C1(n_328),
.C2(n_331),
.Y(n_3603)
);

INVx2_ASAP7_75t_SL g3604 ( 
.A(n_3204),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3092),
.B(n_331),
.Y(n_3605)
);

INVx3_ASAP7_75t_L g3606 ( 
.A(n_2918),
.Y(n_3606)
);

AOI21xp5_ASAP7_75t_SL g3607 ( 
.A1(n_3201),
.A2(n_334),
.B(n_335),
.Y(n_3607)
);

INVx1_ASAP7_75t_SL g3608 ( 
.A(n_3153),
.Y(n_3608)
);

AOI22xp33_ASAP7_75t_L g3609 ( 
.A1(n_3249),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3047),
.Y(n_3610)
);

HB1xp67_ASAP7_75t_L g3611 ( 
.A(n_3093),
.Y(n_3611)
);

INVx3_ASAP7_75t_L g3612 ( 
.A(n_2918),
.Y(n_3612)
);

NOR2xp33_ASAP7_75t_L g3613 ( 
.A(n_3111),
.B(n_336),
.Y(n_3613)
);

HB1xp67_ASAP7_75t_L g3614 ( 
.A(n_3104),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3094),
.B(n_337),
.Y(n_3615)
);

BUFx4f_ASAP7_75t_SL g3616 ( 
.A(n_2949),
.Y(n_3616)
);

INVx6_ASAP7_75t_L g3617 ( 
.A(n_2974),
.Y(n_3617)
);

OAI21x1_ASAP7_75t_L g3618 ( 
.A1(n_3314),
.A2(n_3205),
.B(n_2902),
.Y(n_3618)
);

BUFx6f_ASAP7_75t_L g3619 ( 
.A(n_3343),
.Y(n_3619)
);

BUFx6f_ASAP7_75t_L g3620 ( 
.A(n_3343),
.Y(n_3620)
);

OAI221xp5_ASAP7_75t_L g3621 ( 
.A1(n_3297),
.A2(n_3048),
.B1(n_3060),
.B2(n_3143),
.C(n_3072),
.Y(n_3621)
);

INVx2_ASAP7_75t_SL g3622 ( 
.A(n_3282),
.Y(n_3622)
);

OAI21x1_ASAP7_75t_L g3623 ( 
.A1(n_3314),
.A2(n_3151),
.B(n_3259),
.Y(n_3623)
);

AOI21x1_ASAP7_75t_L g3624 ( 
.A1(n_3433),
.A2(n_2985),
.B(n_3183),
.Y(n_3624)
);

OAI21x1_ASAP7_75t_L g3625 ( 
.A1(n_3342),
.A2(n_3151),
.B(n_3259),
.Y(n_3625)
);

OAI21x1_ASAP7_75t_L g3626 ( 
.A1(n_3374),
.A2(n_3197),
.B(n_3213),
.Y(n_3626)
);

AOI221xp5_ASAP7_75t_L g3627 ( 
.A1(n_3375),
.A2(n_3147),
.B1(n_3176),
.B2(n_3032),
.C(n_2987),
.Y(n_3627)
);

AND2x2_ASAP7_75t_SL g3628 ( 
.A(n_3473),
.B(n_3246),
.Y(n_3628)
);

AO21x2_ASAP7_75t_L g3629 ( 
.A1(n_3529),
.A2(n_3203),
.B(n_3145),
.Y(n_3629)
);

NAND3xp33_ASAP7_75t_L g3630 ( 
.A(n_3469),
.B(n_3301),
.C(n_3603),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3280),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3281),
.Y(n_3632)
);

AND2x4_ASAP7_75t_L g3633 ( 
.A(n_3565),
.B(n_2949),
.Y(n_3633)
);

NAND3xp33_ASAP7_75t_L g3634 ( 
.A(n_3311),
.B(n_3613),
.C(n_3357),
.Y(n_3634)
);

HB1xp67_ASAP7_75t_L g3635 ( 
.A(n_3305),
.Y(n_3635)
);

INVx1_ASAP7_75t_SL g3636 ( 
.A(n_3406),
.Y(n_3636)
);

OAI21x1_ASAP7_75t_L g3637 ( 
.A1(n_3433),
.A2(n_3197),
.B(n_3213),
.Y(n_3637)
);

HB1xp67_ASAP7_75t_L g3638 ( 
.A(n_3292),
.Y(n_3638)
);

INVx2_ASAP7_75t_L g3639 ( 
.A(n_3379),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3439),
.Y(n_3640)
);

OAI21x1_ASAP7_75t_L g3641 ( 
.A1(n_3427),
.A2(n_3138),
.B(n_3135),
.Y(n_3641)
);

OAI21xp5_ASAP7_75t_L g3642 ( 
.A1(n_3367),
.A2(n_2861),
.B(n_3116),
.Y(n_3642)
);

A2O1A1Ixp33_ASAP7_75t_L g3643 ( 
.A1(n_3291),
.A2(n_3246),
.B(n_3228),
.C(n_3075),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3391),
.Y(n_3644)
);

INVx1_ASAP7_75t_SL g3645 ( 
.A(n_3423),
.Y(n_3645)
);

OAI21x1_ASAP7_75t_L g3646 ( 
.A1(n_3480),
.A2(n_3138),
.B(n_3135),
.Y(n_3646)
);

BUFx12f_ASAP7_75t_L g3647 ( 
.A(n_3318),
.Y(n_3647)
);

CKINVDCx20_ASAP7_75t_R g3648 ( 
.A(n_3302),
.Y(n_3648)
);

OR2x2_ASAP7_75t_L g3649 ( 
.A(n_3290),
.B(n_3059),
.Y(n_3649)
);

OAI21x1_ASAP7_75t_L g3650 ( 
.A1(n_3486),
.A2(n_3107),
.B(n_3019),
.Y(n_3650)
);

AOI221xp5_ASAP7_75t_L g3651 ( 
.A1(n_3286),
.A2(n_3097),
.B1(n_2953),
.B2(n_2973),
.C(n_3178),
.Y(n_3651)
);

NOR2xp67_ASAP7_75t_L g3652 ( 
.A(n_3329),
.B(n_3019),
.Y(n_3652)
);

AOI21x1_ASAP7_75t_L g3653 ( 
.A1(n_3501),
.A2(n_3241),
.B(n_3239),
.Y(n_3653)
);

INVx3_ASAP7_75t_L g3654 ( 
.A(n_3329),
.Y(n_3654)
);

INVx1_ASAP7_75t_SL g3655 ( 
.A(n_3438),
.Y(n_3655)
);

OAI21x1_ASAP7_75t_L g3656 ( 
.A1(n_3502),
.A2(n_3107),
.B(n_3204),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3288),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3393),
.Y(n_3658)
);

NAND2x1p5_ASAP7_75t_L g3659 ( 
.A(n_3310),
.B(n_3228),
.Y(n_3659)
);

AOI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3371),
.A2(n_2891),
.B1(n_2907),
.B2(n_3122),
.Y(n_3660)
);

HB1xp67_ASAP7_75t_L g3661 ( 
.A(n_3400),
.Y(n_3661)
);

AOI221xp5_ASAP7_75t_L g3662 ( 
.A1(n_3316),
.A2(n_3002),
.B1(n_3155),
.B2(n_3154),
.C(n_3139),
.Y(n_3662)
);

OAI21x1_ASAP7_75t_L g3663 ( 
.A1(n_3294),
.A2(n_3243),
.B(n_3126),
.Y(n_3663)
);

OA21x2_ASAP7_75t_L g3664 ( 
.A1(n_3426),
.A2(n_2895),
.B(n_3120),
.Y(n_3664)
);

NOR2xp33_ASAP7_75t_L g3665 ( 
.A(n_3600),
.B(n_2946),
.Y(n_3665)
);

INVx2_ASAP7_75t_SL g3666 ( 
.A(n_3328),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3325),
.A2(n_3044),
.B(n_3005),
.Y(n_3667)
);

NAND2x1p5_ASAP7_75t_L g3668 ( 
.A(n_3330),
.B(n_3372),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3289),
.Y(n_3669)
);

AOI221xp5_ASAP7_75t_L g3670 ( 
.A1(n_3553),
.A2(n_3164),
.B1(n_3200),
.B2(n_3195),
.C(n_3177),
.Y(n_3670)
);

INVx3_ASAP7_75t_L g3671 ( 
.A(n_3329),
.Y(n_3671)
);

INVx2_ASAP7_75t_L g3672 ( 
.A(n_3412),
.Y(n_3672)
);

OAI21x1_ASAP7_75t_L g3673 ( 
.A1(n_3514),
.A2(n_3123),
.B(n_3134),
.Y(n_3673)
);

OAI22xp5_ASAP7_75t_L g3674 ( 
.A1(n_3565),
.A2(n_2879),
.B1(n_2936),
.B2(n_3056),
.Y(n_3674)
);

NAND2x1p5_ASAP7_75t_L g3675 ( 
.A(n_3378),
.B(n_3236),
.Y(n_3675)
);

BUFx4_ASAP7_75t_R g3676 ( 
.A(n_3481),
.Y(n_3676)
);

CKINVDCx20_ASAP7_75t_R g3677 ( 
.A(n_3411),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3431),
.Y(n_3678)
);

INVx3_ASAP7_75t_L g3679 ( 
.A(n_3380),
.Y(n_3679)
);

NOR2xp67_ASAP7_75t_SL g3680 ( 
.A(n_3380),
.B(n_3436),
.Y(n_3680)
);

INVx3_ASAP7_75t_L g3681 ( 
.A(n_3380),
.Y(n_3681)
);

NAND2x1p5_ASAP7_75t_L g3682 ( 
.A(n_3296),
.B(n_3236),
.Y(n_3682)
);

INVx2_ASAP7_75t_L g3683 ( 
.A(n_3446),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3451),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_3474),
.B(n_3053),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3496),
.A2(n_2888),
.B(n_2887),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3461),
.B(n_3062),
.Y(n_3687)
);

BUFx3_ASAP7_75t_L g3688 ( 
.A(n_3401),
.Y(n_3688)
);

AO21x2_ASAP7_75t_L g3689 ( 
.A1(n_3591),
.A2(n_3076),
.B(n_2921),
.Y(n_3689)
);

AOI22xp33_ASAP7_75t_L g3690 ( 
.A1(n_3363),
.A2(n_3146),
.B1(n_3127),
.B2(n_3209),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3459),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3300),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3283),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3306),
.Y(n_3694)
);

INVx6_ASAP7_75t_SL g3695 ( 
.A(n_3363),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_3313),
.B(n_3003),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3364),
.B(n_3073),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3366),
.Y(n_3698)
);

BUFx2_ASAP7_75t_L g3699 ( 
.A(n_3507),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3376),
.Y(n_3700)
);

OA21x2_ASAP7_75t_L g3701 ( 
.A1(n_3418),
.A2(n_2901),
.B(n_2898),
.Y(n_3701)
);

AO21x2_ASAP7_75t_L g3702 ( 
.A1(n_3303),
.A2(n_2998),
.B(n_2892),
.Y(n_3702)
);

OAI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_3399),
.A2(n_3021),
.B(n_3227),
.Y(n_3703)
);

AND2x4_ASAP7_75t_L g3704 ( 
.A(n_3436),
.B(n_3005),
.Y(n_3704)
);

NAND2x1p5_ASAP7_75t_L g3705 ( 
.A(n_3274),
.B(n_3044),
.Y(n_3705)
);

INVx3_ASAP7_75t_L g3706 ( 
.A(n_3436),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3381),
.Y(n_3707)
);

BUFx2_ASAP7_75t_R g3708 ( 
.A(n_3273),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3285),
.Y(n_3709)
);

HB1xp67_ASAP7_75t_L g3710 ( 
.A(n_3532),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3390),
.Y(n_3711)
);

OAI21x1_ASAP7_75t_L g3712 ( 
.A1(n_3414),
.A2(n_3159),
.B(n_3162),
.Y(n_3712)
);

AND2x4_ASAP7_75t_L g3713 ( 
.A(n_3561),
.B(n_3044),
.Y(n_3713)
);

NOR2xp33_ASAP7_75t_SL g3714 ( 
.A(n_3509),
.B(n_3065),
.Y(n_3714)
);

O2A1O1Ixp33_ASAP7_75t_SL g3715 ( 
.A1(n_3505),
.A2(n_2943),
.B(n_2942),
.C(n_3110),
.Y(n_3715)
);

OAI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_3322),
.A2(n_3235),
.B(n_3232),
.Y(n_3716)
);

OAI21x1_ASAP7_75t_L g3717 ( 
.A1(n_3472),
.A2(n_3193),
.B(n_3185),
.Y(n_3717)
);

OR2x2_ASAP7_75t_L g3718 ( 
.A(n_3563),
.B(n_3206),
.Y(n_3718)
);

OAI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3355),
.A2(n_3254),
.B(n_3251),
.Y(n_3719)
);

NOR3xp33_ASAP7_75t_SL g3720 ( 
.A(n_3333),
.B(n_3217),
.C(n_3218),
.Y(n_3720)
);

OAI21x1_ASAP7_75t_L g3721 ( 
.A1(n_3454),
.A2(n_3382),
.B(n_3319),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3398),
.Y(n_3722)
);

AOI21x1_ASAP7_75t_L g3723 ( 
.A1(n_3501),
.A2(n_3114),
.B(n_3263),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_3416),
.B(n_2910),
.Y(n_3724)
);

INVx1_ASAP7_75t_SL g3725 ( 
.A(n_3401),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3419),
.Y(n_3726)
);

OAI21x1_ASAP7_75t_L g3727 ( 
.A1(n_3307),
.A2(n_3210),
.B(n_2948),
.Y(n_3727)
);

AO31x2_ASAP7_75t_L g3728 ( 
.A1(n_3327),
.A2(n_2951),
.A3(n_2917),
.B(n_2857),
.Y(n_3728)
);

OAI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_3276),
.A2(n_3042),
.B(n_2967),
.Y(n_3729)
);

AOI22xp33_ASAP7_75t_SL g3730 ( 
.A1(n_3617),
.A2(n_2863),
.B1(n_2867),
.B2(n_2856),
.Y(n_3730)
);

BUFx10_ASAP7_75t_L g3731 ( 
.A(n_3277),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_SL g3732 ( 
.A1(n_3457),
.A2(n_3109),
.B1(n_2870),
.B2(n_2878),
.Y(n_3732)
);

INVxp67_ASAP7_75t_L g3733 ( 
.A(n_3584),
.Y(n_3733)
);

OAI21x1_ASAP7_75t_L g3734 ( 
.A1(n_3320),
.A2(n_2884),
.B(n_2869),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3425),
.B(n_3071),
.Y(n_3735)
);

OA21x2_ASAP7_75t_L g3736 ( 
.A1(n_3327),
.A2(n_3077),
.B(n_3068),
.Y(n_3736)
);

OAI21x1_ASAP7_75t_L g3737 ( 
.A1(n_3335),
.A2(n_3086),
.B(n_3080),
.Y(n_3737)
);

OAI21x1_ASAP7_75t_L g3738 ( 
.A1(n_3339),
.A2(n_3090),
.B(n_3070),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3428),
.Y(n_3739)
);

AO21x2_ASAP7_75t_L g3740 ( 
.A1(n_3395),
.A2(n_3070),
.B(n_3065),
.Y(n_3740)
);

BUFx3_ASAP7_75t_L g3741 ( 
.A(n_3334),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3359),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3437),
.B(n_3065),
.Y(n_3743)
);

OAI21x1_ASAP7_75t_L g3744 ( 
.A1(n_3323),
.A2(n_3121),
.B(n_3070),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3533),
.Y(n_3745)
);

AND2x2_ASAP7_75t_L g3746 ( 
.A(n_3504),
.B(n_337),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3453),
.B(n_3121),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3543),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3556),
.Y(n_3749)
);

OAI221xp5_ASAP7_75t_L g3750 ( 
.A1(n_3498),
.A2(n_3133),
.B1(n_3137),
.B2(n_3125),
.C(n_3121),
.Y(n_3750)
);

AOI21xp5_ASAP7_75t_L g3751 ( 
.A1(n_3488),
.A2(n_3133),
.B(n_3125),
.Y(n_3751)
);

INVx4_ASAP7_75t_L g3752 ( 
.A(n_3445),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_L g3753 ( 
.A1(n_3340),
.A2(n_3133),
.B(n_3125),
.Y(n_3753)
);

OAI21x1_ASAP7_75t_L g3754 ( 
.A1(n_3599),
.A2(n_3174),
.B(n_3137),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3458),
.Y(n_3755)
);

AO21x2_ASAP7_75t_L g3756 ( 
.A1(n_3601),
.A2(n_3174),
.B(n_3137),
.Y(n_3756)
);

BUFx2_ASAP7_75t_L g3757 ( 
.A(n_3572),
.Y(n_3757)
);

AND2x2_ASAP7_75t_SL g3758 ( 
.A(n_3554),
.B(n_3174),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3575),
.Y(n_3759)
);

BUFx2_ASAP7_75t_L g3760 ( 
.A(n_3616),
.Y(n_3760)
);

OAI21x1_ASAP7_75t_L g3761 ( 
.A1(n_3490),
.A2(n_3238),
.B(n_3229),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3478),
.B(n_3517),
.Y(n_3762)
);

NOR2xp33_ASAP7_75t_SL g3763 ( 
.A(n_3523),
.B(n_3229),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3586),
.Y(n_3764)
);

OAI22xp5_ASAP7_75t_L g3765 ( 
.A1(n_3526),
.A2(n_3238),
.B1(n_3229),
.B2(n_340),
.Y(n_3765)
);

OAI21x1_ASAP7_75t_L g3766 ( 
.A1(n_3503),
.A2(n_3238),
.B(n_730),
.Y(n_3766)
);

OR2x2_ASAP7_75t_L g3767 ( 
.A(n_3470),
.B(n_338),
.Y(n_3767)
);

BUFx3_ASAP7_75t_L g3768 ( 
.A(n_3349),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3521),
.Y(n_3769)
);

AO21x1_ASAP7_75t_L g3770 ( 
.A1(n_3583),
.A2(n_338),
.B(n_339),
.Y(n_3770)
);

AOI21x1_ASAP7_75t_L g3771 ( 
.A1(n_3370),
.A2(n_3368),
.B(n_3356),
.Y(n_3771)
);

AOI22xp5_ASAP7_75t_L g3772 ( 
.A1(n_3526),
.A2(n_342),
.B1(n_339),
.B2(n_341),
.Y(n_3772)
);

NOR2xp33_ASAP7_75t_L g3773 ( 
.A(n_3440),
.B(n_342),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3487),
.Y(n_3774)
);

CKINVDCx20_ASAP7_75t_R g3775 ( 
.A(n_3441),
.Y(n_3775)
);

OAI21xp5_ASAP7_75t_L g3776 ( 
.A1(n_3551),
.A2(n_343),
.B(n_344),
.Y(n_3776)
);

INVx6_ASAP7_75t_L g3777 ( 
.A(n_3404),
.Y(n_3777)
);

NAND2x1p5_ASAP7_75t_L g3778 ( 
.A(n_3309),
.B(n_3331),
.Y(n_3778)
);

AOI22xp5_ASAP7_75t_L g3779 ( 
.A1(n_3545),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_3779)
);

BUFx12f_ASAP7_75t_L g3780 ( 
.A(n_3383),
.Y(n_3780)
);

OAI21x1_ASAP7_75t_L g3781 ( 
.A1(n_3518),
.A2(n_732),
.B(n_729),
.Y(n_3781)
);

BUFx2_ASAP7_75t_R g3782 ( 
.A(n_3388),
.Y(n_3782)
);

HB1xp67_ASAP7_75t_L g3783 ( 
.A(n_3522),
.Y(n_3783)
);

AO21x2_ASAP7_75t_L g3784 ( 
.A1(n_3332),
.A2(n_345),
.B(n_346),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3524),
.B(n_346),
.Y(n_3785)
);

INVx1_ASAP7_75t_SL g3786 ( 
.A(n_3452),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3479),
.Y(n_3787)
);

NOR2x1_ASAP7_75t_R g3788 ( 
.A(n_3338),
.B(n_347),
.Y(n_3788)
);

AO22x1_ASAP7_75t_L g3789 ( 
.A1(n_3561),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_3789)
);

OAI21x1_ASAP7_75t_L g3790 ( 
.A1(n_3525),
.A2(n_736),
.B(n_733),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3568),
.B(n_348),
.Y(n_3791)
);

OAI21x1_ASAP7_75t_L g3792 ( 
.A1(n_3508),
.A2(n_740),
.B(n_739),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3315),
.B(n_349),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3513),
.Y(n_3794)
);

OAI21x1_ASAP7_75t_L g3795 ( 
.A1(n_3520),
.A2(n_742),
.B(n_741),
.Y(n_3795)
);

INVx6_ASAP7_75t_L g3796 ( 
.A(n_3331),
.Y(n_3796)
);

OAI21xp5_ASAP7_75t_L g3797 ( 
.A1(n_3324),
.A2(n_350),
.B(n_351),
.Y(n_3797)
);

OAI21x1_ASAP7_75t_L g3798 ( 
.A1(n_3559),
.A2(n_744),
.B(n_743),
.Y(n_3798)
);

OAI21x1_ASAP7_75t_L g3799 ( 
.A1(n_3564),
.A2(n_747),
.B(n_746),
.Y(n_3799)
);

OAI21x1_ASAP7_75t_SL g3800 ( 
.A1(n_3465),
.A2(n_351),
.B(n_352),
.Y(n_3800)
);

OAI21x1_ASAP7_75t_L g3801 ( 
.A1(n_3569),
.A2(n_3573),
.B(n_3515),
.Y(n_3801)
);

BUFx2_ASAP7_75t_L g3802 ( 
.A(n_3445),
.Y(n_3802)
);

INVx2_ASAP7_75t_L g3803 ( 
.A(n_3337),
.Y(n_3803)
);

INVx1_ASAP7_75t_SL g3804 ( 
.A(n_3475),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3347),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3534),
.Y(n_3806)
);

CKINVDCx6p67_ASAP7_75t_R g3807 ( 
.A(n_3336),
.Y(n_3807)
);

OAI21x1_ASAP7_75t_L g3808 ( 
.A1(n_3495),
.A2(n_752),
.B(n_751),
.Y(n_3808)
);

OA21x2_ASAP7_75t_L g3809 ( 
.A1(n_3356),
.A2(n_756),
.B(n_754),
.Y(n_3809)
);

AOI31xp33_ASAP7_75t_L g3810 ( 
.A1(n_3304),
.A2(n_355),
.A3(n_353),
.B(n_354),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3549),
.Y(n_3811)
);

AND2x4_ASAP7_75t_L g3812 ( 
.A(n_3561),
.B(n_353),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3574),
.Y(n_3813)
);

AND2x4_ASAP7_75t_SL g3814 ( 
.A(n_3336),
.B(n_354),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3579),
.Y(n_3815)
);

OA21x2_ASAP7_75t_L g3816 ( 
.A1(n_3373),
.A2(n_760),
.B(n_757),
.Y(n_3816)
);

AOI21x1_ASAP7_75t_L g3817 ( 
.A1(n_3368),
.A2(n_762),
.B(n_761),
.Y(n_3817)
);

OAI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3354),
.A2(n_355),
.B(n_356),
.Y(n_3818)
);

AOI21xp5_ASAP7_75t_L g3819 ( 
.A1(n_3488),
.A2(n_769),
.B(n_768),
.Y(n_3819)
);

OAI21x1_ASAP7_75t_L g3820 ( 
.A1(n_3429),
.A2(n_772),
.B(n_770),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3587),
.Y(n_3821)
);

OAI21x1_ASAP7_75t_L g3822 ( 
.A1(n_3432),
.A2(n_778),
.B(n_776),
.Y(n_3822)
);

NOR2xp67_ASAP7_75t_L g3823 ( 
.A(n_3552),
.B(n_356),
.Y(n_3823)
);

NAND2x1_ASAP7_75t_L g3824 ( 
.A(n_3373),
.B(n_3445),
.Y(n_3824)
);

AOI21xp5_ASAP7_75t_L g3825 ( 
.A1(n_3548),
.A2(n_780),
.B(n_779),
.Y(n_3825)
);

NOR2xp33_ASAP7_75t_L g3826 ( 
.A(n_3510),
.B(n_357),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_L g3827 ( 
.A1(n_3583),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_3827)
);

AO21x2_ASAP7_75t_L g3828 ( 
.A1(n_3407),
.A2(n_358),
.B(n_359),
.Y(n_3828)
);

INVx4_ASAP7_75t_L g3829 ( 
.A(n_3499),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3547),
.B(n_361),
.Y(n_3830)
);

OAI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_3537),
.A2(n_361),
.B(n_362),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3439),
.Y(n_3832)
);

OAI21x1_ASAP7_75t_L g3833 ( 
.A1(n_3588),
.A2(n_783),
.B(n_782),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3589),
.Y(n_3834)
);

OAI21x1_ASAP7_75t_SL g3835 ( 
.A1(n_3604),
.A2(n_362),
.B(n_364),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3595),
.Y(n_3836)
);

BUFx6f_ASAP7_75t_L g3837 ( 
.A(n_3348),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3610),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3476),
.Y(n_3839)
);

OAI21x1_ASAP7_75t_L g3840 ( 
.A1(n_3596),
.A2(n_785),
.B(n_784),
.Y(n_3840)
);

INVx4_ASAP7_75t_L g3841 ( 
.A(n_3499),
.Y(n_3841)
);

O2A1O1Ixp33_ASAP7_75t_L g3842 ( 
.A1(n_3272),
.A2(n_366),
.B(n_364),
.C(n_365),
.Y(n_3842)
);

NOR2xp67_ASAP7_75t_L g3843 ( 
.A(n_3506),
.B(n_365),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3544),
.B(n_367),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3410),
.Y(n_3845)
);

OAI21x1_ASAP7_75t_L g3846 ( 
.A1(n_3606),
.A2(n_787),
.B(n_786),
.Y(n_3846)
);

BUFx3_ASAP7_75t_L g3847 ( 
.A(n_3389),
.Y(n_3847)
);

BUFx2_ASAP7_75t_L g3848 ( 
.A(n_3499),
.Y(n_3848)
);

OA21x2_ASAP7_75t_L g3849 ( 
.A1(n_3408),
.A2(n_792),
.B(n_791),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3312),
.Y(n_3850)
);

OAI21x1_ASAP7_75t_L g3851 ( 
.A1(n_3612),
.A2(n_796),
.B(n_795),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3410),
.Y(n_3852)
);

CKINVDCx5p33_ASAP7_75t_R g3853 ( 
.A(n_3477),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3444),
.Y(n_3854)
);

BUFx2_ASAP7_75t_L g3855 ( 
.A(n_3396),
.Y(n_3855)
);

HB1xp67_ASAP7_75t_L g3856 ( 
.A(n_3435),
.Y(n_3856)
);

OR2x2_ASAP7_75t_L g3857 ( 
.A(n_3541),
.B(n_367),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3491),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3444),
.Y(n_3859)
);

HB1xp67_ASAP7_75t_L g3860 ( 
.A(n_3527),
.Y(n_3860)
);

A2O1A1Ixp33_ASAP7_75t_L g3861 ( 
.A1(n_3597),
.A2(n_370),
.B(n_368),
.C(n_369),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3293),
.B(n_368),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3614),
.Y(n_3863)
);

OAI21xp5_ASAP7_75t_L g3864 ( 
.A1(n_3420),
.A2(n_369),
.B(n_370),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3578),
.Y(n_3865)
);

OAI21x1_ASAP7_75t_SL g3866 ( 
.A1(n_3511),
.A2(n_371),
.B(n_372),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3448),
.Y(n_3867)
);

INVx4_ASAP7_75t_L g3868 ( 
.A(n_3348),
.Y(n_3868)
);

OA21x2_ASAP7_75t_L g3869 ( 
.A1(n_3555),
.A2(n_800),
.B(n_799),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3447),
.B(n_372),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3448),
.Y(n_3871)
);

AND2x4_ASAP7_75t_L g3872 ( 
.A(n_3284),
.B(n_373),
.Y(n_3872)
);

NOR2xp33_ASAP7_75t_L g3873 ( 
.A(n_3422),
.B(n_373),
.Y(n_3873)
);

OAI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3512),
.A2(n_374),
.B(n_375),
.Y(n_3874)
);

HB1xp67_ASAP7_75t_L g3875 ( 
.A(n_3560),
.Y(n_3875)
);

BUFx2_ASAP7_75t_L g3876 ( 
.A(n_3396),
.Y(n_3876)
);

AND3x1_ASAP7_75t_L g3877 ( 
.A(n_3484),
.B(n_374),
.C(n_376),
.Y(n_3877)
);

BUFx8_ASAP7_75t_L g3878 ( 
.A(n_3409),
.Y(n_3878)
);

AND2x4_ASAP7_75t_L g3879 ( 
.A(n_3284),
.B(n_376),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3608),
.B(n_377),
.Y(n_3880)
);

INVxp67_ASAP7_75t_SL g3881 ( 
.A(n_3397),
.Y(n_3881)
);

OA21x2_ASAP7_75t_L g3882 ( 
.A1(n_3341),
.A2(n_807),
.B(n_806),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3605),
.Y(n_3883)
);

OA21x2_ASAP7_75t_L g3884 ( 
.A1(n_3397),
.A2(n_3430),
.B(n_3442),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3615),
.Y(n_3885)
);

NAND2x1p5_ASAP7_75t_L g3886 ( 
.A(n_3377),
.B(n_377),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_3468),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3468),
.Y(n_3888)
);

OAI21x1_ASAP7_75t_L g3889 ( 
.A1(n_3424),
.A2(n_809),
.B(n_808),
.Y(n_3889)
);

OA21x2_ASAP7_75t_L g3890 ( 
.A1(n_3430),
.A2(n_812),
.B(n_811),
.Y(n_3890)
);

HB1xp67_ASAP7_75t_L g3891 ( 
.A(n_3611),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3350),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3287),
.Y(n_3893)
);

INVxp67_ASAP7_75t_L g3894 ( 
.A(n_3545),
.Y(n_3894)
);

A2O1A1Ixp33_ASAP7_75t_L g3895 ( 
.A1(n_3576),
.A2(n_380),
.B(n_378),
.C(n_379),
.Y(n_3895)
);

OR2x6_ASAP7_75t_L g3896 ( 
.A(n_3607),
.B(n_379),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3494),
.Y(n_3897)
);

INVx1_ASAP7_75t_SL g3898 ( 
.A(n_3562),
.Y(n_3898)
);

AO21x2_ASAP7_75t_L g3899 ( 
.A1(n_3443),
.A2(n_381),
.B(n_382),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3538),
.Y(n_3900)
);

OAI22xp5_ASAP7_75t_SL g3901 ( 
.A1(n_3775),
.A2(n_3463),
.B1(n_3385),
.B2(n_3392),
.Y(n_3901)
);

OAI21x1_ASAP7_75t_L g3902 ( 
.A1(n_3625),
.A2(n_3751),
.B(n_3623),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3693),
.Y(n_3903)
);

CKINVDCx5p33_ASAP7_75t_R g3904 ( 
.A(n_3677),
.Y(n_3904)
);

INVx6_ASAP7_75t_L g3905 ( 
.A(n_3878),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3709),
.Y(n_3906)
);

AOI22xp33_ASAP7_75t_L g3907 ( 
.A1(n_3630),
.A2(n_3352),
.B1(n_3542),
.B2(n_3558),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3631),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3863),
.B(n_3592),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_3742),
.Y(n_3910)
);

INVx6_ASAP7_75t_L g3911 ( 
.A(n_3878),
.Y(n_3911)
);

NAND2xp33_ASAP7_75t_R g3912 ( 
.A(n_3757),
.B(n_3760),
.Y(n_3912)
);

AND2x4_ASAP7_75t_L g3913 ( 
.A(n_3881),
.B(n_3362),
.Y(n_3913)
);

AOI221xp5_ASAP7_75t_L g3914 ( 
.A1(n_3810),
.A2(n_3528),
.B1(n_3492),
.B2(n_3602),
.C(n_3550),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_L g3915 ( 
.A1(n_3634),
.A2(n_3299),
.B1(n_3317),
.B2(n_3326),
.Y(n_3915)
);

OAI22xp5_ASAP7_75t_L g3916 ( 
.A1(n_3628),
.A2(n_3617),
.B1(n_3609),
.B2(n_3535),
.Y(n_3916)
);

NAND2xp33_ASAP7_75t_R g3917 ( 
.A(n_3699),
.B(n_3275),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3632),
.Y(n_3918)
);

AOI22xp33_ASAP7_75t_L g3919 ( 
.A1(n_3674),
.A2(n_3345),
.B1(n_3566),
.B2(n_3570),
.Y(n_3919)
);

AOI221xp5_ASAP7_75t_L g3920 ( 
.A1(n_3670),
.A2(n_3394),
.B1(n_3386),
.B2(n_3530),
.C(n_3298),
.Y(n_3920)
);

OAI22xp33_ASAP7_75t_L g3921 ( 
.A1(n_3896),
.A2(n_3360),
.B1(n_3516),
.B2(n_3546),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3893),
.B(n_3415),
.Y(n_3922)
);

AOI221xp5_ASAP7_75t_L g3923 ( 
.A1(n_3877),
.A2(n_3402),
.B1(n_3413),
.B2(n_3361),
.C(n_3531),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3657),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_3803),
.B(n_3321),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3687),
.B(n_3403),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3669),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3692),
.Y(n_3928)
);

AOI22xp33_ASAP7_75t_SL g3929 ( 
.A1(n_3872),
.A2(n_3369),
.B1(n_3350),
.B2(n_3360),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3694),
.Y(n_3930)
);

NAND2x1_ASAP7_75t_L g3931 ( 
.A(n_3680),
.B(n_3752),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3698),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3700),
.Y(n_3933)
);

AND2x4_ASAP7_75t_L g3934 ( 
.A(n_3847),
.B(n_3585),
.Y(n_3934)
);

AOI21xp5_ASAP7_75t_L g3935 ( 
.A1(n_3643),
.A2(n_3417),
.B(n_3442),
.Y(n_3935)
);

AND2x4_ASAP7_75t_L g3936 ( 
.A(n_3633),
.B(n_3598),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3707),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3685),
.B(n_3464),
.Y(n_3938)
);

OAI22xp33_ASAP7_75t_L g3939 ( 
.A1(n_3896),
.A2(n_3818),
.B1(n_3695),
.B2(n_3864),
.Y(n_3939)
);

INVx6_ASAP7_75t_L g3940 ( 
.A(n_3731),
.Y(n_3940)
);

OR2x2_ASAP7_75t_L g3941 ( 
.A(n_3635),
.B(n_3450),
.Y(n_3941)
);

AOI22xp33_ASAP7_75t_L g3942 ( 
.A1(n_3642),
.A2(n_3567),
.B1(n_3449),
.B2(n_3351),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3774),
.Y(n_3943)
);

AOI22xp5_ASAP7_75t_SL g3944 ( 
.A1(n_3768),
.A2(n_3369),
.B1(n_3308),
.B2(n_3384),
.Y(n_3944)
);

OAI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3695),
.A2(n_3421),
.B1(n_3493),
.B2(n_3365),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3711),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3805),
.B(n_3460),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3722),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3794),
.Y(n_3949)
);

OAI22xp5_ASAP7_75t_L g3950 ( 
.A1(n_3690),
.A2(n_3462),
.B1(n_3455),
.B2(n_3387),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3639),
.Y(n_3951)
);

AOI211xp5_ASAP7_75t_L g3952 ( 
.A1(n_3788),
.A2(n_3353),
.B(n_3344),
.C(n_3467),
.Y(n_3952)
);

OAI22xp5_ASAP7_75t_L g3953 ( 
.A1(n_3894),
.A2(n_3365),
.B1(n_3278),
.B2(n_3271),
.Y(n_3953)
);

AND2x2_ASAP7_75t_L g3954 ( 
.A(n_3891),
.B(n_3456),
.Y(n_3954)
);

AOI22xp33_ASAP7_75t_L g3955 ( 
.A1(n_3651),
.A2(n_3483),
.B1(n_3358),
.B2(n_3466),
.Y(n_3955)
);

AOI22xp33_ASAP7_75t_L g3956 ( 
.A1(n_3770),
.A2(n_3627),
.B1(n_3732),
.B2(n_3621),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3726),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3644),
.Y(n_3958)
);

INVx1_ASAP7_75t_SL g3959 ( 
.A(n_3777),
.Y(n_3959)
);

AOI211xp5_ASAP7_75t_L g3960 ( 
.A1(n_3826),
.A2(n_3482),
.B(n_3358),
.C(n_3295),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3739),
.Y(n_3961)
);

AOI22xp33_ASAP7_75t_SL g3962 ( 
.A1(n_3872),
.A2(n_3497),
.B1(n_3500),
.B2(n_3456),
.Y(n_3962)
);

OAI22xp5_ASAP7_75t_L g3963 ( 
.A1(n_3772),
.A2(n_3580),
.B1(n_3405),
.B2(n_3500),
.Y(n_3963)
);

AOI221xp5_ASAP7_75t_L g3964 ( 
.A1(n_3662),
.A2(n_3279),
.B1(n_3434),
.B2(n_3489),
.C(n_3485),
.Y(n_3964)
);

CKINVDCx5p33_ASAP7_75t_R g3965 ( 
.A(n_3648),
.Y(n_3965)
);

AOI22xp33_ASAP7_75t_L g3966 ( 
.A1(n_3879),
.A2(n_3497),
.B1(n_3571),
.B2(n_3540),
.Y(n_3966)
);

OAI21x1_ASAP7_75t_L g3967 ( 
.A1(n_3618),
.A2(n_3346),
.B(n_3580),
.Y(n_3967)
);

AOI22xp33_ASAP7_75t_L g3968 ( 
.A1(n_3879),
.A2(n_3571),
.B1(n_3582),
.B2(n_3540),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3658),
.Y(n_3969)
);

BUFx3_ASAP7_75t_L g3970 ( 
.A(n_3777),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3672),
.Y(n_3971)
);

INVx6_ASAP7_75t_L g3972 ( 
.A(n_3731),
.Y(n_3972)
);

AND2x4_ASAP7_75t_L g3973 ( 
.A(n_3633),
.B(n_3582),
.Y(n_3973)
);

AND2x2_ASAP7_75t_L g3974 ( 
.A(n_3718),
.B(n_3638),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3755),
.Y(n_3975)
);

BUFx8_ASAP7_75t_SL g3976 ( 
.A(n_3647),
.Y(n_3976)
);

INVx2_ASAP7_75t_L g3977 ( 
.A(n_3678),
.Y(n_3977)
);

AOI22xp33_ASAP7_75t_L g3978 ( 
.A1(n_3729),
.A2(n_3594),
.B1(n_3580),
.B2(n_3519),
.Y(n_3978)
);

HB1xp67_ASAP7_75t_L g3979 ( 
.A(n_3661),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_SL g3980 ( 
.A(n_3758),
.B(n_3471),
.Y(n_3980)
);

INVx4_ASAP7_75t_SL g3981 ( 
.A(n_3812),
.Y(n_3981)
);

AOI22xp33_ASAP7_75t_L g3982 ( 
.A1(n_3797),
.A2(n_3594),
.B1(n_3519),
.B2(n_3536),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_3715),
.A2(n_3593),
.B(n_3536),
.Y(n_3983)
);

INVxp67_ASAP7_75t_SL g3984 ( 
.A(n_3710),
.Y(n_3984)
);

NAND3x1_ASAP7_75t_L g3985 ( 
.A(n_3773),
.B(n_381),
.C(n_382),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3806),
.B(n_3471),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_SL g3987 ( 
.A(n_3752),
.B(n_3593),
.Y(n_3987)
);

OA21x2_ASAP7_75t_L g3988 ( 
.A1(n_3637),
.A2(n_3557),
.B(n_3539),
.Y(n_3988)
);

AOI22xp33_ASAP7_75t_L g3989 ( 
.A1(n_3716),
.A2(n_3874),
.B1(n_3831),
.B2(n_3702),
.Y(n_3989)
);

BUFx6f_ASAP7_75t_L g3990 ( 
.A(n_3619),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3769),
.Y(n_3991)
);

OAI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3779),
.A2(n_3557),
.B1(n_3577),
.B2(n_3539),
.Y(n_3992)
);

BUFx6f_ASAP7_75t_L g3993 ( 
.A(n_3619),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3787),
.Y(n_3994)
);

AOI222xp33_ASAP7_75t_L g3995 ( 
.A1(n_3865),
.A2(n_385),
.B1(n_387),
.B2(n_383),
.C1(n_384),
.C2(n_386),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3815),
.B(n_3590),
.Y(n_3996)
);

AND2x4_ASAP7_75t_L g3997 ( 
.A(n_3868),
.B(n_3577),
.Y(n_3997)
);

INVx5_ASAP7_75t_L g3998 ( 
.A(n_3619),
.Y(n_3998)
);

OAI22xp5_ASAP7_75t_L g3999 ( 
.A1(n_3827),
.A2(n_3590),
.B1(n_3581),
.B2(n_385),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3683),
.Y(n_4000)
);

NAND2x1p5_ASAP7_75t_L g4001 ( 
.A(n_3666),
.B(n_3581),
.Y(n_4001)
);

OAI21x1_ASAP7_75t_SL g4002 ( 
.A1(n_3771),
.A2(n_383),
.B(n_384),
.Y(n_4002)
);

AOI21x1_ASAP7_75t_L g4003 ( 
.A1(n_3890),
.A2(n_387),
.B(n_388),
.Y(n_4003)
);

NAND3x1_ASAP7_75t_L g4004 ( 
.A(n_3676),
.B(n_388),
.C(n_389),
.Y(n_4004)
);

A2O1A1Ixp33_ASAP7_75t_L g4005 ( 
.A1(n_3843),
.A2(n_392),
.B(n_390),
.C(n_391),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3762),
.Y(n_4006)
);

OAI22xp33_ASAP7_75t_L g4007 ( 
.A1(n_3659),
.A2(n_395),
.B1(n_391),
.B2(n_394),
.Y(n_4007)
);

OR2x6_ASAP7_75t_L g4008 ( 
.A(n_3829),
.B(n_394),
.Y(n_4008)
);

AOI22xp5_ASAP7_75t_L g4009 ( 
.A1(n_3660),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_4009)
);

AOI22xp33_ASAP7_75t_L g4010 ( 
.A1(n_3689),
.A2(n_399),
.B1(n_396),
.B2(n_398),
.Y(n_4010)
);

AOI22xp33_ASAP7_75t_SL g4011 ( 
.A1(n_3855),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_4011)
);

BUFx6f_ASAP7_75t_SL g4012 ( 
.A(n_3622),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3801),
.Y(n_4013)
);

AO21x2_ASAP7_75t_L g4014 ( 
.A1(n_3800),
.A2(n_400),
.B(n_401),
.Y(n_4014)
);

CKINVDCx5p33_ASAP7_75t_R g4015 ( 
.A(n_3780),
.Y(n_4015)
);

HB1xp67_ASAP7_75t_L g4016 ( 
.A(n_3783),
.Y(n_4016)
);

OAI22xp5_ASAP7_75t_L g4017 ( 
.A1(n_3823),
.A2(n_405),
.B1(n_401),
.B2(n_402),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3850),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3811),
.B(n_402),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3856),
.B(n_406),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3813),
.B(n_3821),
.Y(n_4021)
);

NAND2x1_ASAP7_75t_L g4022 ( 
.A(n_3680),
.B(n_406),
.Y(n_4022)
);

OR2x2_ASAP7_75t_L g4023 ( 
.A(n_3640),
.B(n_407),
.Y(n_4023)
);

OAI22xp5_ASAP7_75t_L g4024 ( 
.A1(n_3861),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_4024)
);

AND2x4_ASAP7_75t_L g4025 ( 
.A(n_3868),
.B(n_408),
.Y(n_4025)
);

AO31x2_ASAP7_75t_L g4026 ( 
.A1(n_3892),
.A2(n_411),
.A3(n_409),
.B(n_410),
.Y(n_4026)
);

AOI22xp33_ASAP7_75t_L g4027 ( 
.A1(n_3800),
.A2(n_415),
.B1(n_413),
.B2(n_414),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3684),
.Y(n_4028)
);

CKINVDCx5p33_ASAP7_75t_R g4029 ( 
.A(n_3708),
.Y(n_4029)
);

OAI22xp5_ASAP7_75t_L g4030 ( 
.A1(n_3765),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_4030)
);

NAND3xp33_ASAP7_75t_L g4031 ( 
.A(n_3720),
.B(n_416),
.C(n_418),
.Y(n_4031)
);

CKINVDCx5p33_ASAP7_75t_R g4032 ( 
.A(n_3853),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3834),
.Y(n_4033)
);

CKINVDCx11_ASAP7_75t_R g4034 ( 
.A(n_3807),
.Y(n_4034)
);

AOI22xp33_ASAP7_75t_L g4035 ( 
.A1(n_3730),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3836),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3838),
.B(n_420),
.Y(n_4037)
);

OAI22xp5_ASAP7_75t_L g4038 ( 
.A1(n_3895),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_4038)
);

AND2x4_ASAP7_75t_L g4039 ( 
.A(n_3733),
.B(n_425),
.Y(n_4039)
);

AOI22xp33_ASAP7_75t_L g4040 ( 
.A1(n_3665),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_4040)
);

INVx3_ASAP7_75t_L g4041 ( 
.A(n_3668),
.Y(n_4041)
);

CKINVDCx16_ASAP7_75t_R g4042 ( 
.A(n_3688),
.Y(n_4042)
);

OAI221xp5_ASAP7_75t_L g4043 ( 
.A1(n_3886),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.C(n_430),
.Y(n_4043)
);

NAND2xp33_ASAP7_75t_SL g4044 ( 
.A(n_3824),
.B(n_429),
.Y(n_4044)
);

NAND2x1_ASAP7_75t_L g4045 ( 
.A(n_3829),
.B(n_431),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3860),
.Y(n_4046)
);

CKINVDCx8_ASAP7_75t_R g4047 ( 
.A(n_3620),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3691),
.Y(n_4048)
);

NOR2x1_ASAP7_75t_SL g4049 ( 
.A(n_3841),
.B(n_431),
.Y(n_4049)
);

NOR2xp33_ASAP7_75t_L g4050 ( 
.A(n_3636),
.B(n_432),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_3745),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3640),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3832),
.Y(n_4053)
);

INVx4_ASAP7_75t_L g4054 ( 
.A(n_3741),
.Y(n_4054)
);

BUFx4f_ASAP7_75t_L g4055 ( 
.A(n_3778),
.Y(n_4055)
);

NOR2xp33_ASAP7_75t_L g4056 ( 
.A(n_3645),
.B(n_433),
.Y(n_4056)
);

AOI22xp33_ASAP7_75t_L g4057 ( 
.A1(n_3784),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_4057)
);

AOI22xp33_ASAP7_75t_L g4058 ( 
.A1(n_3703),
.A2(n_437),
.B1(n_434),
.B2(n_435),
.Y(n_4058)
);

INVx3_ASAP7_75t_L g4059 ( 
.A(n_3620),
.Y(n_4059)
);

AOI22xp33_ASAP7_75t_L g4060 ( 
.A1(n_3746),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_4060)
);

OAI211xp5_ASAP7_75t_SL g4061 ( 
.A1(n_3883),
.A2(n_441),
.B(n_439),
.C(n_440),
.Y(n_4061)
);

OAI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_3842),
.A2(n_440),
.B(n_441),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_SL g4063 ( 
.A(n_3841),
.B(n_442),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3832),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3748),
.Y(n_4065)
);

AOI22xp5_ASAP7_75t_L g4066 ( 
.A1(n_3885),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3649),
.B(n_443),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_L g4068 ( 
.A1(n_3844),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3749),
.Y(n_4069)
);

AOI22xp33_ASAP7_75t_L g4070 ( 
.A1(n_3899),
.A2(n_448),
.B1(n_445),
.B2(n_447),
.Y(n_4070)
);

OR2x2_ASAP7_75t_L g4071 ( 
.A(n_3759),
.B(n_447),
.Y(n_4071)
);

AND2x4_ASAP7_75t_L g4072 ( 
.A(n_3876),
.B(n_448),
.Y(n_4072)
);

NAND2x1p5_ASAP7_75t_L g4073 ( 
.A(n_3655),
.B(n_3786),
.Y(n_4073)
);

OAI221xp5_ASAP7_75t_L g4074 ( 
.A1(n_3900),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.C(n_453),
.Y(n_4074)
);

INVxp67_ASAP7_75t_SL g4075 ( 
.A(n_3884),
.Y(n_4075)
);

OAI22xp5_ASAP7_75t_L g4076 ( 
.A1(n_3804),
.A2(n_455),
.B1(n_450),
.B2(n_454),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3764),
.Y(n_4077)
);

AOI221xp5_ASAP7_75t_L g4078 ( 
.A1(n_3897),
.A2(n_458),
.B1(n_454),
.B2(n_457),
.C(n_459),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_3839),
.B(n_457),
.Y(n_4079)
);

OAI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_3812),
.A2(n_3898),
.B1(n_3824),
.B2(n_3767),
.Y(n_4080)
);

AO21x2_ASAP7_75t_L g4081 ( 
.A1(n_3835),
.A2(n_459),
.B(n_460),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3875),
.Y(n_4082)
);

OAI22xp5_ASAP7_75t_L g4083 ( 
.A1(n_3802),
.A2(n_463),
.B1(n_460),
.B2(n_461),
.Y(n_4083)
);

INVx4_ASAP7_75t_L g4084 ( 
.A(n_3682),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_3870),
.B(n_463),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3743),
.Y(n_4086)
);

AOI21xp33_ASAP7_75t_L g4087 ( 
.A1(n_3701),
.A2(n_464),
.B(n_465),
.Y(n_4087)
);

AOI22xp33_ASAP7_75t_L g4088 ( 
.A1(n_3835),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3747),
.Y(n_4089)
);

AOI221xp5_ASAP7_75t_L g4090 ( 
.A1(n_3858),
.A2(n_3873),
.B1(n_3830),
.B2(n_3791),
.C(n_3880),
.Y(n_4090)
);

AOI22xp33_ASAP7_75t_L g4091 ( 
.A1(n_3866),
.A2(n_470),
.B1(n_466),
.B2(n_467),
.Y(n_4091)
);

AOI22xp33_ASAP7_75t_L g4092 ( 
.A1(n_3866),
.A2(n_3719),
.B1(n_3776),
.B2(n_3862),
.Y(n_4092)
);

BUFx6f_ASAP7_75t_L g4093 ( 
.A(n_3620),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4021),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3908),
.Y(n_4095)
);

CKINVDCx16_ASAP7_75t_R g4096 ( 
.A(n_3917),
.Y(n_4096)
);

AO31x2_ASAP7_75t_L g4097 ( 
.A1(n_4013),
.A2(n_3892),
.A3(n_3667),
.B(n_3819),
.Y(n_4097)
);

BUFx4f_ASAP7_75t_L g4098 ( 
.A(n_3905),
.Y(n_4098)
);

XOR2x2_ASAP7_75t_SL g4099 ( 
.A(n_4073),
.B(n_3675),
.Y(n_4099)
);

NOR2x1_ASAP7_75t_SL g4100 ( 
.A(n_4008),
.B(n_3771),
.Y(n_4100)
);

BUFx2_ASAP7_75t_L g4101 ( 
.A(n_3981),
.Y(n_4101)
);

CKINVDCx16_ASAP7_75t_R g4102 ( 
.A(n_4042),
.Y(n_4102)
);

BUFx12f_ASAP7_75t_L g4103 ( 
.A(n_4034),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3918),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_3974),
.B(n_3884),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_3954),
.B(n_3725),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_3938),
.B(n_3845),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_SL g4108 ( 
.A1(n_3944),
.A2(n_3848),
.B1(n_3890),
.B2(n_3814),
.Y(n_4108)
);

AOI22xp33_ASAP7_75t_SL g4109 ( 
.A1(n_4080),
.A2(n_3671),
.B1(n_3679),
.B2(n_3654),
.Y(n_4109)
);

A2O1A1Ixp33_ASAP7_75t_L g4110 ( 
.A1(n_3952),
.A2(n_4044),
.B(n_4031),
.C(n_3956),
.Y(n_4110)
);

AOI22xp33_ASAP7_75t_L g4111 ( 
.A1(n_3939),
.A2(n_3701),
.B1(n_3796),
.B2(n_3629),
.Y(n_4111)
);

NOR3xp33_ASAP7_75t_SL g4112 ( 
.A(n_4029),
.B(n_3750),
.C(n_3785),
.Y(n_4112)
);

AND2x4_ASAP7_75t_L g4113 ( 
.A(n_3981),
.B(n_3654),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3924),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_3927),
.Y(n_4115)
);

CKINVDCx16_ASAP7_75t_R g4116 ( 
.A(n_4012),
.Y(n_4116)
);

HB1xp67_ASAP7_75t_L g4117 ( 
.A(n_3979),
.Y(n_4117)
);

INVx3_ASAP7_75t_L g4118 ( 
.A(n_3905),
.Y(n_4118)
);

INVx2_ASAP7_75t_SL g4119 ( 
.A(n_3911),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3928),
.Y(n_4120)
);

OAI21xp33_ASAP7_75t_L g4121 ( 
.A1(n_3907),
.A2(n_3857),
.B(n_3793),
.Y(n_4121)
);

INVx2_ASAP7_75t_L g4122 ( 
.A(n_3903),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_3926),
.B(n_3852),
.Y(n_4123)
);

INVx2_ASAP7_75t_L g4124 ( 
.A(n_3906),
.Y(n_4124)
);

NAND2x1p5_ASAP7_75t_L g4125 ( 
.A(n_4055),
.B(n_3837),
.Y(n_4125)
);

INVx3_ASAP7_75t_SL g4126 ( 
.A(n_3911),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_3930),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_SL g4128 ( 
.A(n_3929),
.B(n_3837),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_3910),
.Y(n_4129)
);

NAND2xp33_ASAP7_75t_R g4130 ( 
.A(n_4041),
.B(n_3809),
.Y(n_4130)
);

CKINVDCx5p33_ASAP7_75t_R g4131 ( 
.A(n_3904),
.Y(n_4131)
);

OAI22xp5_ASAP7_75t_L g4132 ( 
.A1(n_3919),
.A2(n_3652),
.B1(n_3679),
.B2(n_3671),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3932),
.Y(n_4133)
);

NAND3xp33_ASAP7_75t_L g4134 ( 
.A(n_4090),
.B(n_3789),
.C(n_3724),
.Y(n_4134)
);

NOR3xp33_ASAP7_75t_SL g4135 ( 
.A(n_3945),
.B(n_3782),
.C(n_3697),
.Y(n_4135)
);

AND2x4_ASAP7_75t_L g4136 ( 
.A(n_3913),
.B(n_3681),
.Y(n_4136)
);

NAND2xp33_ASAP7_75t_SL g4137 ( 
.A(n_3912),
.B(n_3681),
.Y(n_4137)
);

NAND2xp33_ASAP7_75t_R g4138 ( 
.A(n_4008),
.B(n_3809),
.Y(n_4138)
);

AND2x2_ASAP7_75t_SL g4139 ( 
.A(n_4054),
.B(n_3816),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_3933),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3937),
.Y(n_4141)
);

AOI22xp33_ASAP7_75t_L g4142 ( 
.A1(n_3921),
.A2(n_3796),
.B1(n_3828),
.B2(n_3756),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_3951),
.Y(n_4143)
);

CKINVDCx5p33_ASAP7_75t_R g4144 ( 
.A(n_3976),
.Y(n_4144)
);

INVx2_ASAP7_75t_L g4145 ( 
.A(n_3958),
.Y(n_4145)
);

AND2x2_ASAP7_75t_L g4146 ( 
.A(n_4082),
.B(n_3854),
.Y(n_4146)
);

AND2x2_ASAP7_75t_L g4147 ( 
.A(n_4046),
.B(n_3859),
.Y(n_4147)
);

NOR2xp33_ASAP7_75t_R g4148 ( 
.A(n_4032),
.B(n_4015),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_4006),
.B(n_3728),
.Y(n_4149)
);

AOI22xp33_ASAP7_75t_L g4150 ( 
.A1(n_3915),
.A2(n_3736),
.B1(n_3849),
.B2(n_3816),
.Y(n_4150)
);

INVx1_ASAP7_75t_SL g4151 ( 
.A(n_3959),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_4016),
.B(n_3728),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3946),
.Y(n_4153)
);

AOI211xp5_ASAP7_75t_L g4154 ( 
.A1(n_3963),
.A2(n_3789),
.B(n_3714),
.C(n_3763),
.Y(n_4154)
);

OR2x6_ASAP7_75t_L g4155 ( 
.A(n_3931),
.B(n_3706),
.Y(n_4155)
);

INVx8_ASAP7_75t_L g4156 ( 
.A(n_3934),
.Y(n_4156)
);

BUFx6f_ASAP7_75t_L g4157 ( 
.A(n_4093),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_3984),
.B(n_3867),
.Y(n_4158)
);

NOR2xp33_ASAP7_75t_R g4159 ( 
.A(n_3940),
.B(n_3837),
.Y(n_4159)
);

BUFx2_ASAP7_75t_L g4160 ( 
.A(n_3970),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_4018),
.B(n_3871),
.Y(n_4161)
);

NOR2x1p5_ASAP7_75t_L g4162 ( 
.A(n_4045),
.B(n_3706),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_4086),
.B(n_3887),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3948),
.Y(n_4164)
);

CKINVDCx16_ASAP7_75t_R g4165 ( 
.A(n_3901),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_3957),
.B(n_3888),
.Y(n_4166)
);

CKINVDCx5p33_ASAP7_75t_R g4167 ( 
.A(n_3965),
.Y(n_4167)
);

AND2x2_ASAP7_75t_L g4168 ( 
.A(n_3961),
.B(n_3721),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_3975),
.Y(n_4169)
);

CKINVDCx5p33_ASAP7_75t_R g4170 ( 
.A(n_3940),
.Y(n_4170)
);

INVx5_ASAP7_75t_SL g4171 ( 
.A(n_4025),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3991),
.Y(n_4172)
);

CKINVDCx12_ASAP7_75t_R g4173 ( 
.A(n_3941),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_L g4174 ( 
.A1(n_3916),
.A2(n_3736),
.B1(n_3849),
.B2(n_3686),
.Y(n_4174)
);

HB1xp67_ASAP7_75t_L g4175 ( 
.A(n_3947),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_3969),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3994),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4033),
.Y(n_4178)
);

INVx4_ASAP7_75t_L g4179 ( 
.A(n_3972),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4036),
.Y(n_4180)
);

CKINVDCx5p33_ASAP7_75t_R g4181 ( 
.A(n_3972),
.Y(n_4181)
);

HB1xp67_ASAP7_75t_L g4182 ( 
.A(n_3943),
.Y(n_4182)
);

OR2x6_ASAP7_75t_L g4183 ( 
.A(n_4072),
.B(n_4084),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_3971),
.Y(n_4184)
);

O2A1O1Ixp33_ASAP7_75t_SL g4185 ( 
.A1(n_4005),
.A2(n_3696),
.B(n_3735),
.C(n_3825),
.Y(n_4185)
);

NAND2xp33_ASAP7_75t_R g4186 ( 
.A(n_4072),
.B(n_3869),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3909),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4052),
.Y(n_4188)
);

NAND2xp33_ASAP7_75t_R g4189 ( 
.A(n_4039),
.B(n_3869),
.Y(n_4189)
);

NAND2xp33_ASAP7_75t_R g4190 ( 
.A(n_3913),
.B(n_3882),
.Y(n_4190)
);

AND2x4_ASAP7_75t_L g4191 ( 
.A(n_4105),
.B(n_4075),
.Y(n_4191)
);

INVx1_ASAP7_75t_SL g4192 ( 
.A(n_4126),
.Y(n_4192)
);

INVx2_ASAP7_75t_L g4193 ( 
.A(n_4122),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4095),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_4168),
.B(n_4053),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_4124),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4182),
.B(n_4064),
.Y(n_4197)
);

AND2x2_ASAP7_75t_L g4198 ( 
.A(n_4094),
.B(n_3949),
.Y(n_4198)
);

HB1xp67_ASAP7_75t_L g4199 ( 
.A(n_4117),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4104),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_4187),
.B(n_4089),
.Y(n_4201)
);

OR2x2_ASAP7_75t_L g4202 ( 
.A(n_4149),
.B(n_3977),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_4129),
.Y(n_4203)
);

NAND3xp33_ASAP7_75t_L g4204 ( 
.A(n_4111),
.B(n_3989),
.C(n_4050),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4114),
.Y(n_4205)
);

BUFx3_ASAP7_75t_L g4206 ( 
.A(n_4156),
.Y(n_4206)
);

NOR2xp33_ASAP7_75t_L g4207 ( 
.A(n_4102),
.B(n_4056),
.Y(n_4207)
);

INVx2_ASAP7_75t_L g4208 ( 
.A(n_4143),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_4145),
.B(n_4000),
.Y(n_4209)
);

INVx2_ASAP7_75t_L g4210 ( 
.A(n_4176),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_4184),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_4188),
.Y(n_4212)
);

HB1xp67_ASAP7_75t_L g4213 ( 
.A(n_4173),
.Y(n_4213)
);

HB1xp67_ASAP7_75t_L g4214 ( 
.A(n_4175),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4115),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_4152),
.B(n_4065),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_4120),
.B(n_4028),
.Y(n_4217)
);

HB1xp67_ASAP7_75t_L g4218 ( 
.A(n_4151),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_4127),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_4133),
.B(n_4048),
.Y(n_4220)
);

AND2x2_ASAP7_75t_L g4221 ( 
.A(n_4140),
.B(n_4051),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_4166),
.B(n_4141),
.Y(n_4222)
);

AND2x2_ASAP7_75t_L g4223 ( 
.A(n_4153),
.B(n_4164),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_4169),
.Y(n_4224)
);

AOI221xp5_ASAP7_75t_L g4225 ( 
.A1(n_4134),
.A2(n_4043),
.B1(n_3920),
.B2(n_4076),
.C(n_4074),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_4172),
.B(n_4069),
.Y(n_4226)
);

INVx3_ASAP7_75t_L g4227 ( 
.A(n_4155),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4177),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4178),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4180),
.Y(n_4230)
);

HB1xp67_ASAP7_75t_L g4231 ( 
.A(n_4158),
.Y(n_4231)
);

INVx3_ASAP7_75t_L g4232 ( 
.A(n_4155),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_4161),
.Y(n_4233)
);

HB1xp67_ASAP7_75t_L g4234 ( 
.A(n_4107),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_4163),
.B(n_4077),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4147),
.Y(n_4236)
);

AND2x4_ASAP7_75t_L g4237 ( 
.A(n_4101),
.B(n_3740),
.Y(n_4237)
);

OA21x2_ASAP7_75t_L g4238 ( 
.A1(n_4142),
.A2(n_3902),
.B(n_4087),
.Y(n_4238)
);

INVx4_ASAP7_75t_L g4239 ( 
.A(n_4098),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_SL g4240 ( 
.A(n_4099),
.B(n_3960),
.Y(n_4240)
);

AND2x2_ASAP7_75t_L g4241 ( 
.A(n_4146),
.B(n_3922),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_4106),
.B(n_3664),
.Y(n_4242)
);

BUFx3_ASAP7_75t_L g4243 ( 
.A(n_4156),
.Y(n_4243)
);

HB1xp67_ASAP7_75t_L g4244 ( 
.A(n_4160),
.Y(n_4244)
);

AND2x4_ASAP7_75t_L g4245 ( 
.A(n_4136),
.B(n_4100),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_4123),
.B(n_3664),
.Y(n_4246)
);

AND2x2_ASAP7_75t_L g4247 ( 
.A(n_4136),
.B(n_3988),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4157),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4139),
.Y(n_4249)
);

AND2x2_ASAP7_75t_L g4250 ( 
.A(n_4096),
.B(n_3988),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_4097),
.B(n_3925),
.Y(n_4251)
);

AO21x2_ASAP7_75t_L g4252 ( 
.A1(n_4110),
.A2(n_4002),
.B(n_4003),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4097),
.B(n_3986),
.Y(n_4253)
);

AND2x4_ASAP7_75t_L g4254 ( 
.A(n_4113),
.B(n_4183),
.Y(n_4254)
);

AND2x2_ASAP7_75t_L g4255 ( 
.A(n_4097),
.B(n_3996),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4137),
.Y(n_4256)
);

AOI221xp5_ASAP7_75t_L g4257 ( 
.A1(n_4121),
.A2(n_4007),
.B1(n_4020),
.B2(n_3923),
.C(n_4083),
.Y(n_4257)
);

INVx2_ASAP7_75t_SL g4258 ( 
.A(n_4159),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_4157),
.Y(n_4259)
);

HB1xp67_ASAP7_75t_L g4260 ( 
.A(n_4183),
.Y(n_4260)
);

INVx2_ASAP7_75t_L g4261 ( 
.A(n_4157),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_4109),
.B(n_3973),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4113),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_4162),
.Y(n_4264)
);

OAI22xp5_ASAP7_75t_L g4265 ( 
.A1(n_4240),
.A2(n_4108),
.B1(n_4135),
.B2(n_4165),
.Y(n_4265)
);

AND2x2_ASAP7_75t_L g4266 ( 
.A(n_4231),
.B(n_4119),
.Y(n_4266)
);

NOR2xp33_ASAP7_75t_L g4267 ( 
.A(n_4239),
.B(n_4116),
.Y(n_4267)
);

OAI21xp33_ASAP7_75t_L g4268 ( 
.A1(n_4256),
.A2(n_4174),
.B(n_4112),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4195),
.B(n_4150),
.Y(n_4269)
);

AND2x2_ASAP7_75t_L g4270 ( 
.A(n_4250),
.B(n_4179),
.Y(n_4270)
);

OAI21xp5_ASAP7_75t_SL g4271 ( 
.A1(n_4254),
.A2(n_4125),
.B(n_4118),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_4195),
.B(n_4092),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_4197),
.B(n_3728),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4250),
.B(n_4179),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_4234),
.B(n_4171),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_4197),
.B(n_4023),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_L g4277 ( 
.A(n_4199),
.B(n_4026),
.Y(n_4277)
);

OA21x2_ASAP7_75t_L g4278 ( 
.A1(n_4256),
.A2(n_4128),
.B(n_3935),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4214),
.B(n_4026),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_L g4280 ( 
.A(n_4198),
.B(n_4132),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4198),
.B(n_4067),
.Y(n_4281)
);

OAI22xp5_ASAP7_75t_L g4282 ( 
.A1(n_4260),
.A2(n_4171),
.B1(n_4154),
.B2(n_3962),
.Y(n_4282)
);

OAI21xp5_ASAP7_75t_L g4283 ( 
.A1(n_4204),
.A2(n_4004),
.B(n_3985),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4223),
.B(n_4216),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_4223),
.B(n_4079),
.Y(n_4285)
);

NAND3xp33_ASAP7_75t_L g4286 ( 
.A(n_4249),
.B(n_4138),
.C(n_4189),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_4217),
.B(n_4071),
.Y(n_4287)
);

OA21x2_ASAP7_75t_L g4288 ( 
.A1(n_4249),
.A2(n_3983),
.B(n_3967),
.Y(n_4288)
);

NAND3xp33_ASAP7_75t_L g4289 ( 
.A(n_4257),
.B(n_4238),
.C(n_4225),
.Y(n_4289)
);

AND2x2_ASAP7_75t_L g4290 ( 
.A(n_4191),
.B(n_4170),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_4217),
.B(n_4085),
.Y(n_4291)
);

AND2x2_ASAP7_75t_L g4292 ( 
.A(n_4191),
.B(n_4181),
.Y(n_4292)
);

AND2x2_ASAP7_75t_SL g4293 ( 
.A(n_4245),
.B(n_4254),
.Y(n_4293)
);

AND2x2_ASAP7_75t_L g4294 ( 
.A(n_4191),
.B(n_3936),
.Y(n_4294)
);

AOI22xp33_ASAP7_75t_L g4295 ( 
.A1(n_4262),
.A2(n_3964),
.B1(n_4014),
.B2(n_3914),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_4220),
.B(n_4221),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_4241),
.B(n_4059),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4220),
.B(n_4221),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4226),
.B(n_4019),
.Y(n_4299)
);

NAND3xp33_ASAP7_75t_L g4300 ( 
.A(n_4239),
.B(n_4244),
.C(n_4218),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_4226),
.B(n_4037),
.Y(n_4301)
);

NAND3xp33_ASAP7_75t_L g4302 ( 
.A(n_4238),
.B(n_4186),
.C(n_4130),
.Y(n_4302)
);

OAI21xp5_ASAP7_75t_SL g4303 ( 
.A1(n_4254),
.A2(n_4011),
.B(n_3942),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_4246),
.B(n_3966),
.Y(n_4304)
);

NOR2xp33_ASAP7_75t_L g4305 ( 
.A(n_4239),
.B(n_4103),
.Y(n_4305)
);

AND2x2_ASAP7_75t_L g4306 ( 
.A(n_4241),
.B(n_3968),
.Y(n_4306)
);

AND2x2_ASAP7_75t_L g4307 ( 
.A(n_4263),
.B(n_3990),
.Y(n_4307)
);

NAND4xp25_ASAP7_75t_L g4308 ( 
.A(n_4207),
.B(n_3955),
.C(n_4190),
.D(n_3995),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_4246),
.B(n_4009),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_4242),
.B(n_3978),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4242),
.B(n_3982),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_4202),
.B(n_4081),
.Y(n_4312)
);

AND2x2_ASAP7_75t_L g4313 ( 
.A(n_4247),
.B(n_3990),
.Y(n_4313)
);

OAI22xp5_ASAP7_75t_L g4314 ( 
.A1(n_4258),
.A2(n_4022),
.B1(n_4047),
.B2(n_4027),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_SL g4315 ( 
.A(n_4245),
.B(n_4148),
.Y(n_4315)
);

NOR2xp33_ASAP7_75t_L g4316 ( 
.A(n_4192),
.B(n_4131),
.Y(n_4316)
);

AND2x2_ASAP7_75t_L g4317 ( 
.A(n_4247),
.B(n_3993),
.Y(n_4317)
);

OA21x2_ASAP7_75t_L g4318 ( 
.A1(n_4264),
.A2(n_4237),
.B(n_4251),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_4202),
.B(n_4057),
.Y(n_4319)
);

OAI221xp5_ASAP7_75t_L g4320 ( 
.A1(n_4264),
.A2(n_4035),
.B1(n_4062),
.B2(n_4040),
.C(n_3950),
.Y(n_4320)
);

OAI22xp5_ASAP7_75t_L g4321 ( 
.A1(n_4258),
.A2(n_3953),
.B1(n_4088),
.B2(n_4091),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4235),
.B(n_4070),
.Y(n_4322)
);

NAND3xp33_ASAP7_75t_L g4323 ( 
.A(n_4238),
.B(n_4010),
.C(n_4017),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_4235),
.B(n_4185),
.Y(n_4324)
);

INVx3_ASAP7_75t_L g4325 ( 
.A(n_4245),
.Y(n_4325)
);

OAI221xp5_ASAP7_75t_SL g4326 ( 
.A1(n_4262),
.A2(n_3992),
.B1(n_4068),
.B2(n_4060),
.C(n_4066),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4233),
.B(n_3993),
.Y(n_4327)
);

AOI22xp33_ASAP7_75t_SL g4328 ( 
.A1(n_4206),
.A2(n_4049),
.B1(n_4144),
.B2(n_3997),
.Y(n_4328)
);

AOI221xp5_ASAP7_75t_L g4329 ( 
.A1(n_4201),
.A2(n_4030),
.B1(n_4024),
.B2(n_4078),
.C(n_4038),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4236),
.B(n_4093),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_SL g4331 ( 
.A(n_4227),
.B(n_3998),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_4325),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4296),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4298),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4325),
.Y(n_4335)
);

O2A1O1Ixp33_ASAP7_75t_L g4336 ( 
.A1(n_4289),
.A2(n_4206),
.B(n_4243),
.C(n_4213),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4293),
.B(n_4227),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4284),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4300),
.Y(n_4339)
);

AND2x2_ASAP7_75t_L g4340 ( 
.A(n_4270),
.B(n_4227),
.Y(n_4340)
);

INVx2_ASAP7_75t_L g4341 ( 
.A(n_4318),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4300),
.Y(n_4342)
);

AND2x2_ASAP7_75t_L g4343 ( 
.A(n_4274),
.B(n_4232),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_4273),
.B(n_4219),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4272),
.Y(n_4345)
);

AND2x4_ASAP7_75t_SL g4346 ( 
.A(n_4290),
.B(n_4232),
.Y(n_4346)
);

AND2x4_ASAP7_75t_SL g4347 ( 
.A(n_4292),
.B(n_4232),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_4277),
.B(n_4219),
.Y(n_4348)
);

OR2x2_ASAP7_75t_L g4349 ( 
.A(n_4269),
.B(n_4222),
.Y(n_4349)
);

INVx2_ASAP7_75t_L g4350 ( 
.A(n_4318),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4279),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4313),
.B(n_4251),
.Y(n_4352)
);

INVx2_ASAP7_75t_L g4353 ( 
.A(n_4266),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4312),
.B(n_4224),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4317),
.B(n_4237),
.Y(n_4355)
);

AND2x2_ASAP7_75t_L g4356 ( 
.A(n_4294),
.B(n_4237),
.Y(n_4356)
);

NAND2x1_ASAP7_75t_L g4357 ( 
.A(n_4286),
.B(n_4253),
.Y(n_4357)
);

AND2x2_ASAP7_75t_L g4358 ( 
.A(n_4306),
.B(n_4253),
.Y(n_4358)
);

OAI221xp5_ASAP7_75t_SL g4359 ( 
.A1(n_4303),
.A2(n_4243),
.B1(n_4255),
.B2(n_4058),
.C(n_4229),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_SL g4360 ( 
.A(n_4265),
.B(n_4255),
.Y(n_4360)
);

OR2x2_ASAP7_75t_L g4361 ( 
.A(n_4311),
.B(n_4193),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4287),
.Y(n_4362)
);

AND2x4_ASAP7_75t_SL g4363 ( 
.A(n_4275),
.B(n_4209),
.Y(n_4363)
);

OR2x2_ASAP7_75t_L g4364 ( 
.A(n_4304),
.B(n_4193),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4324),
.Y(n_4365)
);

OR2x2_ASAP7_75t_L g4366 ( 
.A(n_4310),
.B(n_4196),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4276),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4299),
.Y(n_4368)
);

HB1xp67_ASAP7_75t_L g4369 ( 
.A(n_4315),
.Y(n_4369)
);

AND2x2_ASAP7_75t_L g4370 ( 
.A(n_4297),
.B(n_4209),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4301),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4319),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4268),
.B(n_4224),
.Y(n_4373)
);

INVx3_ASAP7_75t_L g4374 ( 
.A(n_4288),
.Y(n_4374)
);

AND2x2_ASAP7_75t_L g4375 ( 
.A(n_4280),
.B(n_4248),
.Y(n_4375)
);

HB1xp67_ASAP7_75t_L g4376 ( 
.A(n_4339),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4333),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4341),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4334),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4338),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4362),
.Y(n_4381)
);

AND2x2_ASAP7_75t_L g4382 ( 
.A(n_4369),
.B(n_4271),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_4350),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4364),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_4372),
.B(n_4268),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_L g4386 ( 
.A(n_4345),
.B(n_4205),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_4351),
.B(n_4205),
.Y(n_4387)
);

INVx2_ASAP7_75t_L g4388 ( 
.A(n_4366),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4368),
.Y(n_4389)
);

AND2x2_ASAP7_75t_L g4390 ( 
.A(n_4369),
.B(n_4282),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4371),
.Y(n_4391)
);

AND2x2_ASAP7_75t_L g4392 ( 
.A(n_4337),
.B(n_4346),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4346),
.B(n_4278),
.Y(n_4393)
);

INVx2_ASAP7_75t_SL g4394 ( 
.A(n_4347),
.Y(n_4394)
);

AND2x2_ASAP7_75t_L g4395 ( 
.A(n_4347),
.B(n_4278),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4356),
.B(n_4307),
.Y(n_4396)
);

AND2x2_ASAP7_75t_L g4397 ( 
.A(n_4355),
.B(n_4330),
.Y(n_4397)
);

INVxp67_ASAP7_75t_L g4398 ( 
.A(n_4342),
.Y(n_4398)
);

INVx2_ASAP7_75t_SL g4399 ( 
.A(n_4363),
.Y(n_4399)
);

AND2x2_ASAP7_75t_L g4400 ( 
.A(n_4340),
.B(n_4267),
.Y(n_4400)
);

OR2x2_ASAP7_75t_L g4401 ( 
.A(n_4344),
.B(n_4309),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4343),
.B(n_4285),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_4365),
.B(n_4215),
.Y(n_4403)
);

OR2x2_ASAP7_75t_L g4404 ( 
.A(n_4344),
.B(n_4322),
.Y(n_4404)
);

OR2x2_ASAP7_75t_L g4405 ( 
.A(n_4354),
.B(n_4281),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4367),
.Y(n_4406)
);

INVx4_ASAP7_75t_L g4407 ( 
.A(n_4363),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4361),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_4348),
.B(n_4215),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_4375),
.B(n_4288),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_4332),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4348),
.Y(n_4412)
);

INVx3_ASAP7_75t_L g4413 ( 
.A(n_4357),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4358),
.B(n_4302),
.Y(n_4414)
);

AND2x2_ASAP7_75t_L g4415 ( 
.A(n_4352),
.B(n_4291),
.Y(n_4415)
);

OR2x2_ASAP7_75t_L g4416 ( 
.A(n_4354),
.B(n_4212),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_4349),
.B(n_4228),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4403),
.Y(n_4418)
);

NOR2x1p5_ASAP7_75t_L g4419 ( 
.A(n_4407),
.B(n_4373),
.Y(n_4419)
);

NOR2xp67_ASAP7_75t_L g4420 ( 
.A(n_4413),
.B(n_4374),
.Y(n_4420)
);

OR2x6_ASAP7_75t_L g4421 ( 
.A(n_4407),
.B(n_4336),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4390),
.B(n_4336),
.Y(n_4422)
);

INVx1_ASAP7_75t_SL g4423 ( 
.A(n_4376),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4403),
.Y(n_4424)
);

AND2x2_ASAP7_75t_L g4425 ( 
.A(n_4392),
.B(n_4335),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_4386),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_4385),
.B(n_4360),
.Y(n_4427)
);

OAI211xp5_ASAP7_75t_L g4428 ( 
.A1(n_4398),
.A2(n_4283),
.B(n_4360),
.C(n_4359),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4386),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_4417),
.Y(n_4430)
);

AND2x2_ASAP7_75t_L g4431 ( 
.A(n_4394),
.B(n_4332),
.Y(n_4431)
);

AOI32xp33_ASAP7_75t_L g4432 ( 
.A1(n_4382),
.A2(n_4374),
.A3(n_4328),
.B1(n_4373),
.B2(n_4295),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4417),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4384),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_4385),
.B(n_4398),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4408),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4387),
.Y(n_4437)
);

HB1xp67_ASAP7_75t_L g4438 ( 
.A(n_4376),
.Y(n_4438)
);

AND2x2_ASAP7_75t_L g4439 ( 
.A(n_4394),
.B(n_4370),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4387),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_4381),
.B(n_4406),
.Y(n_4441)
);

AND2x2_ASAP7_75t_L g4442 ( 
.A(n_4399),
.B(n_4353),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4378),
.Y(n_4443)
);

OR2x2_ASAP7_75t_L g4444 ( 
.A(n_4404),
.B(n_4359),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4405),
.Y(n_4445)
);

HB1xp67_ASAP7_75t_L g4446 ( 
.A(n_4378),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4427),
.B(n_4380),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4438),
.Y(n_4448)
);

OR2x2_ASAP7_75t_L g4449 ( 
.A(n_4445),
.B(n_4401),
.Y(n_4449)
);

OR2x2_ASAP7_75t_L g4450 ( 
.A(n_4435),
.B(n_4388),
.Y(n_4450)
);

AND2x2_ASAP7_75t_L g4451 ( 
.A(n_4421),
.B(n_4399),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4423),
.B(n_4377),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_4423),
.B(n_4442),
.Y(n_4453)
);

NAND3xp33_ASAP7_75t_L g4454 ( 
.A(n_4432),
.B(n_4413),
.C(n_4383),
.Y(n_4454)
);

AND2x2_ASAP7_75t_L g4455 ( 
.A(n_4421),
.B(n_4400),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_4421),
.B(n_4393),
.Y(n_4456)
);

NOR2xp33_ASAP7_75t_L g4457 ( 
.A(n_4422),
.B(n_4305),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4439),
.B(n_4395),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4446),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_4444),
.B(n_4389),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4431),
.Y(n_4461)
);

INVx2_ASAP7_75t_L g4462 ( 
.A(n_4443),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4441),
.Y(n_4463)
);

INVxp67_ASAP7_75t_SL g4464 ( 
.A(n_4419),
.Y(n_4464)
);

AND2x4_ASAP7_75t_SL g4465 ( 
.A(n_4425),
.B(n_4316),
.Y(n_4465)
);

OR2x2_ASAP7_75t_L g4466 ( 
.A(n_4434),
.B(n_4388),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4418),
.B(n_4379),
.Y(n_4467)
);

NOR2xp33_ASAP7_75t_L g4468 ( 
.A(n_4428),
.B(n_4391),
.Y(n_4468)
);

INVx2_ASAP7_75t_L g4469 ( 
.A(n_4436),
.Y(n_4469)
);

AND2x4_ASAP7_75t_L g4470 ( 
.A(n_4451),
.B(n_4465),
.Y(n_4470)
);

INVx2_ASAP7_75t_L g4471 ( 
.A(n_4459),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4450),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4453),
.Y(n_4473)
);

AND2x2_ASAP7_75t_L g4474 ( 
.A(n_4458),
.B(n_4414),
.Y(n_4474)
);

AND2x2_ASAP7_75t_L g4475 ( 
.A(n_4456),
.B(n_4430),
.Y(n_4475)
);

AOI21xp5_ASAP7_75t_L g4476 ( 
.A1(n_4464),
.A2(n_4420),
.B(n_4383),
.Y(n_4476)
);

AOI22xp5_ASAP7_75t_L g4477 ( 
.A1(n_4457),
.A2(n_4433),
.B1(n_4420),
.B2(n_4440),
.Y(n_4477)
);

AOI22xp33_ASAP7_75t_L g4478 ( 
.A1(n_4455),
.A2(n_4426),
.B1(n_4429),
.B2(n_4424),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4452),
.Y(n_4479)
);

AOI21xp33_ASAP7_75t_SL g4480 ( 
.A1(n_4454),
.A2(n_4437),
.B(n_4167),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_L g4481 ( 
.A(n_4468),
.B(n_4412),
.Y(n_4481)
);

AOI21xp5_ASAP7_75t_L g4482 ( 
.A1(n_4454),
.A2(n_4411),
.B(n_4314),
.Y(n_4482)
);

NOR2xp33_ASAP7_75t_L g4483 ( 
.A(n_4461),
.B(n_4410),
.Y(n_4483)
);

AOI21xp33_ASAP7_75t_L g4484 ( 
.A1(n_4448),
.A2(n_4323),
.B(n_4411),
.Y(n_4484)
);

NOR2x1_ASAP7_75t_L g4485 ( 
.A(n_4460),
.B(n_4308),
.Y(n_4485)
);

AOI22xp5_ASAP7_75t_L g4486 ( 
.A1(n_4463),
.A2(n_4321),
.B1(n_4323),
.B2(n_4252),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_4462),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4449),
.B(n_4415),
.Y(n_4488)
);

AND2x4_ASAP7_75t_L g4489 ( 
.A(n_4469),
.B(n_4466),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4447),
.B(n_4402),
.Y(n_4490)
);

AOI211x1_ASAP7_75t_L g4491 ( 
.A1(n_4452),
.A2(n_4409),
.B(n_4320),
.C(n_4331),
.Y(n_4491)
);

OAI22xp33_ASAP7_75t_L g4492 ( 
.A1(n_4467),
.A2(n_4409),
.B1(n_4416),
.B2(n_4327),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4467),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_4468),
.B(n_4252),
.Y(n_4494)
);

AOI22xp5_ASAP7_75t_L g4495 ( 
.A1(n_4457),
.A2(n_4252),
.B1(n_4397),
.B2(n_4396),
.Y(n_4495)
);

INVx1_ASAP7_75t_SL g4496 ( 
.A(n_4470),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_4470),
.B(n_4194),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_4488),
.B(n_4200),
.Y(n_4498)
);

OAI211xp5_ASAP7_75t_SL g4499 ( 
.A1(n_4473),
.A2(n_4329),
.B(n_4063),
.C(n_3999),
.Y(n_4499)
);

INVx1_ASAP7_75t_SL g4500 ( 
.A(n_4487),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4472),
.Y(n_4501)
);

NOR2x1_ASAP7_75t_L g4502 ( 
.A(n_4471),
.B(n_4061),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4489),
.Y(n_4503)
);

INVx2_ASAP7_75t_L g4504 ( 
.A(n_4489),
.Y(n_4504)
);

AND2x4_ASAP7_75t_L g4505 ( 
.A(n_4475),
.B(n_4230),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4479),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4483),
.Y(n_4507)
);

INVx2_ASAP7_75t_L g4508 ( 
.A(n_4474),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4490),
.B(n_4228),
.Y(n_4509)
);

OAI22xp5_ASAP7_75t_L g4510 ( 
.A1(n_4486),
.A2(n_4326),
.B1(n_4001),
.B2(n_4259),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4493),
.Y(n_4511)
);

AOI22xp5_ASAP7_75t_L g4512 ( 
.A1(n_4485),
.A2(n_4248),
.B1(n_4261),
.B2(n_4259),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4481),
.Y(n_4513)
);

AND2x2_ASAP7_75t_L g4514 ( 
.A(n_4482),
.B(n_4477),
.Y(n_4514)
);

OAI21xp5_ASAP7_75t_L g4515 ( 
.A1(n_4476),
.A2(n_3705),
.B(n_3734),
.Y(n_4515)
);

NOR2xp33_ASAP7_75t_L g4516 ( 
.A(n_4480),
.B(n_4484),
.Y(n_4516)
);

A2O1A1Ixp33_ASAP7_75t_L g4517 ( 
.A1(n_4494),
.A2(n_4261),
.B(n_3987),
.C(n_4212),
.Y(n_4517)
);

INVx1_ASAP7_75t_SL g4518 ( 
.A(n_4495),
.Y(n_4518)
);

OAI21xp5_ASAP7_75t_L g4519 ( 
.A1(n_4478),
.A2(n_3723),
.B(n_3673),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4491),
.B(n_4196),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4492),
.Y(n_4521)
);

OAI22xp5_ASAP7_75t_L g4522 ( 
.A1(n_4486),
.A2(n_4203),
.B1(n_4210),
.B2(n_4208),
.Y(n_4522)
);

OAI21xp33_ASAP7_75t_SL g4523 ( 
.A1(n_4496),
.A2(n_3980),
.B(n_4203),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_SL g4524 ( 
.A(n_4514),
.B(n_3998),
.Y(n_4524)
);

OR2x2_ASAP7_75t_L g4525 ( 
.A(n_4500),
.B(n_4208),
.Y(n_4525)
);

AOI221x1_ASAP7_75t_L g4526 ( 
.A1(n_4506),
.A2(n_472),
.B1(n_470),
.B2(n_471),
.C(n_473),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4508),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_4503),
.Y(n_4528)
);

OAI221xp5_ASAP7_75t_L g4529 ( 
.A1(n_4510),
.A2(n_3998),
.B1(n_3723),
.B2(n_3882),
.C(n_3653),
.Y(n_4529)
);

NOR3xp33_ASAP7_75t_L g4530 ( 
.A(n_4516),
.B(n_3817),
.C(n_3840),
.Y(n_4530)
);

OAI21xp33_ASAP7_75t_SL g4531 ( 
.A1(n_4521),
.A2(n_4211),
.B(n_4210),
.Y(n_4531)
);

AOI22xp5_ASAP7_75t_L g4532 ( 
.A1(n_4507),
.A2(n_4504),
.B1(n_4513),
.B2(n_4518),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_4497),
.B(n_4211),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_SL g4534 ( 
.A(n_4501),
.B(n_3653),
.Y(n_4534)
);

AOI22xp5_ASAP7_75t_L g4535 ( 
.A1(n_4499),
.A2(n_3713),
.B1(n_3704),
.B2(n_3737),
.Y(n_4535)
);

OAI221xp5_ASAP7_75t_L g4536 ( 
.A1(n_4502),
.A2(n_3817),
.B1(n_3624),
.B2(n_474),
.C(n_471),
.Y(n_4536)
);

AOI22xp5_ASAP7_75t_L g4537 ( 
.A1(n_4520),
.A2(n_3713),
.B1(n_3704),
.B2(n_3650),
.Y(n_4537)
);

OAI31xp33_ASAP7_75t_L g4538 ( 
.A1(n_4511),
.A2(n_475),
.A3(n_472),
.B(n_474),
.Y(n_4538)
);

AOI221xp5_ASAP7_75t_L g4539 ( 
.A1(n_4522),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.C(n_478),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_SL g4540 ( 
.A(n_4512),
.B(n_3624),
.Y(n_4540)
);

OAI22xp33_ASAP7_75t_L g4541 ( 
.A1(n_4498),
.A2(n_479),
.B1(n_476),
.B2(n_478),
.Y(n_4541)
);

AOI22xp5_ASAP7_75t_L g4542 ( 
.A1(n_4502),
.A2(n_3656),
.B1(n_3663),
.B2(n_3846),
.Y(n_4542)
);

OAI21xp5_ASAP7_75t_L g4543 ( 
.A1(n_4515),
.A2(n_3851),
.B(n_3790),
.Y(n_4543)
);

AOI22xp5_ASAP7_75t_L g4544 ( 
.A1(n_4505),
.A2(n_3781),
.B1(n_3822),
.B2(n_3820),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_L g4545 ( 
.A(n_4505),
.B(n_479),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_4509),
.Y(n_4546)
);

AOI322xp5_ASAP7_75t_L g4547 ( 
.A1(n_4517),
.A2(n_480),
.A3(n_481),
.B1(n_482),
.B2(n_483),
.C1(n_484),
.C2(n_485),
.Y(n_4547)
);

AO22x1_ASAP7_75t_L g4548 ( 
.A1(n_4519),
.A2(n_484),
.B1(n_480),
.B2(n_481),
.Y(n_4548)
);

XOR2x2_ASAP7_75t_L g4549 ( 
.A(n_4496),
.B(n_486),
.Y(n_4549)
);

INVxp67_ASAP7_75t_L g4550 ( 
.A(n_4496),
.Y(n_4550)
);

AOI21xp5_ASAP7_75t_L g4551 ( 
.A1(n_4496),
.A2(n_3799),
.B(n_3798),
.Y(n_4551)
);

OAI322xp33_ASAP7_75t_SL g4552 ( 
.A1(n_4513),
.A2(n_487),
.A3(n_488),
.B1(n_489),
.B2(n_490),
.C1(n_491),
.C2(n_492),
.Y(n_4552)
);

NOR2xp33_ASAP7_75t_L g4553 ( 
.A(n_4496),
.B(n_487),
.Y(n_4553)
);

NOR3x1_ASAP7_75t_L g4554 ( 
.A(n_4524),
.B(n_3808),
.C(n_3766),
.Y(n_4554)
);

NAND3xp33_ASAP7_75t_L g4555 ( 
.A(n_4550),
.B(n_489),
.C(n_492),
.Y(n_4555)
);

HB1xp67_ASAP7_75t_L g4556 ( 
.A(n_4528),
.Y(n_4556)
);

AOI22xp5_ASAP7_75t_L g4557 ( 
.A1(n_4553),
.A2(n_3626),
.B1(n_3727),
.B2(n_3738),
.Y(n_4557)
);

NOR3xp33_ASAP7_75t_L g4558 ( 
.A(n_4541),
.B(n_493),
.C(n_494),
.Y(n_4558)
);

AOI211x1_ASAP7_75t_L g4559 ( 
.A1(n_4527),
.A2(n_499),
.B(n_493),
.C(n_498),
.Y(n_4559)
);

AOI22xp5_ASAP7_75t_L g4560 ( 
.A1(n_4549),
.A2(n_3889),
.B1(n_3712),
.B2(n_3646),
.Y(n_4560)
);

AOI21xp5_ASAP7_75t_L g4561 ( 
.A1(n_4545),
.A2(n_3833),
.B(n_3795),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4525),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4532),
.Y(n_4563)
);

OAI21xp5_ASAP7_75t_L g4564 ( 
.A1(n_4531),
.A2(n_3792),
.B(n_3641),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_SL g4565 ( 
.A(n_4538),
.B(n_3761),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4548),
.B(n_4547),
.Y(n_4566)
);

NOR3x1_ASAP7_75t_L g4567 ( 
.A(n_4536),
.B(n_498),
.C(n_499),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4546),
.Y(n_4568)
);

NOR3xp33_ASAP7_75t_SL g4569 ( 
.A(n_4539),
.B(n_4523),
.C(n_4529),
.Y(n_4569)
);

AOI211xp5_ASAP7_75t_L g4570 ( 
.A1(n_4551),
.A2(n_502),
.B(n_500),
.C(n_501),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4526),
.Y(n_4571)
);

OAI22xp33_ASAP7_75t_L g4572 ( 
.A1(n_4537),
.A2(n_504),
.B1(n_500),
.B2(n_503),
.Y(n_4572)
);

NOR3xp33_ASAP7_75t_SL g4573 ( 
.A(n_4534),
.B(n_505),
.C(n_506),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_SL g4574 ( 
.A(n_4540),
.B(n_3717),
.Y(n_4574)
);

INVx3_ASAP7_75t_L g4575 ( 
.A(n_4533),
.Y(n_4575)
);

AOI21xp5_ASAP7_75t_L g4576 ( 
.A1(n_4552),
.A2(n_505),
.B(n_506),
.Y(n_4576)
);

XNOR2x1_ASAP7_75t_SL g4577 ( 
.A(n_4535),
.B(n_4530),
.Y(n_4577)
);

NOR4xp25_ASAP7_75t_L g4578 ( 
.A(n_4543),
.B(n_510),
.C(n_507),
.D(n_508),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_4542),
.B(n_507),
.Y(n_4579)
);

NOR2x1_ASAP7_75t_L g4580 ( 
.A(n_4544),
.B(n_510),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4556),
.Y(n_4581)
);

NAND4xp25_ASAP7_75t_L g4582 ( 
.A(n_4576),
.B(n_513),
.C(n_511),
.D(n_512),
.Y(n_4582)
);

OR3x1_ASAP7_75t_L g4583 ( 
.A(n_4563),
.B(n_511),
.C(n_512),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4571),
.Y(n_4584)
);

NAND3xp33_ASAP7_75t_L g4585 ( 
.A(n_4555),
.B(n_513),
.C(n_515),
.Y(n_4585)
);

O2A1O1Ixp5_ASAP7_75t_SL g4586 ( 
.A1(n_4568),
.A2(n_518),
.B(n_516),
.C(n_517),
.Y(n_4586)
);

AOI221xp5_ASAP7_75t_L g4587 ( 
.A1(n_4578),
.A2(n_516),
.B1(n_518),
.B2(n_519),
.C(n_520),
.Y(n_4587)
);

O2A1O1Ixp33_ASAP7_75t_L g4588 ( 
.A1(n_4558),
.A2(n_522),
.B(n_519),
.C(n_521),
.Y(n_4588)
);

NAND3xp33_ASAP7_75t_SL g4589 ( 
.A(n_4570),
.B(n_4566),
.C(n_4579),
.Y(n_4589)
);

NAND4xp75_ASAP7_75t_L g4590 ( 
.A(n_4567),
.B(n_523),
.C(n_521),
.D(n_522),
.Y(n_4590)
);

NOR2xp33_ASAP7_75t_L g4591 ( 
.A(n_4562),
.B(n_524),
.Y(n_4591)
);

BUFx6f_ASAP7_75t_L g4592 ( 
.A(n_4565),
.Y(n_4592)
);

NAND3xp33_ASAP7_75t_L g4593 ( 
.A(n_4559),
.B(n_524),
.C(n_525),
.Y(n_4593)
);

AOI21x1_ASAP7_75t_L g4594 ( 
.A1(n_4580),
.A2(n_525),
.B(n_526),
.Y(n_4594)
);

NAND4xp25_ASAP7_75t_SL g4595 ( 
.A(n_4560),
.B(n_531),
.C(n_527),
.D(n_530),
.Y(n_4595)
);

INVx2_ASAP7_75t_L g4596 ( 
.A(n_4554),
.Y(n_4596)
);

NAND2xp5_ASAP7_75t_SL g4597 ( 
.A(n_4572),
.B(n_527),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4575),
.Y(n_4598)
);

NAND3xp33_ASAP7_75t_L g4599 ( 
.A(n_4573),
.B(n_531),
.C(n_532),
.Y(n_4599)
);

NOR3xp33_ASAP7_75t_L g4600 ( 
.A(n_4575),
.B(n_533),
.C(n_534),
.Y(n_4600)
);

OAI22xp33_ASAP7_75t_L g4601 ( 
.A1(n_4557),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_4601)
);

A2O1A1Ixp33_ASAP7_75t_L g4602 ( 
.A1(n_4569),
.A2(n_3754),
.B(n_3753),
.C(n_3744),
.Y(n_4602)
);

NOR2xp33_ASAP7_75t_L g4603 ( 
.A(n_4574),
.B(n_537),
.Y(n_4603)
);

NAND3xp33_ASAP7_75t_SL g4604 ( 
.A(n_4561),
.B(n_538),
.C(n_539),
.Y(n_4604)
);

NOR2xp33_ASAP7_75t_L g4605 ( 
.A(n_4577),
.B(n_538),
.Y(n_4605)
);

NOR3xp33_ASAP7_75t_L g4606 ( 
.A(n_4564),
.B(n_540),
.C(n_541),
.Y(n_4606)
);

NOR3xp33_ASAP7_75t_L g4607 ( 
.A(n_4584),
.B(n_540),
.C(n_541),
.Y(n_4607)
);

NOR2x1_ASAP7_75t_L g4608 ( 
.A(n_4583),
.B(n_542),
.Y(n_4608)
);

NOR2x1p5_ASAP7_75t_L g4609 ( 
.A(n_4590),
.B(n_4604),
.Y(n_4609)
);

XNOR2x1_ASAP7_75t_L g4610 ( 
.A(n_4599),
.B(n_542),
.Y(n_4610)
);

OAI211xp5_ASAP7_75t_SL g4611 ( 
.A1(n_4581),
.A2(n_546),
.B(n_543),
.C(n_544),
.Y(n_4611)
);

AOI22xp33_ASAP7_75t_SL g4612 ( 
.A1(n_4605),
.A2(n_548),
.B1(n_546),
.B2(n_547),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_4592),
.B(n_549),
.Y(n_4613)
);

NOR2x1_ASAP7_75t_L g4614 ( 
.A(n_4598),
.B(n_549),
.Y(n_4614)
);

AND2x2_ASAP7_75t_L g4615 ( 
.A(n_4591),
.B(n_4596),
.Y(n_4615)
);

NOR3xp33_ASAP7_75t_L g4616 ( 
.A(n_4593),
.B(n_550),
.C(n_551),
.Y(n_4616)
);

INVx2_ASAP7_75t_L g4617 ( 
.A(n_4592),
.Y(n_4617)
);

NAND4xp75_ASAP7_75t_L g4618 ( 
.A(n_4587),
.B(n_553),
.C(n_551),
.D(n_552),
.Y(n_4618)
);

NAND3xp33_ASAP7_75t_SL g4619 ( 
.A(n_4600),
.B(n_552),
.C(n_553),
.Y(n_4619)
);

NOR3x1_ASAP7_75t_L g4620 ( 
.A(n_4582),
.B(n_554),
.C(n_555),
.Y(n_4620)
);

NAND4xp25_ASAP7_75t_L g4621 ( 
.A(n_4589),
.B(n_556),
.C(n_554),
.D(n_555),
.Y(n_4621)
);

AO22x1_ASAP7_75t_L g4622 ( 
.A1(n_4606),
.A2(n_4603),
.B1(n_4592),
.B2(n_4594),
.Y(n_4622)
);

INVxp67_ASAP7_75t_L g4623 ( 
.A(n_4597),
.Y(n_4623)
);

NOR3xp33_ASAP7_75t_L g4624 ( 
.A(n_4588),
.B(n_557),
.C(n_558),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_SL g4625 ( 
.A(n_4601),
.B(n_557),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4585),
.B(n_558),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4586),
.B(n_559),
.Y(n_4627)
);

NOR2x1_ASAP7_75t_L g4628 ( 
.A(n_4595),
.B(n_559),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4602),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4583),
.Y(n_4630)
);

NAND4xp75_ASAP7_75t_L g4631 ( 
.A(n_4605),
.B(n_562),
.C(n_560),
.D(n_561),
.Y(n_4631)
);

AOI22xp5_ASAP7_75t_L g4632 ( 
.A1(n_4582),
.A2(n_566),
.B1(n_562),
.B2(n_564),
.Y(n_4632)
);

AOI22xp5_ASAP7_75t_L g4633 ( 
.A1(n_4630),
.A2(n_568),
.B1(n_564),
.B2(n_567),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4608),
.Y(n_4634)
);

AOI22xp5_ASAP7_75t_L g4635 ( 
.A1(n_4616),
.A2(n_573),
.B1(n_567),
.B2(n_571),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_4617),
.B(n_571),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4628),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_4609),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4613),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4626),
.B(n_574),
.Y(n_4640)
);

HB1xp67_ASAP7_75t_L g4641 ( 
.A(n_4614),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4631),
.Y(n_4642)
);

INVx2_ASAP7_75t_L g4643 ( 
.A(n_4610),
.Y(n_4643)
);

INVxp67_ASAP7_75t_SL g4644 ( 
.A(n_4627),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4625),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4618),
.Y(n_4646)
);

AOI22xp5_ASAP7_75t_L g4647 ( 
.A1(n_4624),
.A2(n_578),
.B1(n_575),
.B2(n_577),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4623),
.Y(n_4648)
);

AO22x1_ASAP7_75t_L g4649 ( 
.A1(n_4620),
.A2(n_578),
.B1(n_575),
.B2(n_577),
.Y(n_4649)
);

AOI22xp5_ASAP7_75t_L g4650 ( 
.A1(n_4632),
.A2(n_579),
.B1(n_580),
.B2(n_581),
.Y(n_4650)
);

AOI22xp5_ASAP7_75t_L g4651 ( 
.A1(n_4621),
.A2(n_579),
.B1(n_580),
.B2(n_581),
.Y(n_4651)
);

OAI21xp5_ASAP7_75t_L g4652 ( 
.A1(n_4612),
.A2(n_582),
.B(n_583),
.Y(n_4652)
);

AOI22xp5_ASAP7_75t_L g4653 ( 
.A1(n_4619),
.A2(n_582),
.B1(n_583),
.B2(n_584),
.Y(n_4653)
);

INVx1_ASAP7_75t_SL g4654 ( 
.A(n_4615),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4607),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4611),
.Y(n_4656)
);

BUFx4f_ASAP7_75t_SL g4657 ( 
.A(n_4654),
.Y(n_4657)
);

BUFx2_ASAP7_75t_L g4658 ( 
.A(n_4636),
.Y(n_4658)
);

NAND4xp75_ASAP7_75t_L g4659 ( 
.A(n_4633),
.B(n_4629),
.C(n_4622),
.D(n_589),
.Y(n_4659)
);

NAND3x1_ASAP7_75t_L g4660 ( 
.A(n_4656),
.B(n_4652),
.C(n_4634),
.Y(n_4660)
);

NOR3xp33_ASAP7_75t_L g4661 ( 
.A(n_4649),
.B(n_586),
.C(n_587),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4640),
.Y(n_4662)
);

NAND4xp75_ASAP7_75t_L g4663 ( 
.A(n_4647),
.B(n_586),
.C(n_589),
.D(n_590),
.Y(n_4663)
);

NOR3xp33_ASAP7_75t_L g4664 ( 
.A(n_4648),
.B(n_592),
.C(n_593),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4651),
.Y(n_4665)
);

NOR4xp75_ASAP7_75t_SL g4666 ( 
.A(n_4653),
.B(n_593),
.C(n_595),
.D(n_596),
.Y(n_4666)
);

OR2x2_ASAP7_75t_L g4667 ( 
.A(n_4638),
.B(n_595),
.Y(n_4667)
);

NOR2xp33_ASAP7_75t_L g4668 ( 
.A(n_4637),
.B(n_596),
.Y(n_4668)
);

AOI31xp33_ASAP7_75t_L g4669 ( 
.A1(n_4642),
.A2(n_597),
.A3(n_598),
.B(n_599),
.Y(n_4669)
);

AND2x2_ASAP7_75t_SL g4670 ( 
.A(n_4655),
.B(n_598),
.Y(n_4670)
);

NOR4xp25_ASAP7_75t_L g4671 ( 
.A(n_4646),
.B(n_600),
.C(n_601),
.D(n_602),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_4635),
.Y(n_4672)
);

NOR3xp33_ASAP7_75t_L g4673 ( 
.A(n_4644),
.B(n_600),
.C(n_601),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4641),
.Y(n_4674)
);

CKINVDCx16_ASAP7_75t_R g4675 ( 
.A(n_4667),
.Y(n_4675)
);

NOR2xp67_ASAP7_75t_L g4676 ( 
.A(n_4674),
.B(n_4645),
.Y(n_4676)
);

NOR2x1_ASAP7_75t_L g4677 ( 
.A(n_4659),
.B(n_4665),
.Y(n_4677)
);

AOI222xp33_ASAP7_75t_L g4678 ( 
.A1(n_4657),
.A2(n_4639),
.B1(n_4643),
.B2(n_4650),
.C1(n_605),
.C2(n_606),
.Y(n_4678)
);

CKINVDCx20_ASAP7_75t_R g4679 ( 
.A(n_4658),
.Y(n_4679)
);

CKINVDCx5p33_ASAP7_75t_R g4680 ( 
.A(n_4668),
.Y(n_4680)
);

INVx1_ASAP7_75t_SL g4681 ( 
.A(n_4670),
.Y(n_4681)
);

BUFx2_ASAP7_75t_L g4682 ( 
.A(n_4660),
.Y(n_4682)
);

NAND2xp33_ASAP7_75t_R g4683 ( 
.A(n_4672),
.B(n_602),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4669),
.Y(n_4684)
);

BUFx2_ASAP7_75t_L g4685 ( 
.A(n_4662),
.Y(n_4685)
);

CKINVDCx20_ASAP7_75t_R g4686 ( 
.A(n_4666),
.Y(n_4686)
);

HB1xp67_ASAP7_75t_L g4687 ( 
.A(n_4663),
.Y(n_4687)
);

CKINVDCx5p33_ASAP7_75t_R g4688 ( 
.A(n_4671),
.Y(n_4688)
);

INVx1_ASAP7_75t_SL g4689 ( 
.A(n_4664),
.Y(n_4689)
);

AOI21xp5_ASAP7_75t_L g4690 ( 
.A1(n_4661),
.A2(n_603),
.B(n_604),
.Y(n_4690)
);

NOR2xp33_ASAP7_75t_R g4691 ( 
.A(n_4673),
.B(n_603),
.Y(n_4691)
);

CKINVDCx5p33_ASAP7_75t_R g4692 ( 
.A(n_4691),
.Y(n_4692)
);

INVx1_ASAP7_75t_SL g4693 ( 
.A(n_4685),
.Y(n_4693)
);

NAND3xp33_ASAP7_75t_SL g4694 ( 
.A(n_4688),
.B(n_605),
.C(n_606),
.Y(n_4694)
);

NOR2x1p5_ASAP7_75t_L g4695 ( 
.A(n_4684),
.B(n_607),
.Y(n_4695)
);

CKINVDCx5p33_ASAP7_75t_R g4696 ( 
.A(n_4683),
.Y(n_4696)
);

AND2x2_ASAP7_75t_L g4697 ( 
.A(n_4675),
.B(n_608),
.Y(n_4697)
);

NAND2x1p5_ASAP7_75t_L g4698 ( 
.A(n_4676),
.B(n_608),
.Y(n_4698)
);

HB1xp67_ASAP7_75t_L g4699 ( 
.A(n_4677),
.Y(n_4699)
);

INVx1_ASAP7_75t_SL g4700 ( 
.A(n_4682),
.Y(n_4700)
);

NAND3xp33_ASAP7_75t_L g4701 ( 
.A(n_4678),
.B(n_609),
.C(n_610),
.Y(n_4701)
);

CKINVDCx5p33_ASAP7_75t_R g4702 ( 
.A(n_4686),
.Y(n_4702)
);

CKINVDCx5p33_ASAP7_75t_R g4703 ( 
.A(n_4680),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_L g4704 ( 
.A(n_4690),
.B(n_610),
.Y(n_4704)
);

AOI211xp5_ASAP7_75t_L g4705 ( 
.A1(n_4694),
.A2(n_4689),
.B(n_4687),
.C(n_4681),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_L g4706 ( 
.A(n_4693),
.B(n_4679),
.Y(n_4706)
);

HB1xp67_ASAP7_75t_L g4707 ( 
.A(n_4702),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4698),
.Y(n_4708)
);

OAI22xp5_ASAP7_75t_SL g4709 ( 
.A1(n_4704),
.A2(n_611),
.B1(n_612),
.B2(n_613),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4698),
.Y(n_4710)
);

NOR2x1_ASAP7_75t_L g4711 ( 
.A(n_4701),
.B(n_611),
.Y(n_4711)
);

HB1xp67_ASAP7_75t_L g4712 ( 
.A(n_4699),
.Y(n_4712)
);

OA22x2_ASAP7_75t_L g4713 ( 
.A1(n_4700),
.A2(n_612),
.B1(n_613),
.B2(n_614),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4697),
.Y(n_4714)
);

OAI222xp33_ASAP7_75t_L g4715 ( 
.A1(n_4706),
.A2(n_4696),
.B1(n_4703),
.B2(n_4692),
.C1(n_4695),
.C2(n_618),
.Y(n_4715)
);

AOI22xp33_ASAP7_75t_L g4716 ( 
.A1(n_4712),
.A2(n_614),
.B1(n_615),
.B2(n_616),
.Y(n_4716)
);

AOI21xp5_ASAP7_75t_L g4717 ( 
.A1(n_4707),
.A2(n_616),
.B(n_617),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4713),
.Y(n_4718)
);

XNOR2x1_ASAP7_75t_L g4719 ( 
.A(n_4711),
.B(n_4708),
.Y(n_4719)
);

AOI21xp5_ASAP7_75t_L g4720 ( 
.A1(n_4709),
.A2(n_617),
.B(n_618),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4710),
.Y(n_4721)
);

AOI22xp5_ASAP7_75t_L g4722 ( 
.A1(n_4714),
.A2(n_619),
.B1(n_620),
.B2(n_621),
.Y(n_4722)
);

AOI22xp5_ASAP7_75t_L g4723 ( 
.A1(n_4721),
.A2(n_4705),
.B1(n_621),
.B2(n_622),
.Y(n_4723)
);

INVx1_ASAP7_75t_SL g4724 ( 
.A(n_4719),
.Y(n_4724)
);

OAI21xp5_ASAP7_75t_L g4725 ( 
.A1(n_4720),
.A2(n_619),
.B(n_624),
.Y(n_4725)
);

HB1xp67_ASAP7_75t_L g4726 ( 
.A(n_4724),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4723),
.Y(n_4727)
);

XNOR2xp5_ASAP7_75t_L g4728 ( 
.A(n_4726),
.B(n_4722),
.Y(n_4728)
);

AOI22xp5_ASAP7_75t_L g4729 ( 
.A1(n_4728),
.A2(n_4727),
.B1(n_4718),
.B2(n_4725),
.Y(n_4729)
);

AOI322xp5_ASAP7_75t_L g4730 ( 
.A1(n_4729),
.A2(n_4715),
.A3(n_4717),
.B1(n_4716),
.B2(n_628),
.C1(n_629),
.C2(n_630),
.Y(n_4730)
);

OAI22xp5_ASAP7_75t_L g4731 ( 
.A1(n_4730),
.A2(n_625),
.B1(n_626),
.B2(n_627),
.Y(n_4731)
);

AOI211xp5_ASAP7_75t_L g4732 ( 
.A1(n_4731),
.A2(n_625),
.B(n_626),
.C(n_630),
.Y(n_4732)
);


endmodule