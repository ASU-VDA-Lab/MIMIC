module fake_aes_12534_n_705 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_705);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_705;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g106 ( .A(n_105), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_32), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_21), .Y(n_108) );
NOR2xp67_ASAP7_75t_L g109 ( .A(n_72), .B(n_22), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_65), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_23), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_100), .Y(n_113) );
BUFx10_ASAP7_75t_L g114 ( .A(n_104), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_12), .Y(n_115) );
OR2x2_ASAP7_75t_L g116 ( .A(n_86), .B(n_39), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_68), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_81), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_63), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_20), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_42), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_85), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_4), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_97), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_13), .Y(n_125) );
INVx1_ASAP7_75t_SL g126 ( .A(n_88), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_28), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_5), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_66), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_6), .Y(n_130) );
INVx1_ASAP7_75t_SL g131 ( .A(n_56), .Y(n_131) );
NOR2xp67_ASAP7_75t_L g132 ( .A(n_27), .B(n_48), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_57), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_93), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_96), .Y(n_135) );
INVx1_ASAP7_75t_SL g136 ( .A(n_89), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_78), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_74), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_101), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_47), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_3), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_33), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_34), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_38), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_20), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_82), .Y(n_146) );
INVxp67_ASAP7_75t_L g147 ( .A(n_17), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_83), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_43), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_25), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_125), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_133), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_110), .Y(n_153) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_112), .A2(n_46), .B(n_102), .Y(n_154) );
NOR2x1_ASAP7_75t_L g155 ( .A(n_121), .B(n_0), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_114), .B(n_0), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_144), .B(n_1), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_134), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_106), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_137), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_115), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_106), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_106), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_133), .B(n_1), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_106), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_108), .B(n_2), .Y(n_167) );
CKINVDCx8_ASAP7_75t_R g168 ( .A(n_107), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_153), .B(n_119), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_165), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_153), .B(n_115), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_165), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_165), .Y(n_174) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_165), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_156), .B(n_127), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
OR2x2_ASAP7_75t_L g178 ( .A(n_151), .B(n_123), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_160), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_160), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_160), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_156), .B(n_123), .Y(n_182) );
BUFx10_ASAP7_75t_L g183 ( .A(n_162), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
NAND2xp33_ASAP7_75t_L g185 ( .A(n_159), .B(n_161), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_168), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_163), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_159), .B(n_130), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_163), .Y(n_189) );
OR2x6_ASAP7_75t_L g190 ( .A(n_157), .B(n_111), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_151), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_166), .Y(n_192) );
NAND3xp33_ASAP7_75t_L g193 ( .A(n_161), .B(n_150), .C(n_142), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_169), .B(n_148), .Y(n_194) );
AND2x4_ASAP7_75t_SL g195 ( .A(n_158), .B(n_117), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_166), .Y(n_196) );
NAND3xp33_ASAP7_75t_SL g197 ( .A(n_191), .B(n_168), .C(n_129), .Y(n_197) );
NAND2x1_ASAP7_75t_L g198 ( .A(n_171), .B(n_169), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_172), .B(n_158), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_175), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_171), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_182), .B(n_168), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_178), .B(n_167), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_175), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_178), .B(n_167), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_179), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_188), .B(n_152), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_183), .B(n_130), .Y(n_209) );
NAND2xp33_ASAP7_75t_L g210 ( .A(n_173), .B(n_116), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_173), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_174), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_181), .Y(n_213) );
NOR2xp33_ASAP7_75t_SL g214 ( .A(n_175), .B(n_186), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_174), .A2(n_154), .B(n_152), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_183), .B(n_145), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_170), .B(n_107), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_183), .B(n_176), .Y(n_218) );
AND2x6_ASAP7_75t_SL g219 ( .A(n_190), .B(n_120), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_190), .A2(n_128), .B1(n_141), .B2(n_145), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_185), .B(n_113), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_194), .B(n_113), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_177), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_186), .A2(n_147), .B1(n_155), .B2(n_138), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_181), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_183), .B(n_122), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_180), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_190), .A2(n_155), .B1(n_138), .B2(n_135), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_177), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_190), .B(n_154), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_195), .B(n_122), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_204), .B(n_190), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_230), .B(n_177), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_204), .A2(n_195), .B1(n_193), .B2(n_143), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_202), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_206), .B(n_114), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_206), .A2(n_193), .B1(n_143), .B2(n_139), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_209), .A2(n_139), .B1(n_135), .B2(n_146), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_209), .B(n_146), .Y(n_239) );
NAND2x1p5_ASAP7_75t_L g240 ( .A(n_205), .B(n_154), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_215), .A2(n_196), .B(n_192), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_198), .A2(n_196), .B(n_192), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_218), .B(n_114), .Y(n_243) );
INVx2_ASAP7_75t_SL g244 ( .A(n_216), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_198), .Y(n_245) );
INVxp67_ASAP7_75t_L g246 ( .A(n_216), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_229), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_205), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_201), .A2(n_112), .B(n_149), .C(n_132), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_201), .A2(n_149), .B1(n_106), .B2(n_166), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_230), .A2(n_187), .B(n_184), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_202), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_199), .B(n_118), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_203), .B(n_126), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_226), .B(n_131), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_211), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_211), .A2(n_136), .B1(n_109), .B2(n_184), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_230), .B(n_180), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_205), .B(n_2), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_212), .A2(n_189), .B(n_187), .Y(n_260) );
AOI22xp33_ASAP7_75t_SL g261 ( .A1(n_220), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_261) );
INVxp67_ASAP7_75t_SL g262 ( .A(n_205), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_251), .A2(n_230), .B(n_212), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_236), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_258), .A2(n_210), .B(n_208), .Y(n_265) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_241), .A2(n_223), .B(n_207), .Y(n_266) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_240), .A2(n_223), .B(n_207), .Y(n_267) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_249), .A2(n_220), .A3(n_228), .B(n_213), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g269 ( .A1(n_246), .A2(n_224), .B(n_197), .C(n_222), .Y(n_269) );
CKINVDCx16_ASAP7_75t_R g270 ( .A(n_239), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_235), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_235), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_232), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_256), .Y(n_274) );
INVx6_ASAP7_75t_L g275 ( .A(n_248), .Y(n_275) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_240), .A2(n_202), .B(n_207), .Y(n_276) );
AO31x2_ASAP7_75t_L g277 ( .A1(n_252), .A2(n_225), .A3(n_213), .B(n_227), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_244), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_252), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_238), .A2(n_231), .B1(n_200), .B2(n_214), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_234), .B(n_217), .Y(n_281) );
AO21x1_ASAP7_75t_L g282 ( .A1(n_233), .A2(n_214), .B(n_225), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_258), .A2(n_221), .B(n_200), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_233), .A2(n_229), .B(n_225), .Y(n_284) );
NAND3xp33_ASAP7_75t_SL g285 ( .A(n_261), .B(n_219), .C(n_213), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_242), .A2(n_229), .B(n_227), .Y(n_286) );
AO31x2_ASAP7_75t_L g287 ( .A1(n_259), .A2(n_227), .A3(n_189), .B(n_164), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_270), .B(n_259), .Y(n_288) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_276), .A2(n_260), .B(n_245), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_263), .A2(n_255), .B(n_247), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_271), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_286), .A2(n_247), .B(n_243), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_277), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_275), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_282), .A2(n_250), .B(n_257), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_273), .B(n_237), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_274), .B(n_254), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_271), .B(n_248), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_277), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_265), .A2(n_247), .B(n_254), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_284), .A2(n_247), .B(n_262), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_277), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_267), .A2(n_250), .B(n_253), .Y(n_303) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_266), .A2(n_229), .B(n_164), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_281), .A2(n_219), .B(n_229), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_266), .A2(n_229), .B(n_164), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_277), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_279), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_266), .A2(n_164), .B(n_52), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_298), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_304), .Y(n_311) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_306), .A2(n_285), .B(n_283), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_296), .B(n_264), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_304), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_298), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_302), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_293), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_296), .B(n_278), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_302), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_293), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_298), .Y(n_321) );
AO21x2_ASAP7_75t_L g322 ( .A1(n_299), .A2(n_281), .B(n_272), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_308), .B(n_268), .Y(n_323) );
OR2x6_ASAP7_75t_L g324 ( .A(n_305), .B(n_299), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_291), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_298), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_307), .B(n_272), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_291), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_289), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_307), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_291), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_308), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_302), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_289), .B(n_287), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_295), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_317), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_311), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_311), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_327), .B(n_288), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_317), .B(n_287), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_314), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_314), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_320), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_331), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_332), .B(n_268), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_318), .A2(n_305), .B1(n_297), .B2(n_294), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_331), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_314), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_320), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_328), .B(n_287), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_330), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_323), .B(n_297), .C(n_300), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_330), .B(n_287), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_316), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_323), .B(n_295), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_325), .B(n_295), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_332), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_329), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_327), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_329), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_325), .B(n_295), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_325), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_333), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_315), .B(n_268), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_333), .B(n_292), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_316), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_333), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_322), .B(n_268), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_315), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_334), .B(n_309), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_322), .B(n_290), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_324), .B(n_322), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_315), .B(n_294), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_322), .B(n_294), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_315), .B(n_303), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_334), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_326), .B(n_303), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_324), .B(n_278), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_352), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_361), .B(n_313), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_361), .B(n_310), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_366), .B(n_324), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_366), .B(n_324), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_342), .B(n_324), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_356), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_360), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_359), .B(n_321), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_359), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_337), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_337), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_345), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_342), .B(n_334), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_371), .B(n_335), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_342), .B(n_319), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_355), .B(n_319), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_364), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_364), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_380), .B(n_6), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_355), .B(n_335), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_345), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_380), .B(n_7), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_340), .B(n_326), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_355), .B(n_335), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_352), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_371), .B(n_335), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_371), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_351), .B(n_329), .Y(n_409) );
NOR2xp67_ASAP7_75t_L g410 ( .A(n_374), .B(n_336), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_347), .B(n_336), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_351), .B(n_336), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_340), .B(n_326), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_353), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_353), .B(n_326), .Y(n_415) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_356), .B(n_329), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_357), .B(n_329), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_357), .B(n_329), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_357), .B(n_312), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_347), .B(n_312), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_368), .B(n_312), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_368), .B(n_312), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_365), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_365), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_369), .B(n_164), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_348), .B(n_7), .Y(n_426) );
INVxp67_ASAP7_75t_L g427 ( .A(n_375), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_375), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_369), .B(n_164), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_377), .B(n_301), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_378), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_358), .B(n_363), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_378), .B(n_8), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_358), .B(n_8), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_376), .B(n_9), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_358), .B(n_9), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_376), .B(n_10), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_363), .B(n_10), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_346), .B(n_11), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_377), .B(n_58), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_363), .B(n_11), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_338), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_346), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_354), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_379), .B(n_12), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_379), .B(n_59), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_391), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_387), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_401), .B(n_374), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_401), .B(n_367), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_391), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_405), .B(n_367), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_442), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_395), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_405), .B(n_367), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_400), .A2(n_349), .B1(n_354), .B2(n_370), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_417), .B(n_367), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_392), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_382), .B(n_370), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_402), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_402), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_442), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_417), .B(n_338), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_390), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_393), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_387), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_418), .B(n_419), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_418), .B(n_338), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_381), .B(n_349), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_403), .A2(n_269), .B(n_373), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_419), .B(n_350), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_443), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_386), .B(n_350), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_386), .B(n_350), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_427), .B(n_13), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_394), .B(n_344), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_394), .B(n_344), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_398), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_414), .Y(n_479) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_439), .B(n_344), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_384), .B(n_343), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_384), .B(n_343), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_436), .B(n_373), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_385), .B(n_396), .Y(n_484) );
INVxp67_ASAP7_75t_SL g485 ( .A(n_410), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_385), .B(n_396), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_408), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_436), .B(n_343), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_397), .B(n_341), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_438), .B(n_341), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_397), .B(n_341), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_406), .B(n_339), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_432), .B(n_339), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_398), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_423), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_399), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_399), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_441), .B(n_372), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_431), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_431), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_424), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_439), .Y(n_502) );
NOR2xp67_ASAP7_75t_SL g503 ( .A(n_435), .B(n_437), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_428), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_411), .B(n_372), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_441), .B(n_372), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_408), .Y(n_507) );
NOR2x1_ASAP7_75t_SL g508 ( .A(n_435), .B(n_362), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_383), .B(n_14), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_395), .B(n_372), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_425), .Y(n_511) );
NOR2xp67_ASAP7_75t_L g512 ( .A(n_421), .B(n_14), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_437), .B(n_15), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_395), .B(n_360), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_407), .B(n_360), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_445), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_407), .B(n_409), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_445), .B(n_15), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_434), .B(n_16), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_407), .B(n_362), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_389), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_409), .B(n_362), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_404), .B(n_362), .Y(n_523) );
BUFx2_ASAP7_75t_SL g524 ( .A(n_440), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_425), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_467), .B(n_484), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_458), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_467), .B(n_413), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_493), .B(n_415), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_504), .Y(n_530) );
NOR4xp25_ASAP7_75t_L g531 ( .A(n_513), .B(n_444), .C(n_426), .D(n_433), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_458), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_492), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_484), .B(n_430), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_469), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_486), .B(n_430), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_472), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_487), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_479), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_479), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_502), .B(n_444), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_487), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_507), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_492), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_500), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_493), .B(n_420), .Y(n_546) );
OAI211xp5_ASAP7_75t_L g547 ( .A1(n_470), .A2(n_433), .B(n_421), .C(n_422), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_469), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_486), .B(n_430), .Y(n_549) );
OAI21xp33_ASAP7_75t_SL g550 ( .A1(n_485), .A2(n_422), .B(n_412), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_521), .B(n_501), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_483), .B(n_488), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_464), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_449), .B(n_412), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_490), .B(n_420), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_449), .B(n_409), .Y(n_556) );
NAND4xp25_ASAP7_75t_L g557 ( .A(n_475), .B(n_446), .C(n_440), .D(n_280), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_507), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_459), .B(n_429), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_465), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_456), .A2(n_446), .B(n_440), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_505), .B(n_416), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_471), .B(n_429), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_503), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_447), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_512), .B(n_446), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_517), .B(n_416), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_471), .B(n_416), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_451), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g570 ( .A1(n_480), .A2(n_388), .B(n_17), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_453), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_460), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_489), .B(n_388), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_524), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_495), .B(n_388), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_454), .B(n_362), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_453), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_461), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_489), .B(n_360), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_516), .B(n_360), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_499), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_448), .B(n_360), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_466), .B(n_16), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_491), .B(n_18), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_476), .B(n_19), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_509), .B(n_19), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_503), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_476), .B(n_21), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_518), .B(n_275), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_491), .B(n_24), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_481), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_481), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_543), .Y(n_593) );
NAND2x1p5_ASAP7_75t_L g594 ( .A(n_574), .B(n_524), .Y(n_594) );
O2A1O1Ixp33_ASAP7_75t_SL g595 ( .A1(n_566), .A2(n_454), .B(n_525), .C(n_511), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_574), .B(n_454), .Y(n_596) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_538), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_551), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_558), .B(n_450), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_541), .B(n_482), .Y(n_600) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_570), .B(n_519), .Y(n_601) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_542), .Y(n_602) );
AOI21xp33_ASAP7_75t_SL g603 ( .A1(n_550), .A2(n_498), .B(n_506), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_564), .A2(n_455), .B1(n_450), .B2(n_452), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_561), .A2(n_452), .B1(n_455), .B2(n_510), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_551), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_571), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_584), .A2(n_457), .B1(n_482), .B2(n_473), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_534), .B(n_474), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_535), .Y(n_610) );
AOI21x1_ASAP7_75t_L g611 ( .A1(n_570), .A2(n_494), .B(n_478), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_541), .B(n_473), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_577), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_548), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_531), .B(n_474), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_537), .B(n_508), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_573), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_530), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_579), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_546), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_586), .A2(n_457), .B1(n_468), .B2(n_463), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_539), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_557), .A2(n_468), .B1(n_463), .B2(n_477), .Y(n_623) );
INVx2_ASAP7_75t_SL g624 ( .A(n_554), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_540), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_547), .A2(n_508), .B(n_514), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_585), .A2(n_477), .B1(n_520), .B2(n_515), .Y(n_627) );
INVx1_ASAP7_75t_SL g628 ( .A(n_582), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_553), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_560), .Y(n_630) );
OAI32xp33_ASAP7_75t_L g631 ( .A1(n_552), .A2(n_523), .A3(n_514), .B1(n_520), .B2(n_515), .Y(n_631) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_583), .A2(n_522), .B(n_497), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_527), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_531), .B(n_497), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_528), .B(n_496), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_532), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_591), .B(n_496), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_585), .A2(n_494), .B1(n_478), .B2(n_462), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_576), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_533), .Y(n_640) );
OAI21xp5_ASAP7_75t_L g641 ( .A1(n_588), .A2(n_462), .B(n_522), .Y(n_641) );
AOI211xp5_ASAP7_75t_SL g642 ( .A1(n_595), .A2(n_588), .B(n_583), .C(n_589), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_615), .B(n_526), .Y(n_643) );
NAND3xp33_ASAP7_75t_SL g644 ( .A(n_603), .B(n_590), .C(n_562), .Y(n_644) );
NAND2xp33_ASAP7_75t_L g645 ( .A(n_593), .B(n_536), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_631), .A2(n_572), .B1(n_565), .B2(n_581), .C(n_569), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_605), .A2(n_557), .B1(n_549), .B2(n_567), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_601), .A2(n_582), .B(n_580), .Y(n_648) );
OA21x2_ASAP7_75t_SL g649 ( .A1(n_593), .A2(n_568), .B(n_563), .Y(n_649) );
CKINVDCx14_ASAP7_75t_R g650 ( .A(n_599), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_623), .B(n_592), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_626), .A2(n_559), .B(n_575), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g653 ( .A1(n_621), .A2(n_555), .B1(n_578), .B2(n_529), .C(n_575), .Y(n_653) );
AOI21xp33_ASAP7_75t_L g654 ( .A1(n_634), .A2(n_576), .B(n_545), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_627), .A2(n_608), .B1(n_616), .B2(n_604), .Y(n_655) );
OAI21xp33_ASAP7_75t_SL g656 ( .A1(n_597), .A2(n_556), .B(n_544), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_618), .A2(n_26), .B1(n_29), .B2(n_30), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_638), .A2(n_31), .B(n_35), .Y(n_658) );
OAI211xp5_ASAP7_75t_L g659 ( .A1(n_641), .A2(n_36), .B(n_37), .C(n_40), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_641), .A2(n_41), .B1(n_44), .B2(n_45), .C(n_49), .Y(n_660) );
NOR2xp33_ASAP7_75t_SL g661 ( .A(n_594), .B(n_50), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_638), .A2(n_51), .B(n_53), .Y(n_662) );
O2A1O1Ixp5_ASAP7_75t_L g663 ( .A1(n_602), .A2(n_54), .B(n_55), .C(n_60), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_632), .A2(n_61), .B1(n_62), .B2(n_64), .C(n_67), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_620), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g666 ( .A1(n_594), .A2(n_69), .B1(n_70), .B2(n_71), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_598), .A2(n_73), .B1(n_75), .B2(n_76), .C(n_77), .Y(n_667) );
XOR2x2_ASAP7_75t_L g668 ( .A(n_624), .B(n_79), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_606), .B(n_80), .Y(n_669) );
NAND2xp33_ASAP7_75t_L g670 ( .A(n_640), .B(n_84), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_610), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_628), .A2(n_87), .B1(n_90), .B2(n_91), .C(n_92), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_611), .B(n_94), .C(n_95), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_614), .B(n_98), .C(n_99), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_596), .A2(n_103), .B(n_637), .Y(n_675) );
OAI31xp33_ASAP7_75t_L g676 ( .A1(n_596), .A2(n_628), .A3(n_639), .B(n_599), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_612), .A2(n_600), .B(n_639), .Y(n_677) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_629), .B(n_630), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_635), .A2(n_607), .B(n_613), .Y(n_679) );
AND5x1_ASAP7_75t_L g680 ( .A(n_617), .B(n_619), .C(n_622), .D(n_625), .E(n_633), .Y(n_680) );
AOI211xp5_ASAP7_75t_SL g681 ( .A1(n_636), .A2(n_595), .B(n_564), .C(n_587), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g682 ( .A(n_656), .B(n_644), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_681), .B(n_676), .C(n_642), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_663), .B(n_672), .C(n_660), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_646), .B(n_673), .C(n_655), .Y(n_685) );
NAND3xp33_ASAP7_75t_SL g686 ( .A(n_661), .B(n_663), .C(n_659), .Y(n_686) );
NAND3xp33_ASAP7_75t_SL g687 ( .A(n_658), .B(n_662), .C(n_664), .Y(n_687) );
OAI211xp5_ASAP7_75t_SL g688 ( .A1(n_647), .A2(n_650), .B(n_654), .C(n_645), .Y(n_688) );
NOR3xp33_ASAP7_75t_L g689 ( .A(n_683), .B(n_666), .C(n_667), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_682), .B(n_665), .Y(n_690) );
NOR2x1_ASAP7_75t_L g691 ( .A(n_686), .B(n_674), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_685), .B(n_680), .Y(n_692) );
INVx3_ASAP7_75t_L g693 ( .A(n_692), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_690), .B(n_643), .Y(n_694) );
XNOR2x1_ASAP7_75t_L g695 ( .A(n_691), .B(n_668), .Y(n_695) );
XNOR2xp5_ASAP7_75t_L g696 ( .A(n_695), .B(n_689), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_693), .B(n_671), .Y(n_697) );
OA21x2_ASAP7_75t_L g698 ( .A1(n_696), .A2(n_694), .B(n_684), .Y(n_698) );
OAI22x1_ASAP7_75t_SL g699 ( .A1(n_697), .A2(n_688), .B1(n_649), .B2(n_687), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_698), .A2(n_697), .B1(n_651), .B2(n_653), .Y(n_700) );
AOI31xp67_ASAP7_75t_L g701 ( .A1(n_699), .A2(n_657), .A3(n_669), .B(n_678), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g702 ( .A1(n_701), .A2(n_670), .B1(n_648), .B2(n_652), .Y(n_702) );
NAND2xp33_ASAP7_75t_R g703 ( .A(n_702), .B(n_700), .Y(n_703) );
AO21x2_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_675), .B(n_677), .Y(n_704) );
AO21x2_ASAP7_75t_L g705 ( .A1(n_704), .A2(n_679), .B(n_609), .Y(n_705) );
endmodule