module fake_netlist_6_546_n_1889 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1889);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1889;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_952;
wire n_725;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1851;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_34),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_66),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_98),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_94),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_119),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_79),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_9),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_17),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_38),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_58),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_7),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_111),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_56),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_7),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_40),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_38),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_45),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_116),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_60),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_12),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_120),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_93),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_90),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_4),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_51),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_71),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_47),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_59),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_5),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_72),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_32),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_26),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_152),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_89),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_74),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_15),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_126),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_26),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_61),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_6),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_151),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_107),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_73),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_62),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_101),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_32),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_21),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_42),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_0),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_143),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_96),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_11),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_53),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_18),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_95),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_142),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_52),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_83),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_22),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_41),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_15),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_134),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_147),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_12),
.Y(n_239)
);

BUFx2_ASAP7_75t_SL g240 ( 
.A(n_104),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_133),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_149),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_46),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_11),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_41),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_1),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_82),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_84),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_54),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_150),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_25),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_55),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_36),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_49),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_91),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_103),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_77),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_76),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_65),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_114),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_141),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_1),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_39),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_4),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_70),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_31),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_30),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_33),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_31),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_40),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_9),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_108),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_86),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_125),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_29),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_48),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_105),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_88),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_30),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_146),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_13),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_64),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_2),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_81),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_34),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_18),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_17),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_78),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_5),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_129),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_16),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_123),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_136),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_14),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_44),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_69),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_85),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_43),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_16),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_3),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_121),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_39),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_10),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_6),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_14),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_115),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_24),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_20),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_28),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_3),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_110),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_263),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_223),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_223),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_211),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_223),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_223),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_160),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_164),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_179),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_211),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_186),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_223),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_199),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_223),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_210),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_223),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_176),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_176),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_176),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_231),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_203),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_176),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_202),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_212),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_214),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_221),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_202),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_202),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_202),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_222),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_302),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_191),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_190),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_246),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_267),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_201),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_224),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_227),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_243),
.Y(n_357)
);

BUFx2_ASAP7_75t_SL g358 ( 
.A(n_231),
.Y(n_358)
);

BUFx2_ASAP7_75t_SL g359 ( 
.A(n_232),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_286),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_243),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_229),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_234),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_232),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_158),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_246),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_235),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_239),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_161),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_267),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_285),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_243),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_236),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_285),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_251),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_268),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_244),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_269),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_191),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_285),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_162),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_271),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_245),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_276),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_283),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_243),
.Y(n_386)
);

INVx4_ASAP7_75t_R g387 ( 
.A(n_208),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_208),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_287),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_343),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_320),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_343),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_332),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_200),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_365),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_343),
.B(n_163),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_318),
.B(n_178),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_333),
.Y(n_405)
);

AND2x2_ASAP7_75t_SL g406 ( 
.A(n_322),
.B(n_200),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_317),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_379),
.B(n_205),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_333),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_327),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_334),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_334),
.Y(n_412)
);

NAND2xp33_ASAP7_75t_L g413 ( 
.A(n_321),
.B(n_169),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_327),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_329),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_337),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_338),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_338),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_314),
.A2(n_178),
.B1(n_291),
.B2(n_310),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_336),
.B(n_180),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_388),
.B(n_163),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_344),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_361),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_316),
.A2(n_310),
.B1(n_291),
.B2(n_169),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_346),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_361),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_347),
.B(n_165),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_349),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_382),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_369),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_389),
.B(n_165),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_381),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_372),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_L g445 ( 
.A(n_323),
.B(n_170),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_386),
.A2(n_300),
.B(n_296),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_352),
.B(n_205),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_386),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_351),
.B(n_167),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_384),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_384),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_385),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_352),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_326),
.A2(n_172),
.B1(n_170),
.B2(n_305),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_447),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

BUFx8_ASAP7_75t_SL g461 ( 
.A(n_402),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_390),
.Y(n_462)
);

AND2x2_ASAP7_75t_SL g463 ( 
.A(n_406),
.B(n_220),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_435),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_429),
.B(n_360),
.Y(n_465)
);

NOR2x1p5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_325),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_400),
.B(n_408),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

BUFx10_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_390),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_400),
.A2(n_168),
.B1(n_311),
.B2(n_309),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_406),
.B(n_371),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_447),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_420),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_435),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_430),
.B(n_325),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_400),
.B(n_328),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_447),
.Y(n_479)
);

NAND2xp33_ASAP7_75t_L g480 ( 
.A(n_408),
.B(n_243),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_426),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_330),
.C(n_328),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_420),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_447),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_391),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_391),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_407),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_407),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_391),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_426),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_430),
.B(n_330),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_425),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_425),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_426),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_393),
.B(n_374),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_393),
.B(n_358),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_425),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_L g502 ( 
.A(n_408),
.B(n_243),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_420),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_SL g504 ( 
.A(n_442),
.B(n_168),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_414),
.B(n_380),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_448),
.B(n_354),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_413),
.B(n_339),
.Y(n_507)
);

NAND2xp33_ASAP7_75t_SL g508 ( 
.A(n_450),
.B(n_172),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_392),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_392),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_436),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_436),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_436),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_397),
.Y(n_514)
);

AND3x2_ASAP7_75t_L g515 ( 
.A(n_414),
.B(n_290),
.C(n_166),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_392),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_445),
.B(n_339),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_437),
.B(n_340),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

INVx8_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_443),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_395),
.B(n_340),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_394),
.A2(n_233),
.B(n_220),
.Y(n_523)
);

INVx6_ASAP7_75t_L g524 ( 
.A(n_395),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_426),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_394),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_403),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_448),
.B(n_355),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_394),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_410),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_396),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_432),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_415),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_432),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_415),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_395),
.B(n_341),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_395),
.B(n_341),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_L g539 ( 
.A1(n_433),
.A2(n_270),
.B1(n_282),
.B2(n_280),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_450),
.B(n_348),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_403),
.B(n_348),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_448),
.A2(n_396),
.B1(n_423),
.B2(n_415),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_423),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_398),
.B(n_363),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_423),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_396),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_437),
.B(n_358),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_398),
.B(n_159),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_398),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_444),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_432),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_444),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_398),
.B(n_363),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_444),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_456),
.B(n_356),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_457),
.B(n_359),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_397),
.B(n_367),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_439),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_444),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_397),
.B(n_367),
.Y(n_560)
);

CKINVDCx6p67_ASAP7_75t_R g561 ( 
.A(n_422),
.Y(n_561)
);

AOI21x1_ASAP7_75t_L g562 ( 
.A1(n_399),
.A2(n_405),
.B(n_401),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_432),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_432),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_454),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_432),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_454),
.Y(n_567)
);

AND3x2_ASAP7_75t_L g568 ( 
.A(n_439),
.B(n_233),
.C(n_294),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_457),
.A2(n_383),
.B1(n_377),
.B2(n_368),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_422),
.B(n_368),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_454),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_397),
.B(n_377),
.Y(n_573)
);

AND3x2_ASAP7_75t_L g574 ( 
.A(n_446),
.B(n_177),
.C(n_174),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_397),
.B(n_383),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_451),
.Y(n_576)
);

INVx8_ASAP7_75t_L g577 ( 
.A(n_416),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_404),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_458),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_451),
.A2(n_455),
.B1(n_453),
.B2(n_452),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_458),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_416),
.B(n_187),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_416),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_458),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_416),
.B(n_273),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_452),
.Y(n_586)
);

BUFx8_ASAP7_75t_SL g587 ( 
.A(n_404),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_440),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_399),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_440),
.Y(n_590)
);

BUFx6f_ASAP7_75t_SL g591 ( 
.A(n_453),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_433),
.B(n_167),
.Y(n_592)
);

BUFx6f_ASAP7_75t_SL g593 ( 
.A(n_455),
.Y(n_593)
);

AO21x2_ASAP7_75t_L g594 ( 
.A1(n_401),
.A2(n_185),
.B(n_184),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_405),
.Y(n_595)
);

AND3x1_ASAP7_75t_L g596 ( 
.A(n_456),
.B(n_304),
.C(n_301),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_434),
.B(n_353),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_434),
.B(n_359),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_438),
.B(n_240),
.Y(n_599)
);

AO21x2_ASAP7_75t_L g600 ( 
.A1(n_409),
.A2(n_266),
.B(n_218),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_440),
.Y(n_601)
);

AND3x2_ASAP7_75t_L g602 ( 
.A(n_438),
.B(n_215),
.C(n_194),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_416),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_416),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_409),
.B(n_362),
.C(n_378),
.Y(n_605)
);

AND2x2_ASAP7_75t_SL g606 ( 
.A(n_416),
.B(n_299),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_411),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_477),
.B(n_171),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_459),
.B(n_440),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_464),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_459),
.B(n_460),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_552),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_555),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_473),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_552),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_555),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_473),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_558),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_460),
.B(n_440),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_464),
.B(n_475),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_554),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_463),
.A2(n_306),
.B1(n_307),
.B2(n_305),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_576),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_506),
.B(n_373),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_554),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_559),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_485),
.B(n_440),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_485),
.B(n_440),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_474),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_559),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_461),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_479),
.B(n_528),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_494),
.B(n_324),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_484),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_503),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_463),
.A2(n_313),
.B1(n_335),
.B2(n_364),
.Y(n_636)
);

AO22x2_ASAP7_75t_L g637 ( 
.A1(n_556),
.A2(n_281),
.B1(n_196),
.B2(n_198),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_467),
.B(n_171),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_506),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_462),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_475),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_529),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_471),
.A2(n_307),
.B1(n_293),
.B2(n_253),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_529),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_467),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_589),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_589),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_467),
.B(n_375),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_479),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_562),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_462),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_478),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_518),
.B(n_173),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_528),
.B(n_173),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_586),
.B(n_376),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_595),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_586),
.B(n_411),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_524),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_507),
.B(n_175),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_586),
.B(n_469),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_595),
.Y(n_661)
);

AND2x6_ASAP7_75t_SL g662 ( 
.A(n_500),
.B(n_207),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_470),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_517),
.B(n_299),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_607),
.Y(n_665)
);

INVx5_ASAP7_75t_L g666 ( 
.A(n_524),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_598),
.B(n_412),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_470),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_607),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_500),
.B(n_412),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_562),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_468),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_596),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_540),
.B(n_175),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_550),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_SL g676 ( 
.A(n_569),
.B(n_265),
.C(n_254),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_469),
.B(n_181),
.Y(n_677)
);

AND2x6_ASAP7_75t_L g678 ( 
.A(n_522),
.B(n_299),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_599),
.B(n_226),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_599),
.B(n_241),
.Y(n_680)
);

INVx8_ASAP7_75t_L g681 ( 
.A(n_500),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_556),
.A2(n_312),
.B1(n_288),
.B2(n_264),
.Y(n_682)
);

INVxp33_ASAP7_75t_L g683 ( 
.A(n_587),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_561),
.A2(n_289),
.B1(n_275),
.B2(n_284),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_468),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_483),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_469),
.B(n_182),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_550),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_500),
.B(n_597),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_541),
.B(n_183),
.Y(n_690)
);

OR2x2_ASAP7_75t_SL g691 ( 
.A(n_482),
.B(n_256),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_599),
.B(n_308),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_565),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_547),
.B(n_417),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_472),
.B(n_188),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_542),
.B(n_449),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_468),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_524),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_599),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_537),
.B(n_189),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_483),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_488),
.B(n_449),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_SL g703 ( 
.A(n_591),
.B(n_192),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_488),
.B(n_449),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_538),
.B(n_193),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_565),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_567),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_567),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_524),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_461),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_SL g711 ( 
.A1(n_592),
.A2(n_206),
.B1(n_204),
.B2(n_197),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_480),
.A2(n_243),
.B1(n_299),
.B2(n_303),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_486),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_572),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_568),
.B(n_417),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_547),
.B(n_418),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_572),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_579),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_486),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_579),
.Y(n_720)
);

OAI21xp33_ASAP7_75t_L g721 ( 
.A1(n_580),
.A2(n_418),
.B(n_431),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_504),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_547),
.B(n_419),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_489),
.B(n_449),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_489),
.B(n_449),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_480),
.A2(n_303),
.B1(n_431),
.B2(n_428),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_581),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_547),
.B(n_419),
.Y(n_728)
);

AND2x6_ASAP7_75t_L g729 ( 
.A(n_544),
.B(n_303),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_515),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_521),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_487),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_508),
.A2(n_258),
.B1(n_209),
.B2(n_213),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_581),
.Y(n_734)
);

AO22x2_ASAP7_75t_L g735 ( 
.A1(n_571),
.A2(n_421),
.B1(n_424),
.B2(n_427),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_465),
.B(n_195),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_553),
.B(n_216),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_468),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_584),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_584),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_487),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_495),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_495),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_545),
.Y(n_744)
);

AND2x6_ASAP7_75t_L g745 ( 
.A(n_557),
.B(n_303),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_560),
.B(n_217),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_573),
.B(n_219),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_575),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_466),
.B(n_421),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_545),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_521),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_606),
.B(n_225),
.Y(n_752)
);

OR2x2_ASAP7_75t_SL g753 ( 
.A(n_561),
.B(n_387),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_594),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_605),
.B(n_602),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_549),
.B(n_449),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_491),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_546),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_539),
.A2(n_260),
.B1(n_230),
.B2(n_237),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_546),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_491),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_496),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_L g763 ( 
.A(n_606),
.B(n_449),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_502),
.B(n_428),
.C(n_427),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_591),
.A2(n_259),
.B1(n_298),
.B2(n_297),
.Y(n_765)
);

INVxp33_ASAP7_75t_L g766 ( 
.A(n_587),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_468),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_496),
.Y(n_768)
);

NAND2x1p5_ASAP7_75t_L g769 ( 
.A(n_549),
.B(n_424),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_497),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_594),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_519),
.B(n_295),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_497),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_SL g774 ( 
.A1(n_578),
.A2(n_292),
.B1(n_279),
.B2(n_278),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_591),
.A2(n_277),
.B1(n_274),
.B2(n_262),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_574),
.B(n_261),
.Y(n_776)
);

XOR2xp5_ASAP7_75t_L g777 ( 
.A(n_578),
.B(n_257),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_508),
.A2(n_255),
.B1(n_252),
.B2(n_250),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_501),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_499),
.A2(n_249),
.B1(n_248),
.B2(n_247),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_645),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_611),
.B(n_519),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_645),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_646),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_647),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_656),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_675),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_688),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_661),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_611),
.B(n_527),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_676),
.A2(n_502),
.B1(n_600),
.B2(n_594),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_632),
.B(n_748),
.Y(n_792)
);

OR2x6_ASAP7_75t_L g793 ( 
.A(n_681),
.B(n_505),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_652),
.B(n_504),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_666),
.A2(n_577),
.B(n_520),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_632),
.B(n_527),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_665),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_676),
.A2(n_600),
.B1(n_582),
.B2(n_585),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_748),
.B(n_531),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_614),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_620),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_652),
.B(n_531),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_669),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_610),
.Y(n_804)
);

NOR2x2_ASAP7_75t_L g805 ( 
.A(n_749),
.B(n_593),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_742),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_610),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_641),
.B(n_600),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_731),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_614),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_754),
.A2(n_771),
.B1(n_653),
.B2(n_659),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_614),
.A2(n_593),
.B1(n_548),
.B2(n_583),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_640),
.Y(n_813)
);

NOR2x1_ASAP7_75t_L g814 ( 
.A(n_660),
.B(n_583),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_617),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_624),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_743),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_617),
.B(n_534),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_617),
.A2(n_593),
.B1(n_548),
.B2(n_603),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_649),
.B(n_534),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_674),
.A2(n_603),
.B(n_604),
.C(n_509),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_609),
.A2(n_536),
.B(n_543),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_649),
.B(n_667),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_SL g824 ( 
.A(n_608),
.B(n_228),
.C(n_238),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_649),
.B(n_536),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_609),
.B(n_543),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_672),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_672),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_709),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_641),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_655),
.Y(n_831)
);

INVx5_ASAP7_75t_L g832 ( 
.A(n_666),
.Y(n_832)
);

INVx5_ASAP7_75t_L g833 ( 
.A(n_666),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_751),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_631),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_694),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_673),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_624),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_619),
.B(n_510),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_673),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_666),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_722),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_619),
.B(n_516),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_627),
.B(n_526),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_633),
.B(n_548),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_639),
.A2(n_532),
.B1(n_530),
.B2(n_511),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_654),
.B(n_514),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_695),
.A2(n_722),
.B1(n_644),
.B2(n_642),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_658),
.B(n_476),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_627),
.B(n_501),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_744),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_628),
.B(n_511),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_651),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_750),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_648),
.B(n_512),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_715),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_613),
.A2(n_512),
.B1(n_513),
.B2(n_588),
.Y(n_857)
);

AND2x2_ASAP7_75t_SL g858 ( 
.A(n_636),
.B(n_514),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_691),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_736),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_710),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_672),
.Y(n_862)
);

NAND2xp33_ASAP7_75t_SL g863 ( 
.A(n_689),
.B(n_242),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_657),
.Y(n_864)
);

INVxp67_ASAP7_75t_SL g865 ( 
.A(n_709),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_663),
.Y(n_866)
);

NAND3xp33_ASAP7_75t_SL g867 ( 
.A(n_690),
.B(n_513),
.C(n_514),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_685),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_618),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_668),
.Y(n_870)
);

NOR3xp33_ASAP7_75t_SL g871 ( 
.A(n_682),
.B(n_0),
.C(n_2),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_616),
.A2(n_601),
.B1(n_493),
.B2(n_588),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_628),
.B(n_601),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_749),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_715),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_686),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_716),
.B(n_601),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_670),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_623),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_629),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_696),
.B(n_533),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_696),
.B(n_533),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_716),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_634),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_635),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_658),
.B(n_590),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_780),
.B(n_535),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_701),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_723),
.B(n_749),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_698),
.A2(n_520),
.B(n_577),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_638),
.B(n_8),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_713),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_753),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_730),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_728),
.A2(n_533),
.B1(n_588),
.B2(n_493),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_698),
.B(n_590),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_719),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_758),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_760),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_681),
.B(n_699),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_671),
.B(n_525),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_650),
.B(n_525),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_637),
.A2(n_525),
.B1(n_493),
.B2(n_498),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_723),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_732),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_685),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_693),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_755),
.B(n_679),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_780),
.B(n_590),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_755),
.B(n_551),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_682),
.B(n_551),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_706),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_746),
.A2(n_535),
.B1(n_498),
.B2(n_551),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_707),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_708),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_685),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_714),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_717),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_679),
.B(n_535),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_718),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_L g921 ( 
.A(n_765),
.B(n_498),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_697),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_720),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_681),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_727),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_752),
.A2(n_563),
.B1(n_564),
.B2(n_566),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_622),
.B(n_563),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_699),
.B(n_563),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_734),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_711),
.B(n_566),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_739),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_680),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_662),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_735),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_650),
.B(n_564),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_776),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_777),
.B(n_566),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_776),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_740),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_726),
.B(n_564),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_697),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_697),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_712),
.A2(n_590),
.B1(n_481),
.B2(n_570),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_680),
.B(n_590),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_726),
.B(n_492),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_712),
.B(n_492),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_761),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_735),
.B(n_492),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_637),
.A2(n_492),
.B1(n_570),
.B2(n_481),
.Y(n_949)
);

INVx5_ASAP7_75t_L g950 ( 
.A(n_767),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_692),
.B(n_492),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_735),
.A2(n_570),
.B1(n_481),
.B2(n_476),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_692),
.B(n_570),
.Y(n_953)
);

NAND2x2_ASAP7_75t_L g954 ( 
.A(n_774),
.B(n_523),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_741),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_759),
.B(n_476),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_767),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_767),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_637),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_763),
.B(n_570),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_762),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_733),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_778),
.B(n_481),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_756),
.A2(n_577),
.B(n_520),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_768),
.Y(n_965)
);

OR2x6_ASAP7_75t_L g966 ( 
.A(n_677),
.B(n_577),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_763),
.B(n_481),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_772),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_700),
.A2(n_476),
.B1(n_520),
.B2(n_490),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_687),
.B(n_476),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_759),
.B(n_8),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_779),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_804),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_855),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_968),
.B(n_769),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_834),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_800),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_784),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_902),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_811),
.B(n_769),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_830),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_845),
.A2(n_705),
.B1(n_737),
.B2(n_747),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_902),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_935),
.Y(n_984)
);

NOR2x1p5_ASAP7_75t_L g985 ( 
.A(n_809),
.B(n_683),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_869),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_834),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_968),
.B(n_792),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_864),
.B(n_622),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_971),
.A2(n_684),
.B1(n_721),
.B2(n_643),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_792),
.B(n_772),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_879),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_827),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_823),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_823),
.B(n_757),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_935),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_800),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_859),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_901),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_806),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_827),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_807),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_827),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_817),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_836),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_851),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_901),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_889),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_860),
.B(n_864),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_831),
.A2(n_703),
.B1(n_775),
.B2(n_765),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_924),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_835),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_802),
.B(n_773),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_854),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_787),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_813),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_889),
.Y(n_1017)
);

CKINVDCx8_ASAP7_75t_R g1018 ( 
.A(n_908),
.Y(n_1018)
);

AND2x6_ASAP7_75t_L g1019 ( 
.A(n_952),
.B(n_756),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_802),
.B(n_770),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_831),
.B(n_630),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_801),
.B(n_684),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_847),
.B(n_626),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_861),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_853),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_848),
.B(n_612),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_788),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_810),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_880),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_878),
.A2(n_775),
.B1(n_729),
.B2(n_678),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_866),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_842),
.B(n_766),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_785),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_799),
.B(n_625),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_858),
.B(n_615),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_786),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_789),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_799),
.B(n_621),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_884),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_908),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_808),
.B(n_704),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_910),
.B(n_704),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_885),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_883),
.B(n_764),
.Y(n_1044)
);

INVxp67_ASAP7_75t_SL g1045 ( 
.A(n_943),
.Y(n_1045)
);

AND2x6_ASAP7_75t_L g1046 ( 
.A(n_812),
.B(n_725),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_950),
.Y(n_1047)
);

AND2x4_ASAP7_75t_SL g1048 ( 
.A(n_900),
.B(n_738),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_904),
.B(n_764),
.Y(n_1049)
);

INVx3_ASAP7_75t_SL g1050 ( 
.A(n_805),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_870),
.Y(n_1051)
);

BUFx4f_ASAP7_75t_L g1052 ( 
.A(n_793),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_862),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_862),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_910),
.B(n_702),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_911),
.B(n_702),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_832),
.B(n_725),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_934),
.A2(n_643),
.B1(n_664),
.B2(n_729),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_837),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_839),
.B(n_724),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_840),
.B(n_724),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_898),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_937),
.B(n_729),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_839),
.B(n_729),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_875),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_843),
.B(n_678),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_876),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_899),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_888),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_843),
.B(n_678),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_950),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_844),
.B(n_678),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_810),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_892),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_894),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_832),
.B(n_738),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_907),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_897),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_912),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_815),
.Y(n_1080)
);

INVxp67_ASAP7_75t_SL g1081 ( 
.A(n_943),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_874),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_914),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_905),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_794),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_844),
.B(n_664),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_832),
.B(n_490),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_862),
.Y(n_1088)
);

INVx3_ASAP7_75t_SL g1089 ( 
.A(n_933),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_959),
.B(n_10),
.Y(n_1090)
);

BUFx4f_ASAP7_75t_L g1091 ( 
.A(n_793),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_955),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_815),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_816),
.B(n_19),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_906),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_900),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_873),
.B(n_664),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_856),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_900),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_873),
.B(n_664),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_832),
.B(n_490),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_796),
.B(n_745),
.Y(n_1102)
);

NAND2xp33_ASAP7_75t_L g1103 ( 
.A(n_833),
.B(n_745),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_915),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_833),
.B(n_490),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_917),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_962),
.A2(n_838),
.B1(n_930),
.B2(n_824),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_932),
.B(n_68),
.Y(n_1108)
);

OR2x6_ASAP7_75t_L g1109 ( 
.A(n_793),
.B(n_523),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_918),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_920),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_923),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_906),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_796),
.B(n_745),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_863),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_906),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_881),
.B(n_745),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_925),
.Y(n_1118)
);

AND2x4_ASAP7_75t_SL g1119 ( 
.A(n_877),
.B(n_916),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_916),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_881),
.B(n_490),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_882),
.B(n_19),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_916),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_929),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_882),
.B(n_20),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1060),
.A2(n_833),
.B(n_890),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1047),
.Y(n_1127)
);

AOI21x1_ASAP7_75t_L g1128 ( 
.A1(n_980),
.A2(n_1035),
.B(n_1117),
.Y(n_1128)
);

AND2x6_ASAP7_75t_L g1129 ( 
.A(n_979),
.B(n_948),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_1024),
.Y(n_1130)
);

OAI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_987),
.A2(n_891),
.B1(n_893),
.B2(n_938),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1022),
.B(n_871),
.Y(n_1132)
);

BUFx10_ASAP7_75t_L g1133 ( 
.A(n_1032),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_976),
.B(n_877),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_990),
.A2(n_956),
.B(n_887),
.C(n_791),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_SL g1136 ( 
.A1(n_980),
.A2(n_948),
.B(n_909),
.C(n_824),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_993),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1110),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_986),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_990),
.A2(n_954),
.B1(n_781),
.B2(n_783),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_973),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1110),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1096),
.B(n_936),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_981),
.Y(n_1144)
);

INVx8_ASAP7_75t_L g1145 ( 
.A(n_1001),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_989),
.B(n_919),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_973),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_992),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1032),
.A2(n_919),
.B1(n_970),
.B2(n_966),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_1096),
.B(n_966),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_991),
.B(n_782),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1111),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1045),
.A2(n_1081),
.B1(n_988),
.B2(n_989),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_993),
.Y(n_1154)
);

HAxp5_ASAP7_75t_L g1155 ( 
.A(n_985),
.B(n_21),
.CON(n_1155),
.SN(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1012),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_993),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1029),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1039),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_994),
.B(n_782),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1099),
.B(n_797),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1011),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_1005),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_1005),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1085),
.A2(n_928),
.B1(n_927),
.B2(n_970),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1043),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_1009),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1002),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1000),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_1107),
.B(n_798),
.C(n_821),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1004),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_1047),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1006),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1045),
.A2(n_949),
.B1(n_946),
.B2(n_945),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1099),
.B(n_803),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1010),
.A2(n_819),
.B1(n_966),
.B2(n_939),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1014),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_998),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_982),
.A2(n_921),
.B(n_814),
.C(n_963),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1081),
.A2(n_946),
.B1(n_945),
.B2(n_790),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1008),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_974),
.A2(n_944),
.B1(n_951),
.B2(n_953),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1015),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_974),
.A2(n_972),
.B1(n_965),
.B2(n_961),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1115),
.A2(n_947),
.B1(n_931),
.B2(n_895),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_993),
.Y(n_1186)
);

NOR3xp33_ASAP7_75t_L g1187 ( 
.A(n_1063),
.B(n_867),
.C(n_849),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1017),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1027),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1062),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1059),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_994),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1003),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_975),
.B(n_818),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1065),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1016),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_1001),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_1082),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1044),
.A2(n_867),
.B1(n_903),
.B2(n_825),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_999),
.B(n_790),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1068),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1077),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_1001),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1089),
.Y(n_1204)
);

AOI222xp33_ASAP7_75t_L g1205 ( 
.A1(n_1090),
.A2(n_1091),
.B1(n_1052),
.B2(n_1083),
.C1(n_1079),
.C2(n_1104),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_999),
.B(n_826),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1106),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1056),
.A2(n_833),
.B(n_890),
.Y(n_1208)
);

INVx3_ASAP7_75t_SL g1209 ( 
.A(n_1050),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1061),
.B(n_846),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1023),
.A2(n_795),
.B(n_841),
.Y(n_1211)
);

OAI21xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1035),
.A2(n_940),
.B(n_967),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1011),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1044),
.A2(n_820),
.B1(n_825),
.B2(n_818),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1082),
.B(n_868),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1040),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1003),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1016),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1071),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1049),
.A2(n_820),
.B1(n_872),
.B2(n_960),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1025),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1112),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1090),
.B(n_857),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1116),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1119),
.B(n_868),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1049),
.A2(n_865),
.B1(n_829),
.B2(n_926),
.Y(n_1226)
);

NOR2x1_ASAP7_75t_L g1227 ( 
.A(n_1071),
.B(n_922),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1118),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1007),
.B(n_826),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1119),
.B(n_922),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1021),
.B(n_940),
.Y(n_1231)
);

OAI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1052),
.A2(n_1091),
.B1(n_1018),
.B2(n_1094),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1042),
.A2(n_967),
.B1(n_960),
.B2(n_828),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1098),
.B(n_828),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1124),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1003),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1031),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1048),
.B(n_1108),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1007),
.B(n_850),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1048),
.B(n_941),
.Y(n_1240)
);

BUFx8_ASAP7_75t_SL g1241 ( 
.A(n_1003),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1116),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1108),
.A2(n_886),
.B1(n_896),
.B2(n_913),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1058),
.A2(n_850),
.B1(n_852),
.B2(n_950),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1055),
.A2(n_942),
.B1(n_958),
.B2(n_957),
.Y(n_1245)
);

OAI221xp5_ASAP7_75t_L g1246 ( 
.A1(n_1058),
.A2(n_822),
.B1(n_852),
.B2(n_964),
.C(n_969),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1120),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1041),
.B(n_822),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1122),
.A2(n_950),
.B1(n_958),
.B2(n_957),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_978),
.A2(n_958),
.B1(n_957),
.B2(n_942),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1120),
.Y(n_1251)
);

INVxp67_ASAP7_75t_SL g1252 ( 
.A(n_1073),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1050),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1031),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1053),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1089),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1073),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1051),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1053),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1064),
.A2(n_795),
.B(n_841),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1075),
.A2(n_942),
.B1(n_941),
.B2(n_964),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1093),
.Y(n_1262)
);

NOR2x1_ASAP7_75t_L g1263 ( 
.A(n_1113),
.B(n_941),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1093),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_977),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1053),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_979),
.B(n_22),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1053),
.B(n_75),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_SL g1269 ( 
.A1(n_1030),
.A2(n_67),
.B(n_145),
.C(n_140),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1067),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1069),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_983),
.B(n_984),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1054),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1033),
.A2(n_1036),
.B1(n_1037),
.B2(n_1019),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1001),
.B(n_63),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1266),
.Y(n_1276)
);

BUFx2_ASAP7_75t_SL g1277 ( 
.A(n_1213),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1170),
.A2(n_1114),
.B(n_1102),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1135),
.A2(n_1125),
.B(n_1026),
.C(n_1086),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1192),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1151),
.A2(n_1072),
.B(n_1066),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1179),
.A2(n_1070),
.A3(n_1097),
.B(n_1100),
.Y(n_1282)
);

AO21x2_ASAP7_75t_L g1283 ( 
.A1(n_1170),
.A2(n_1057),
.B(n_1121),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1153),
.B(n_984),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1153),
.A2(n_1205),
.B(n_1136),
.C(n_1176),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1151),
.A2(n_1057),
.B(n_1103),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1208),
.A2(n_1076),
.B(n_1038),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1260),
.A2(n_983),
.B(n_996),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1208),
.A2(n_996),
.A3(n_1013),
.B(n_1020),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1166),
.Y(n_1290)
);

AOI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1260),
.A2(n_1109),
.B(n_1076),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1138),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1126),
.A2(n_1034),
.B(n_995),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1238),
.B(n_1080),
.Y(n_1294)
);

AOI32xp33_ASAP7_75t_L g1295 ( 
.A1(n_1132),
.A2(n_1078),
.A3(n_1092),
.B1(n_1084),
.B2(n_1069),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1126),
.A2(n_1105),
.B(n_1101),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1146),
.B(n_1074),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1167),
.B(n_1074),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1211),
.A2(n_1087),
.B(n_1105),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1211),
.A2(n_1246),
.B(n_1248),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1128),
.A2(n_1087),
.B(n_1101),
.Y(n_1301)
);

CKINVDCx16_ASAP7_75t_R g1302 ( 
.A(n_1156),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1145),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1204),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1155),
.B(n_1078),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1212),
.A2(n_1019),
.B(n_1046),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1223),
.A2(n_1084),
.B1(n_1092),
.B2(n_1123),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1246),
.A2(n_1109),
.B(n_997),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1167),
.A2(n_1109),
.B1(n_977),
.B2(n_997),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1160),
.A2(n_1123),
.B1(n_1054),
.B2(n_1095),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1195),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1144),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1248),
.A2(n_1080),
.B(n_1028),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1180),
.A2(n_1028),
.B(n_1113),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1163),
.B(n_1123),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1142),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1180),
.A2(n_1046),
.B(n_1019),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1139),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1249),
.A2(n_1046),
.B(n_1019),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1160),
.A2(n_1123),
.B1(n_1095),
.B2(n_1088),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1274),
.A2(n_1019),
.B(n_1046),
.Y(n_1321)
);

AOI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1249),
.A2(n_1046),
.B(n_1088),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_SL g1323 ( 
.A1(n_1269),
.A2(n_1095),
.B(n_1088),
.C(n_1054),
.Y(n_1323)
);

OAI21xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1205),
.A2(n_97),
.B(n_156),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1244),
.A2(n_1095),
.B(n_1088),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1244),
.A2(n_1054),
.B(n_57),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1200),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1145),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1172),
.B(n_87),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1163),
.B(n_23),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1232),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1331)
);

CKINVDCx11_ASAP7_75t_R g1332 ( 
.A(n_1209),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1174),
.A2(n_100),
.B(n_128),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1174),
.A2(n_1272),
.B(n_1214),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1147),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1200),
.A2(n_99),
.B(n_122),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1272),
.A2(n_50),
.B(n_118),
.Y(n_1337)
);

AOI21xp33_ASAP7_75t_L g1338 ( 
.A1(n_1194),
.A2(n_27),
.B(n_33),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1148),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1206),
.A2(n_102),
.B(n_117),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1164),
.B(n_35),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1158),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1159),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_SL g1344 ( 
.A1(n_1267),
.A2(n_36),
.B(n_37),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1206),
.A2(n_106),
.B(n_112),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1169),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1229),
.A2(n_139),
.B(n_42),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1268),
.A2(n_37),
.B1(n_43),
.B2(n_1185),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1210),
.A2(n_1165),
.B1(n_1268),
.B2(n_1231),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1267),
.A2(n_1229),
.A3(n_1239),
.B(n_1237),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_SL g1351 ( 
.A1(n_1239),
.A2(n_1243),
.B(n_1261),
.C(n_1222),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1199),
.A2(n_1233),
.B(n_1226),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1238),
.B(n_1215),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1268),
.A2(n_1171),
.B1(n_1207),
.B2(n_1228),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1131),
.A2(n_1187),
.B1(n_1178),
.B2(n_1216),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1191),
.B(n_1168),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1181),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1220),
.A2(n_1140),
.B(n_1129),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1141),
.A2(n_1164),
.B(n_1257),
.C(n_1262),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1270),
.A2(n_1182),
.B(n_1152),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1196),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1173),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1188),
.A2(n_1129),
.B1(n_1253),
.B2(n_1133),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1177),
.A2(n_1202),
.B1(n_1183),
.B2(n_1201),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1149),
.A2(n_1184),
.B(n_1235),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1129),
.B(n_1190),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1215),
.B(n_1143),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1145),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1197),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1189),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1256),
.Y(n_1371)
);

INVx5_ASAP7_75t_L g1372 ( 
.A(n_1197),
.Y(n_1372)
);

AOI222xp33_ASAP7_75t_L g1373 ( 
.A1(n_1134),
.A2(n_1175),
.B1(n_1161),
.B2(n_1143),
.C1(n_1129),
.C2(n_1133),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_1252),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1218),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1203),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1275),
.A2(n_1254),
.B(n_1271),
.Y(n_1377)
);

AOI32xp33_ASAP7_75t_L g1378 ( 
.A1(n_1161),
.A2(n_1175),
.A3(n_1242),
.B1(n_1224),
.B2(n_1234),
.Y(n_1378)
);

CKINVDCx16_ASAP7_75t_R g1379 ( 
.A(n_1130),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1264),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1172),
.A2(n_1150),
.B(n_1275),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1150),
.A2(n_1250),
.B1(n_1245),
.B2(n_1251),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1221),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1258),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1247),
.B(n_1273),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1234),
.A2(n_1265),
.B(n_1230),
.C(n_1225),
.Y(n_1386)
);

AO21x2_ASAP7_75t_L g1387 ( 
.A1(n_1240),
.A2(n_1225),
.B(n_1230),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1227),
.A2(n_1265),
.B(n_1127),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1150),
.B(n_1240),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1241),
.Y(n_1390)
);

NAND2x1p5_ASAP7_75t_L g1391 ( 
.A(n_1172),
.B(n_1203),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1127),
.A2(n_1219),
.B(n_1263),
.Y(n_1392)
);

BUFx2_ASAP7_75t_SL g1393 ( 
.A(n_1162),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1137),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1198),
.A2(n_1172),
.B(n_1219),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1259),
.B(n_1137),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1137),
.A2(n_1154),
.B1(n_1157),
.B2(n_1186),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1154),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1154),
.B(n_1157),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1157),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1186),
.A2(n_1193),
.B(n_1217),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_SL g1402 ( 
.A1(n_1186),
.A2(n_1193),
.B(n_1217),
.C(n_1236),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1193),
.Y(n_1403)
);

NOR2x1_ASAP7_75t_SL g1404 ( 
.A(n_1217),
.B(n_1236),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1236),
.A2(n_1255),
.B1(n_1135),
.B2(n_990),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1255),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1255),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1213),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1146),
.B(n_1132),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1153),
.B(n_1160),
.Y(n_1410)
);

O2A1O1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1135),
.A2(n_653),
.B(n_971),
.C(n_633),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1260),
.A2(n_1126),
.B(n_1211),
.Y(n_1412)
);

AOI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1135),
.A2(n_633),
.B1(n_990),
.B2(n_971),
.C(n_682),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1213),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1195),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1260),
.A2(n_1126),
.B(n_1211),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1260),
.A2(n_1126),
.B(n_1211),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1146),
.B(n_1132),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1260),
.A2(n_1126),
.B(n_1211),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1238),
.B(n_1096),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1318),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1290),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1292),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1332),
.Y(n_1424)
);

AOI21xp33_ASAP7_75t_L g1425 ( 
.A1(n_1411),
.A2(n_1413),
.B(n_1285),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1414),
.Y(n_1426)
);

NOR3xp33_ASAP7_75t_L g1427 ( 
.A(n_1411),
.B(n_1413),
.C(n_1324),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1316),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1389),
.B(n_1387),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1348),
.B(n_1409),
.Y(n_1430)
);

CKINVDCx16_ASAP7_75t_R g1431 ( 
.A(n_1379),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1418),
.B(n_1297),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1305),
.B(n_1298),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1308),
.A2(n_1326),
.B(n_1300),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1348),
.A2(n_1338),
.B1(n_1327),
.B2(n_1349),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1335),
.B(n_1355),
.Y(n_1436)
);

NOR2xp67_ASAP7_75t_L g1437 ( 
.A(n_1371),
.B(n_1408),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1285),
.A2(n_1326),
.B(n_1331),
.C(n_1358),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1327),
.A2(n_1358),
.B1(n_1405),
.B2(n_1306),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1339),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1374),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1389),
.B(n_1387),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1420),
.B(n_1353),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1300),
.A2(n_1286),
.B(n_1351),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1331),
.A2(n_1338),
.B1(n_1344),
.B2(n_1349),
.C(n_1359),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1342),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1352),
.A2(n_1365),
.B1(n_1306),
.B2(n_1405),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1317),
.A2(n_1333),
.B(n_1336),
.C(n_1354),
.Y(n_1448)
);

AOI221xp5_ASAP7_75t_L g1449 ( 
.A1(n_1359),
.A2(n_1279),
.B1(n_1341),
.B2(n_1330),
.C(n_1336),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1373),
.A2(n_1302),
.B1(n_1354),
.B2(n_1363),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1410),
.A2(n_1280),
.B1(n_1370),
.B2(n_1362),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1343),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1378),
.A2(n_1335),
.B1(n_1364),
.B2(n_1410),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1280),
.A2(n_1346),
.B1(n_1357),
.B2(n_1312),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1356),
.B(n_1374),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1398),
.Y(n_1456)
);

NAND2x1p5_ASAP7_75t_L g1457 ( 
.A(n_1372),
.B(n_1381),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1420),
.B(n_1353),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1366),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1373),
.A2(n_1311),
.B1(n_1382),
.B2(n_1304),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1367),
.B(n_1315),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1366),
.Y(n_1462)
);

NAND2xp33_ASAP7_75t_SL g1463 ( 
.A(n_1276),
.B(n_1390),
.Y(n_1463)
);

AO31x2_ASAP7_75t_L g1464 ( 
.A1(n_1308),
.A2(n_1313),
.A3(n_1281),
.B(n_1286),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1367),
.B(n_1380),
.Y(n_1465)
);

BUFx8_ASAP7_75t_SL g1466 ( 
.A(n_1276),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1277),
.A2(n_1276),
.B1(n_1393),
.B2(n_1381),
.Y(n_1467)
);

CKINVDCx11_ASAP7_75t_R g1468 ( 
.A(n_1415),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1412),
.A2(n_1419),
.B(n_1416),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1386),
.B(n_1294),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1364),
.A2(n_1382),
.B1(n_1380),
.B2(n_1284),
.Y(n_1471)
);

OAI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1284),
.A2(n_1329),
.B1(n_1321),
.B2(n_1307),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1375),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1361),
.B(n_1384),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1385),
.B(n_1307),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1321),
.A2(n_1334),
.B1(n_1278),
.B2(n_1283),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1383),
.B(n_1281),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1417),
.A2(n_1293),
.B(n_1313),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1294),
.B(n_1350),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1295),
.B(n_1320),
.C(n_1310),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1368),
.Y(n_1481)
);

AO31x2_ASAP7_75t_L g1482 ( 
.A1(n_1310),
.A2(n_1320),
.A3(n_1397),
.B(n_1291),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1403),
.B(n_1406),
.Y(n_1483)
);

BUFx12f_ASAP7_75t_L g1484 ( 
.A(n_1368),
.Y(n_1484)
);

NOR4xp25_ASAP7_75t_L g1485 ( 
.A(n_1309),
.B(n_1323),
.C(n_1407),
.D(n_1400),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1350),
.B(n_1394),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1368),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1309),
.A2(n_1322),
.B(n_1296),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1396),
.B(n_1399),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1289),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1399),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1360),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1289),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1319),
.A2(n_1329),
.B1(n_1347),
.B2(n_1283),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1391),
.A2(n_1404),
.B(n_1369),
.Y(n_1495)
);

INVxp33_ASAP7_75t_L g1496 ( 
.A(n_1396),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_SL g1497 ( 
.A1(n_1397),
.A2(n_1328),
.B(n_1303),
.C(n_1372),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1303),
.Y(n_1498)
);

NAND2x1_ASAP7_75t_L g1499 ( 
.A(n_1369),
.B(n_1376),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1395),
.B(n_1392),
.Y(n_1500)
);

NOR3xp33_ASAP7_75t_SL g1501 ( 
.A(n_1340),
.B(n_1345),
.C(n_1337),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1401),
.B(n_1395),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1287),
.A2(n_1288),
.B1(n_1314),
.B2(n_1376),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1391),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1388),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1282),
.B(n_1289),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1377),
.B(n_1282),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1282),
.B(n_1325),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1287),
.B(n_1372),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1301),
.B(n_1299),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1402),
.B(n_1297),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1368),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1290),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1297),
.B(n_1298),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1413),
.A2(n_971),
.B1(n_1348),
.B2(n_990),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1409),
.B(n_1418),
.Y(n_1516)
);

OAI211xp5_ASAP7_75t_L g1517 ( 
.A1(n_1413),
.A2(n_1331),
.B(n_1411),
.C(n_971),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1411),
.B(n_1146),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1318),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1413),
.A2(n_971),
.B1(n_1348),
.B2(n_990),
.Y(n_1520)
);

NOR2x1p5_ASAP7_75t_L g1521 ( 
.A(n_1276),
.B(n_1253),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_SL g1522 ( 
.A(n_1411),
.B(n_1413),
.C(n_1205),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1413),
.A2(n_971),
.B1(n_1348),
.B2(n_990),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1409),
.B(n_1418),
.Y(n_1524)
);

OAI211xp5_ASAP7_75t_L g1525 ( 
.A1(n_1413),
.A2(n_1331),
.B(n_1411),
.C(n_971),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1312),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1413),
.A2(n_971),
.B1(n_1348),
.B2(n_990),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1412),
.A2(n_1417),
.B(n_1416),
.Y(n_1528)
);

OAI222xp33_ASAP7_75t_L g1529 ( 
.A1(n_1348),
.A2(n_1411),
.B1(n_1331),
.B2(n_1285),
.C1(n_1327),
.C2(n_990),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1368),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1414),
.Y(n_1531)
);

BUFx12f_ASAP7_75t_L g1532 ( 
.A(n_1332),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1409),
.B(n_1418),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1411),
.A2(n_1135),
.B(n_845),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1389),
.B(n_1387),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1398),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1522),
.A2(n_1460),
.B1(n_1450),
.B2(n_1425),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1421),
.Y(n_1538)
);

CKINVDCx16_ASAP7_75t_R g1539 ( 
.A(n_1431),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1455),
.B(n_1433),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1461),
.B(n_1465),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1429),
.B(n_1442),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1441),
.Y(n_1543)
);

CKINVDCx16_ASAP7_75t_R g1544 ( 
.A(n_1424),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1522),
.A2(n_1523),
.B1(n_1527),
.B2(n_1515),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1441),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1489),
.B(n_1432),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1457),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1459),
.Y(n_1549)
);

NAND2xp33_ASAP7_75t_R g1550 ( 
.A(n_1470),
.B(n_1501),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1440),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1446),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1452),
.Y(n_1553)
);

NAND3xp33_ASAP7_75t_SL g1554 ( 
.A(n_1515),
.B(n_1527),
.C(n_1523),
.Y(n_1554)
);

OR2x6_ASAP7_75t_L g1555 ( 
.A(n_1444),
.B(n_1457),
.Y(n_1555)
);

OR2x6_ASAP7_75t_L g1556 ( 
.A(n_1534),
.B(n_1448),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1516),
.B(n_1524),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1533),
.B(n_1429),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_R g1559 ( 
.A(n_1463),
.B(n_1487),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1442),
.B(n_1535),
.Y(n_1560)
);

NOR3xp33_ASAP7_75t_SL g1561 ( 
.A(n_1517),
.B(n_1525),
.C(n_1529),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1519),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1466),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1535),
.B(n_1462),
.Y(n_1564)
);

INVx4_ASAP7_75t_L g1565 ( 
.A(n_1504),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1479),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1500),
.B(n_1502),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1477),
.Y(n_1568)
);

NOR3xp33_ASAP7_75t_SL g1569 ( 
.A(n_1529),
.B(n_1449),
.C(n_1438),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1483),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1503),
.A2(n_1528),
.B(n_1478),
.Y(n_1571)
);

CKINVDCx16_ASAP7_75t_R g1572 ( 
.A(n_1532),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_R g1573 ( 
.A(n_1491),
.B(n_1468),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1520),
.A2(n_1427),
.B1(n_1435),
.B2(n_1439),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1514),
.B(n_1453),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1480),
.B(n_1448),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1520),
.A2(n_1427),
.B1(n_1435),
.B2(n_1439),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1473),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1518),
.A2(n_1445),
.B1(n_1430),
.B2(n_1436),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1492),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1500),
.B(n_1508),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1486),
.B(n_1454),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1454),
.B(n_1475),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1422),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_R g1585 ( 
.A(n_1484),
.B(n_1481),
.Y(n_1585)
);

CKINVDCx16_ASAP7_75t_R g1586 ( 
.A(n_1531),
.Y(n_1586)
);

OR2x6_ASAP7_75t_L g1587 ( 
.A(n_1509),
.B(n_1495),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_R g1588 ( 
.A(n_1481),
.B(n_1530),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1475),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1518),
.B(n_1474),
.Y(n_1590)
);

CKINVDCx16_ASAP7_75t_R g1591 ( 
.A(n_1456),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1471),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1521),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1506),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1423),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1496),
.B(n_1526),
.Y(n_1596)
);

OR2x6_ASAP7_75t_L g1597 ( 
.A(n_1505),
.B(n_1507),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1451),
.B(n_1513),
.Y(n_1598)
);

NOR3xp33_ASAP7_75t_SL g1599 ( 
.A(n_1438),
.B(n_1430),
.C(n_1511),
.Y(n_1599)
);

XOR2xp5_ASAP7_75t_L g1600 ( 
.A(n_1443),
.B(n_1458),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1510),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_R g1602 ( 
.A(n_1530),
.B(n_1426),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1434),
.A2(n_1447),
.B1(n_1451),
.B2(n_1470),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1512),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_R g1605 ( 
.A(n_1512),
.B(n_1536),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1467),
.B(n_1482),
.Y(n_1606)
);

AND2x6_ASAP7_75t_L g1607 ( 
.A(n_1512),
.B(n_1428),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1580),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1571),
.A2(n_1476),
.B(n_1528),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1601),
.B(n_1567),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1601),
.B(n_1464),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1567),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1589),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1543),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1569),
.A2(n_1447),
.B1(n_1485),
.B2(n_1494),
.C(n_1476),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1581),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1538),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1567),
.B(n_1464),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1554),
.A2(n_1434),
.B1(n_1472),
.B2(n_1494),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1594),
.B(n_1464),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1568),
.B(n_1490),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1551),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1581),
.B(n_1488),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1581),
.B(n_1488),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1594),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1551),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1568),
.B(n_1493),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1556),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1542),
.B(n_1493),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1549),
.B(n_1490),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1542),
.B(n_1469),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1578),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1607),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1582),
.B(n_1478),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1552),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1571),
.Y(n_1637)
);

NAND2xp33_ASAP7_75t_SL g1638 ( 
.A(n_1559),
.B(n_1536),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1560),
.B(n_1528),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1546),
.B(n_1472),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1553),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1597),
.B(n_1469),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1614),
.B(n_1540),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1608),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_L g1645 ( 
.A(n_1620),
.B(n_1576),
.C(n_1579),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1615),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1614),
.B(n_1583),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1616),
.A2(n_1577),
.B1(n_1574),
.B2(n_1545),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1616),
.A2(n_1577),
.B1(n_1574),
.B2(n_1545),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1611),
.B(n_1558),
.Y(n_1650)
);

OAI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1620),
.A2(n_1579),
.B1(n_1561),
.B2(n_1576),
.C(n_1556),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1606),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1609),
.B(n_1590),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1640),
.A2(n_1537),
.B1(n_1599),
.B2(n_1592),
.C(n_1575),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1638),
.B(n_1539),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1609),
.B(n_1636),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1613),
.B(n_1606),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1636),
.B(n_1564),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1638),
.B(n_1586),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1640),
.A2(n_1603),
.B1(n_1570),
.B2(n_1598),
.C(n_1562),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1613),
.B(n_1597),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1615),
.B(n_1547),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1641),
.B(n_1596),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1613),
.B(n_1597),
.Y(n_1664)
);

OAI21xp33_ASAP7_75t_L g1665 ( 
.A1(n_1635),
.A2(n_1576),
.B(n_1556),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1629),
.B(n_1556),
.C(n_1603),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1613),
.B(n_1557),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1641),
.B(n_1541),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1641),
.B(n_1618),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1618),
.B(n_1595),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_SL g1671 ( 
.A1(n_1629),
.A2(n_1559),
.B1(n_1573),
.B2(n_1591),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1629),
.B(n_1550),
.C(n_1584),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1613),
.B(n_1555),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1618),
.B(n_1595),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1675)
);

OAI21xp33_ASAP7_75t_L g1676 ( 
.A1(n_1635),
.A2(n_1573),
.B(n_1602),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1629),
.B(n_1550),
.C(n_1548),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1678)
);

NAND3xp33_ASAP7_75t_L g1679 ( 
.A(n_1629),
.B(n_1635),
.C(n_1621),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1629),
.B(n_1572),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1639),
.B(n_1548),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1627),
.B(n_1548),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1644),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1646),
.B(n_1626),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1677),
.B(n_1634),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1644),
.Y(n_1687)
);

AND2x4_ASAP7_75t_SL g1688 ( 
.A(n_1659),
.B(n_1629),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1669),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1682),
.B(n_1617),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1670),
.Y(n_1691)
);

OAI222xp33_ASAP7_75t_L g1692 ( 
.A1(n_1651),
.A2(n_1617),
.B1(n_1619),
.B2(n_1625),
.C1(n_1624),
.C2(n_1630),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1657),
.B(n_1617),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1647),
.B(n_1626),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1674),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1656),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1677),
.B(n_1634),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1679),
.B(n_1621),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1683),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1681),
.Y(n_1700)
);

NOR2x1_ASAP7_75t_L g1701 ( 
.A(n_1672),
.B(n_1634),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1668),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1653),
.B(n_1630),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1663),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1679),
.A2(n_1610),
.B(n_1625),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1672),
.B(n_1634),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1661),
.B(n_1625),
.Y(n_1707)
);

NAND2x1p5_ASAP7_75t_L g1708 ( 
.A(n_1655),
.B(n_1629),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1662),
.B(n_1621),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1645),
.A2(n_1629),
.B1(n_1593),
.B2(n_1600),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1652),
.B(n_1624),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1675),
.B(n_1631),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1661),
.B(n_1624),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1660),
.B(n_1631),
.Y(n_1714)
);

INVxp33_ASAP7_75t_SL g1715 ( 
.A(n_1710),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1686),
.B(n_1667),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1691),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1691),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1684),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1695),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1714),
.B(n_1654),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1686),
.B(n_1667),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1709),
.B(n_1658),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1695),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1686),
.B(n_1664),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1686),
.B(n_1664),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1697),
.B(n_1650),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1684),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1714),
.B(n_1643),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1684),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1687),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1687),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1697),
.B(n_1650),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_SL g1734 ( 
.A(n_1701),
.B(n_1676),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1687),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1697),
.B(n_1673),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1712),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1709),
.B(n_1680),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1697),
.B(n_1673),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1689),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1706),
.B(n_1665),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1689),
.Y(n_1742)
);

INVxp67_ASAP7_75t_SL g1743 ( 
.A(n_1701),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1706),
.B(n_1632),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1694),
.B(n_1678),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1685),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1706),
.B(n_1665),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1694),
.B(n_1666),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1706),
.B(n_1676),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1696),
.B(n_1612),
.Y(n_1750)
);

INVxp67_ASAP7_75t_SL g1751 ( 
.A(n_1708),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1696),
.B(n_1666),
.Y(n_1752)
);

NAND2xp33_ASAP7_75t_SL g1753 ( 
.A(n_1710),
.B(n_1602),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1711),
.B(n_1632),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1685),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1712),
.B(n_1633),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1721),
.A2(n_1648),
.B(n_1649),
.C(n_1700),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1727),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1729),
.B(n_1699),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1719),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1715),
.B(n_1699),
.Y(n_1761)
);

AND2x2_ASAP7_75t_SL g1762 ( 
.A(n_1734),
.B(n_1544),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1753),
.Y(n_1763)
);

OAI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1734),
.A2(n_1743),
.B1(n_1752),
.B2(n_1748),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_1749),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1736),
.B(n_1739),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1736),
.B(n_1688),
.Y(n_1767)
);

OAI211xp5_ASAP7_75t_SL g1768 ( 
.A1(n_1752),
.A2(n_1671),
.B(n_1704),
.C(n_1698),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1737),
.B(n_1704),
.Y(n_1769)
);

NOR2xp67_ASAP7_75t_L g1770 ( 
.A(n_1749),
.B(n_1698),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1740),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1740),
.Y(n_1772)
);

AOI211xp5_ASAP7_75t_L g1773 ( 
.A1(n_1741),
.A2(n_1692),
.B(n_1700),
.C(n_1702),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1746),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1741),
.B(n_1702),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1742),
.Y(n_1776)
);

OAI322xp33_ASAP7_75t_L g1777 ( 
.A1(n_1748),
.A2(n_1708),
.A3(n_1703),
.B1(n_1628),
.B2(n_1622),
.C1(n_1642),
.C2(n_1627),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1747),
.B(n_1700),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1742),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1717),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1747),
.B(n_1690),
.Y(n_1781)
);

XOR2x2_ASAP7_75t_L g1782 ( 
.A(n_1727),
.B(n_1708),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1746),
.Y(n_1783)
);

AND3x1_ASAP7_75t_SL g1784 ( 
.A(n_1755),
.B(n_1563),
.C(n_1593),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1717),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1718),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1733),
.B(n_1688),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1718),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1720),
.Y(n_1789)
);

OA222x2_ASAP7_75t_L g1790 ( 
.A1(n_1746),
.A2(n_1705),
.B1(n_1642),
.B2(n_1637),
.C1(n_1688),
.C2(n_1605),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1720),
.Y(n_1791)
);

NOR2x1_ASAP7_75t_L g1792 ( 
.A(n_1764),
.B(n_1755),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1762),
.B(n_1739),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1765),
.B(n_1733),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1774),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1757),
.B(n_1716),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1757),
.B(n_1716),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1774),
.Y(n_1798)
);

INVx2_ASAP7_75t_SL g1799 ( 
.A(n_1787),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1762),
.B(n_1725),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1783),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1783),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1781),
.B(n_1724),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1766),
.Y(n_1804)
);

NAND2x1p5_ASAP7_75t_L g1805 ( 
.A(n_1763),
.B(n_1725),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1775),
.B(n_1759),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1769),
.B(n_1724),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1758),
.Y(n_1808)
);

INVx1_ASAP7_75t_SL g1809 ( 
.A(n_1778),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1767),
.B(n_1726),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1787),
.B(n_1726),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1771),
.Y(n_1812)
);

INVxp67_ASAP7_75t_L g1813 ( 
.A(n_1761),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1772),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1768),
.B(n_1563),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1787),
.Y(n_1816)
);

NAND3xp33_ASAP7_75t_L g1817 ( 
.A(n_1792),
.B(n_1764),
.C(n_1773),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1813),
.B(n_1745),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1793),
.B(n_1722),
.Y(n_1819)
);

NOR2xp67_ASAP7_75t_L g1820 ( 
.A(n_1799),
.B(n_1770),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1811),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1809),
.B(n_1722),
.Y(n_1822)
);

AOI21xp33_ASAP7_75t_L g1823 ( 
.A1(n_1793),
.A2(n_1791),
.B(n_1776),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1801),
.Y(n_1824)
);

OAI221xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1796),
.A2(n_1751),
.B1(n_1790),
.B2(n_1788),
.C(n_1786),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1808),
.B(n_1779),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1805),
.A2(n_1744),
.B1(n_1745),
.B2(n_1723),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1797),
.A2(n_1782),
.B(n_1777),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1801),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1800),
.A2(n_1782),
.B1(n_1785),
.B2(n_1789),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1800),
.A2(n_1780),
.B1(n_1705),
.B2(n_1744),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1808),
.B(n_1738),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1811),
.B(n_1744),
.Y(n_1833)
);

AOI222xp33_ASAP7_75t_L g1834 ( 
.A1(n_1815),
.A2(n_1744),
.B1(n_1784),
.B2(n_1750),
.C1(n_1760),
.C2(n_1731),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1804),
.A2(n_1705),
.B1(n_1760),
.B2(n_1738),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1820),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1824),
.Y(n_1837)
);

INVxp67_ASAP7_75t_SL g1838 ( 
.A(n_1817),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1827),
.B(n_1805),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1830),
.A2(n_1799),
.B1(n_1816),
.B2(n_1804),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1828),
.A2(n_1805),
.B(n_1794),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1830),
.A2(n_1816),
.B1(n_1810),
.B2(n_1806),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1821),
.B(n_1810),
.Y(n_1843)
);

AOI32xp33_ASAP7_75t_L g1844 ( 
.A1(n_1819),
.A2(n_1798),
.A3(n_1802),
.B1(n_1795),
.B2(n_1814),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1829),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_SL g1846 ( 
.A(n_1825),
.B(n_1806),
.Y(n_1846)
);

OAI321xp33_ASAP7_75t_L g1847 ( 
.A1(n_1838),
.A2(n_1831),
.A3(n_1835),
.B1(n_1832),
.B2(n_1822),
.C(n_1826),
.Y(n_1847)
);

O2A1O1Ixp33_ASAP7_75t_SL g1848 ( 
.A1(n_1839),
.A2(n_1823),
.B(n_1812),
.C(n_1818),
.Y(n_1848)
);

AOI211xp5_ASAP7_75t_L g1849 ( 
.A1(n_1846),
.A2(n_1841),
.B(n_1842),
.C(n_1836),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1843),
.A2(n_1840),
.B(n_1844),
.Y(n_1850)
);

OAI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1837),
.A2(n_1834),
.B1(n_1831),
.B2(n_1835),
.C(n_1803),
.Y(n_1851)
);

AOI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1845),
.A2(n_1807),
.B1(n_1803),
.B2(n_1833),
.C(n_1731),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1843),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1838),
.A2(n_1784),
.B1(n_1807),
.B2(n_1705),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1843),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1849),
.B(n_1756),
.Y(n_1856)
);

OAI21xp33_ASAP7_75t_L g1857 ( 
.A1(n_1850),
.A2(n_1735),
.B(n_1732),
.Y(n_1857)
);

NOR3xp33_ASAP7_75t_L g1858 ( 
.A(n_1847),
.B(n_1437),
.C(n_1728),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_1851),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1853),
.Y(n_1860)
);

NOR4xp75_ASAP7_75t_L g1861 ( 
.A(n_1856),
.B(n_1848),
.C(n_1855),
.D(n_1852),
.Y(n_1861)
);

NAND4xp25_ASAP7_75t_L g1862 ( 
.A(n_1859),
.B(n_1854),
.C(n_1723),
.D(n_1735),
.Y(n_1862)
);

NOR2xp67_ASAP7_75t_L g1863 ( 
.A(n_1860),
.B(n_1857),
.Y(n_1863)
);

OA211x2_ASAP7_75t_L g1864 ( 
.A1(n_1858),
.A2(n_1499),
.B(n_1585),
.C(n_1605),
.Y(n_1864)
);

NOR2x1_ASAP7_75t_L g1865 ( 
.A(n_1860),
.B(n_1728),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1859),
.B(n_1756),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1865),
.Y(n_1867)
);

A2O1A1Ixp33_ASAP7_75t_SL g1868 ( 
.A1(n_1866),
.A2(n_1728),
.B(n_1719),
.C(n_1730),
.Y(n_1868)
);

OAI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1863),
.A2(n_1862),
.B(n_1861),
.Y(n_1869)
);

NAND3xp33_ASAP7_75t_L g1870 ( 
.A(n_1864),
.B(n_1719),
.C(n_1732),
.Y(n_1870)
);

NOR2x1_ASAP7_75t_L g1871 ( 
.A(n_1863),
.B(n_1730),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1867),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1871),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1869),
.Y(n_1874)
);

INVx1_ASAP7_75t_SL g1875 ( 
.A(n_1873),
.Y(n_1875)
);

OAI211xp5_ASAP7_75t_L g1876 ( 
.A1(n_1875),
.A2(n_1874),
.B(n_1872),
.C(n_1868),
.Y(n_1876)
);

AOI211xp5_ASAP7_75t_L g1877 ( 
.A1(n_1876),
.A2(n_1870),
.B(n_1585),
.C(n_1512),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1876),
.Y(n_1878)
);

XOR2xp5_ASAP7_75t_L g1879 ( 
.A(n_1878),
.B(n_1707),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1877),
.Y(n_1880)
);

OAI221xp5_ASAP7_75t_SL g1881 ( 
.A1(n_1879),
.A2(n_1754),
.B1(n_1693),
.B2(n_1690),
.C(n_1713),
.Y(n_1881)
);

NAND3xp33_ASAP7_75t_SL g1882 ( 
.A(n_1880),
.B(n_1588),
.C(n_1565),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1882),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1883),
.A2(n_1881),
.B1(n_1707),
.B2(n_1754),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1884),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1885),
.B(n_1707),
.Y(n_1886)
);

OAI21xp5_ASAP7_75t_SL g1887 ( 
.A1(n_1886),
.A2(n_1498),
.B(n_1707),
.Y(n_1887)
);

OAI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1887),
.A2(n_1565),
.B1(n_1604),
.B2(n_1713),
.Y(n_1888)
);

AOI211xp5_ASAP7_75t_L g1889 ( 
.A1(n_1888),
.A2(n_1497),
.B(n_1604),
.C(n_1693),
.Y(n_1889)
);


endmodule