module fake_netlist_6_659_n_1941 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1941);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1941;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1888;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_5),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_113),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_34),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_136),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_72),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_163),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_96),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_58),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_44),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_71),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_86),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_127),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_21),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_105),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_109),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_120),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_103),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_90),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_67),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_92),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_44),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_162),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_26),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_34),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_175),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_131),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_145),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_53),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_100),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_8),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_62),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_82),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_135),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_153),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_155),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_130),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_134),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_143),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_183),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_157),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_110),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_29),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_201),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_14),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_167),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_132),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_191),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_91),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_174),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_73),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_111),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_171),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_20),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_81),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_139),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_11),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_30),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_197),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_85),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_65),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_97),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_196),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_190),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_186),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_138),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_173),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_188),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_12),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_45),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_61),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_84),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_177),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_172),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_115),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_75),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_39),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_156),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_38),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_192),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_21),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_6),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_39),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_67),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_47),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_19),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_1),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_74),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_15),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_151),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_182),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_87),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_78),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_31),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_178),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_48),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_77),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_165),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_5),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_79),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_56),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_125),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_95),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_60),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_147),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_16),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_12),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_107),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_37),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_99),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_140),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_198),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_46),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_24),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_160),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_13),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_51),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_66),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_22),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_123),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_31),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_41),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_47),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_11),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_58),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_27),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_159),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_51),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_114),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_18),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_168),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_88),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_104),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_141),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_38),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_65),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_121),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_25),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_0),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_142),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_20),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_13),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_28),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_137),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_17),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_66),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_8),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_48),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_122),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_64),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_15),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_4),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_0),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_119),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_37),
.Y(n_364)
);

BUFx8_ASAP7_75t_SL g365 ( 
.A(n_41),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_146),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_53),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_158),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_118),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_176),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_27),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_161),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_106),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_2),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_133),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_7),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_148),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_69),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_56),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_22),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_24),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_35),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_7),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_16),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_35),
.Y(n_385)
);

BUFx5_ASAP7_75t_L g386 ( 
.A(n_179),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_170),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_144),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_26),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_112),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_180),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_94),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_17),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_50),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_60),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_59),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_25),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_117),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_57),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_187),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_83),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_76),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_9),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_89),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_46),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_365),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_327),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_327),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_359),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_280),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_251),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_327),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_327),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_203),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_248),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_208),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_234),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_254),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_263),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_242),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_298),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_298),
.Y(n_428)
);

INVxp33_ASAP7_75t_SL g429 ( 
.A(n_202),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_298),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_278),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_250),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_298),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_211),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_298),
.Y(n_435)
);

INVxp33_ASAP7_75t_L g436 ( 
.A(n_213),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_360),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_279),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_252),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_252),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_270),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_270),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_330),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_286),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_367),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_236),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_291),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_292),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_386),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_294),
.Y(n_450)
);

INVxp33_ASAP7_75t_SL g451 ( 
.A(n_202),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_236),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_296),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_305),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_271),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_204),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_305),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_285),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_397),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_397),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_341),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_330),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_232),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_308),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_266),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_358),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_310),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_267),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_288),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_313),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_211),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_315),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_290),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_330),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_222),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_293),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_347),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_378),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_347),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_295),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_303),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_262),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_205),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_323),
.Y(n_484)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_325),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_335),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_386),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_345),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_253),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_350),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_351),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_316),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_355),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_357),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_361),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_371),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_318),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_322),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_326),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_367),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_374),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_256),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_260),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_376),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_382),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_284),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_328),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_386),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_331),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_418),
.B(n_423),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_506),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_421),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_427),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_489),
.Y(n_517)
);

INVx6_ASAP7_75t_L g518 ( 
.A(n_506),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_483),
.B(n_235),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_506),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_434),
.B(n_235),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_506),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_428),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_422),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_428),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_430),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_502),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_430),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_434),
.B(n_261),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_506),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_433),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_471),
.B(n_261),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_413),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_503),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_471),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_433),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_409),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_412),
.A2(n_354),
.B1(n_364),
.B2(n_238),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_410),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_414),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_435),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_435),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_446),
.B(n_389),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_415),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_437),
.B(n_246),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_406),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_407),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_406),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_408),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_416),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_426),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_432),
.B(n_246),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_456),
.B(n_247),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_408),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_501),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_501),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_437),
.B(n_247),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_407),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_452),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_454),
.B(n_207),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_449),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_412),
.A2(n_394),
.B1(n_403),
.B2(n_206),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_449),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_459),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_487),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_457),
.B(n_389),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_504),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_487),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_460),
.B(n_384),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_508),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_508),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_413),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_504),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_439),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_505),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_439),
.A2(n_281),
.B(n_258),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_475),
.B(n_249),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_440),
.B(n_258),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_505),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_440),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_420),
.B(n_281),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_441),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_459),
.B(n_317),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_441),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_442),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_455),
.B(n_206),
.Y(n_586)
);

XNOR2x2_ASAP7_75t_L g587 ( 
.A(n_463),
.B(n_332),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_442),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_482),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_514),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_564),
.B(n_411),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_577),
.B(n_589),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_581),
.B(n_317),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_546),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_535),
.B(n_419),
.Y(n_596)
);

AND3x2_ASAP7_75t_L g597 ( 
.A(n_533),
.B(n_399),
.C(n_395),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_586),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_517),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_547),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_513),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_535),
.B(n_424),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_546),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_511),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_524),
.B(n_458),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_548),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_511),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_511),
.Y(n_608)
);

INVx6_ASAP7_75t_L g609 ( 
.A(n_550),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_548),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_512),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_553),
.B(n_284),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_512),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_L g614 ( 
.A(n_519),
.B(n_284),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_512),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_560),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_549),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_552),
.B(n_398),
.Y(n_618)
);

NOR2x1p5_ASAP7_75t_L g619 ( 
.A(n_558),
.B(n_482),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_560),
.B(n_284),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_527),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_561),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_534),
.Y(n_623)
);

AND2x2_ASAP7_75t_SL g624 ( 
.A(n_533),
.B(n_284),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_561),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_561),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_549),
.B(n_424),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_554),
.B(n_425),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_554),
.B(n_212),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_521),
.B(n_429),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_537),
.B(n_425),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_571),
.Y(n_632)
);

INVx8_ASAP7_75t_L g633 ( 
.A(n_510),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_563),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_513),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g636 ( 
.A(n_538),
.B(n_462),
.C(n_443),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_587),
.A2(n_477),
.B1(n_466),
.B2(n_461),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_583),
.B(n_385),
.Y(n_638)
);

CKINVDCx6p67_ASAP7_75t_R g639 ( 
.A(n_551),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_529),
.B(n_431),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_L g641 ( 
.A1(n_562),
.A2(n_396),
.B1(n_337),
.B2(n_334),
.Y(n_641)
);

BUFx10_ASAP7_75t_L g642 ( 
.A(n_572),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_586),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_532),
.B(n_451),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_562),
.B(n_438),
.C(n_431),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_559),
.Y(n_646)
);

NOR2x1p5_ASAP7_75t_L g647 ( 
.A(n_559),
.B(n_438),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_559),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_538),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_543),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_537),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_543),
.Y(n_652)
);

BUFx4f_ASAP7_75t_L g653 ( 
.A(n_550),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_537),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_571),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_563),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_539),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_539),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_566),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_566),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_539),
.B(n_444),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_569),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_563),
.Y(n_663)
);

NOR3xp33_ASAP7_75t_L g664 ( 
.A(n_569),
.B(n_479),
.C(n_474),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_540),
.B(n_447),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_510),
.Y(n_666)
);

AO21x2_ASAP7_75t_L g667 ( 
.A1(n_576),
.A2(n_221),
.B(n_217),
.Y(n_667)
);

XNOR2xp5_ASAP7_75t_L g668 ( 
.A(n_510),
.B(n_478),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_513),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_510),
.B(n_465),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_540),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_571),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_540),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_544),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_545),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_555),
.B(n_447),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_555),
.B(n_448),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_544),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_545),
.B(n_223),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_513),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_513),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_545),
.A2(n_494),
.B1(n_468),
.B2(n_469),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_545),
.B(n_473),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_580),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_550),
.B(n_448),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_557),
.A2(n_488),
.B1(n_496),
.B2(n_495),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_513),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_580),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_550),
.B(n_386),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_580),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_557),
.B(n_450),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_550),
.B(n_450),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_556),
.B(n_453),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_580),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_520),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_557),
.A2(n_492),
.B1(n_507),
.B2(n_499),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_550),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_557),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_518),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_578),
.B(n_453),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_556),
.B(n_464),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_563),
.B(n_464),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_567),
.Y(n_703)
);

INVx6_ASAP7_75t_L g704 ( 
.A(n_580),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_578),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_580),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_563),
.B(n_467),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_520),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_578),
.B(n_476),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_563),
.B(n_467),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_520),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_578),
.A2(n_497),
.B1(n_507),
.B2(n_499),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_520),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_584),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_565),
.B(n_470),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_520),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_584),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_573),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_575),
.B(n_470),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_520),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_584),
.B(n_472),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_584),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_584),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_575),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_579),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_584),
.Y(n_726)
);

BUFx6f_ASAP7_75t_SL g727 ( 
.A(n_579),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_574),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_515),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_515),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_576),
.B(n_480),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_516),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_516),
.Y(n_733)
);

AND2x2_ASAP7_75t_SL g734 ( 
.A(n_582),
.B(n_225),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_582),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_624),
.B(n_565),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_624),
.B(n_472),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_698),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_683),
.B(n_481),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_683),
.B(n_484),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_735),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_734),
.A2(n_386),
.B1(n_392),
.B2(n_391),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_616),
.B(n_565),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_616),
.B(n_593),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_650),
.B(n_492),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_604),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_734),
.B(n_565),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_703),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_628),
.B(n_497),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_591),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_728),
.B(n_565),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_650),
.A2(n_302),
.B1(n_309),
.B2(n_275),
.Y(n_752)
);

NAND2x1_ASAP7_75t_L g753 ( 
.A(n_609),
.B(n_518),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_728),
.B(n_565),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_683),
.B(n_486),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_718),
.B(n_498),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_604),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_627),
.B(n_498),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_633),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_675),
.A2(n_509),
.B1(n_274),
.B2(n_320),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_595),
.B(n_603),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_606),
.B(n_568),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_610),
.B(n_568),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_607),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_617),
.B(n_568),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_633),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_709),
.B(n_490),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_652),
.A2(n_300),
.B1(n_299),
.B2(n_277),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_627),
.B(n_436),
.Y(n_769)
);

NAND2x1p5_ASAP7_75t_L g770 ( 
.A(n_666),
.B(n_228),
.Y(n_770)
);

NAND2x1_ASAP7_75t_L g771 ( 
.A(n_609),
.B(n_518),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_652),
.B(n_568),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_675),
.A2(n_265),
.B1(n_264),
.B2(n_268),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_659),
.B(n_568),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_602),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_647),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_659),
.A2(n_259),
.B1(n_272),
.B2(n_257),
.Y(n_777)
);

BUFx5_ASAP7_75t_L g778 ( 
.A(n_679),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_660),
.B(n_207),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_660),
.B(n_209),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_705),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_631),
.B(n_485),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_719),
.B(n_630),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_591),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_731),
.A2(n_386),
.B1(n_368),
.B2(n_241),
.Y(n_785)
);

BUFx6f_ASAP7_75t_SL g786 ( 
.A(n_600),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_644),
.B(n_568),
.Y(n_787)
);

BUFx6f_ASAP7_75t_SL g788 ( 
.A(n_600),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_661),
.B(n_209),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_607),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_691),
.A2(n_269),
.B1(n_273),
.B2(n_276),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_724),
.B(n_570),
.Y(n_792)
);

NAND2x1p5_ASAP7_75t_L g793 ( 
.A(n_699),
.B(n_237),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_662),
.B(n_347),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_702),
.B(n_570),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_691),
.A2(n_282),
.B1(n_283),
.B2(n_287),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_679),
.B(n_386),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_665),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_608),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_700),
.A2(n_289),
.B1(n_297),
.B2(n_301),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_608),
.Y(n_801)
);

OR2x6_ASAP7_75t_L g802 ( 
.A(n_638),
.B(n_491),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_611),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_705),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_611),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_731),
.A2(n_386),
.B1(n_369),
.B2(n_329),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_646),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_648),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_709),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_707),
.B(n_570),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_676),
.B(n_493),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_710),
.B(n_570),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_677),
.B(n_210),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_715),
.B(n_523),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_693),
.B(n_210),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_685),
.B(n_523),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_709),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_633),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_613),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_701),
.B(n_445),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_692),
.B(n_525),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_729),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_664),
.B(n_500),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_594),
.B(n_526),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_696),
.B(n_215),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_613),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_729),
.B(n_526),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_730),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_730),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_712),
.B(n_215),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_592),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_732),
.B(n_733),
.Y(n_832)
);

O2A1O1Ixp5_ASAP7_75t_L g833 ( 
.A1(n_618),
.A2(n_528),
.B(n_531),
.C(n_542),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_638),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_705),
.B(n_255),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_732),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_733),
.B(n_620),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_640),
.B(n_700),
.Y(n_838)
);

OR2x6_ASAP7_75t_L g839 ( 
.A(n_638),
.B(n_338),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_R g840 ( 
.A(n_649),
.B(n_214),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_721),
.B(n_353),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_731),
.A2(n_372),
.B1(n_390),
.B2(n_401),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_731),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_670),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_721),
.B(n_363),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_615),
.Y(n_846)
);

BUFx6f_ASAP7_75t_SL g847 ( 
.A(n_600),
.Y(n_847)
);

AND2x4_ASAP7_75t_SL g848 ( 
.A(n_639),
.B(n_388),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_SL g849 ( 
.A(n_601),
.B(n_530),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_670),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_620),
.B(n_528),
.Y(n_851)
);

BUFx8_ASAP7_75t_L g852 ( 
.A(n_598),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_618),
.B(n_531),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_670),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_640),
.B(n_645),
.Y(n_855)
);

OAI221xp5_ASAP7_75t_L g856 ( 
.A1(n_682),
.A2(n_686),
.B1(n_638),
.B2(n_670),
.C(n_637),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_697),
.B(n_536),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_596),
.B(n_216),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_684),
.B(n_404),
.Y(n_859)
);

OAI22xp33_ASAP7_75t_L g860 ( 
.A1(n_649),
.A2(n_348),
.B1(n_219),
.B2(n_227),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_674),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_651),
.B(n_536),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_639),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_654),
.B(n_541),
.Y(n_864)
);

NAND2x1_ASAP7_75t_L g865 ( 
.A(n_609),
.B(n_518),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_657),
.B(n_541),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_725),
.B(n_216),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_668),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_684),
.B(n_304),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_688),
.B(n_690),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_688),
.B(n_306),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_641),
.B(n_218),
.Y(n_872)
);

BUFx8_ASAP7_75t_L g873 ( 
.A(n_727),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_658),
.B(n_542),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_671),
.B(n_574),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_629),
.A2(n_574),
.B1(n_588),
.B2(n_214),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_642),
.B(n_220),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_727),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_599),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_622),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_622),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_690),
.B(n_307),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_673),
.B(n_574),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_599),
.Y(n_884)
);

BUFx6f_ASAP7_75t_SL g885 ( 
.A(n_642),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_625),
.Y(n_886)
);

AND2x2_ASAP7_75t_SL g887 ( 
.A(n_636),
.B(n_585),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_678),
.B(n_588),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_634),
.B(n_588),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_642),
.B(n_500),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_633),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_626),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_744),
.B(n_626),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_844),
.B(n_619),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_850),
.B(n_699),
.Y(n_895)
);

BUFx12f_ASAP7_75t_L g896 ( 
.A(n_873),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_822),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_838),
.A2(n_727),
.B1(n_679),
.B2(n_629),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_744),
.B(n_813),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_813),
.B(n_632),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_838),
.B(n_653),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_811),
.B(n_621),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_742),
.A2(n_629),
.B1(n_612),
.B2(n_614),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_828),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_829),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_759),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_736),
.A2(n_612),
.B(n_614),
.C(n_689),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_836),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_855),
.A2(n_679),
.B1(n_629),
.B2(n_722),
.Y(n_909)
);

AOI21xp33_ASAP7_75t_L g910 ( 
.A1(n_758),
.A2(n_623),
.B(n_621),
.Y(n_910)
);

AND2x2_ASAP7_75t_SL g911 ( 
.A(n_742),
.B(n_842),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_746),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_753),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_757),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_782),
.B(n_655),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_771),
.Y(n_916)
);

AND3x1_ASAP7_75t_L g917 ( 
.A(n_872),
.B(n_597),
.C(n_643),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_842),
.A2(n_629),
.B1(n_667),
.B2(n_679),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_759),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_750),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_832),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_748),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_798),
.B(n_623),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_820),
.B(n_655),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_865),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_749),
.B(n_605),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_795),
.A2(n_812),
.B(n_810),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_764),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_R g929 ( 
.A(n_879),
.B(n_220),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_790),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_781),
.Y(n_931)
);

AND2x6_ASAP7_75t_SL g932 ( 
.A(n_872),
.B(n_219),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_785),
.A2(n_629),
.B1(n_667),
.B2(n_679),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_781),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_855),
.B(n_653),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_789),
.B(n_672),
.Y(n_936)
);

NOR3xp33_ASAP7_75t_SL g937 ( 
.A(n_840),
.B(n_229),
.C(n_227),
.Y(n_937)
);

INVxp33_ASAP7_75t_L g938 ( 
.A(n_756),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_769),
.B(n_339),
.C(n_333),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_843),
.B(n_653),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_759),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_785),
.A2(n_672),
.B1(n_229),
.B2(n_393),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_745),
.B(n_231),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_SL g944 ( 
.A1(n_868),
.A2(n_231),
.B1(n_239),
.B2(n_344),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_799),
.Y(n_945)
);

BUFx4f_ASAP7_75t_L g946 ( 
.A(n_887),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_807),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_786),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_801),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_803),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_854),
.B(n_694),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_808),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_778),
.B(n_694),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_805),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_809),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_819),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_826),
.Y(n_957)
);

BUFx12f_ASAP7_75t_SL g958 ( 
.A(n_802),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_890),
.B(n_239),
.Y(n_959)
);

OAI22xp33_ASAP7_75t_L g960 ( 
.A1(n_856),
.A2(n_352),
.B1(n_344),
.B2(n_380),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_787),
.B(n_635),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_759),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_817),
.B(n_706),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_774),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_739),
.B(n_706),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_766),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_846),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_775),
.B(n_224),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_804),
.Y(n_969)
);

INVxp67_ASAP7_75t_L g970 ( 
.A(n_794),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_766),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_784),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_886),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_884),
.Y(n_974)
);

INVx8_ASAP7_75t_L g975 ( 
.A(n_786),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_831),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_SL g977 ( 
.A(n_758),
.B(n_240),
.C(n_224),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_749),
.B(n_634),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_738),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_892),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_741),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_761),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_880),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_816),
.B(n_635),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_823),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_887),
.A2(n_726),
.B1(n_723),
.B2(n_722),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_827),
.Y(n_987)
);

AND2x6_ASAP7_75t_L g988 ( 
.A(n_766),
.B(n_714),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_821),
.B(n_669),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_769),
.B(n_868),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_766),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_861),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_834),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_834),
.Y(n_994)
);

NAND3xp33_ASAP7_75t_SL g995 ( 
.A(n_858),
.B(n_240),
.C(n_230),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_861),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_739),
.Y(n_997)
);

OR2x6_ASAP7_75t_L g998 ( 
.A(n_863),
.B(n_802),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_783),
.A2(n_726),
.B1(n_723),
.B2(n_714),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_858),
.A2(n_717),
.B(n_689),
.C(n_588),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_743),
.B(n_669),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_818),
.B(n_634),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_778),
.B(n_717),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_778),
.B(n_656),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_814),
.B(n_881),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_788),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_740),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_SL g1008 ( 
.A1(n_873),
.A2(n_403),
.B1(n_393),
.B2(n_383),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_740),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_737),
.B(n_656),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_755),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_755),
.B(n_656),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_818),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_776),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_767),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_767),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_751),
.B(n_681),
.Y(n_1017)
);

NAND2xp33_ASAP7_75t_SL g1018 ( 
.A(n_788),
.B(n_226),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_754),
.B(n_681),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_841),
.B(n_681),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_857),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_862),
.Y(n_1022)
);

AND2x4_ASAP7_75t_SL g1023 ( 
.A(n_878),
.B(n_663),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_864),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_SL g1025 ( 
.A1(n_839),
.A2(n_362),
.B1(n_383),
.B2(n_381),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_870),
.Y(n_1026)
);

AND2x6_ASAP7_75t_L g1027 ( 
.A(n_818),
.B(n_695),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_802),
.B(n_663),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_SL g1029 ( 
.A1(n_839),
.A2(n_381),
.B1(n_380),
.B2(n_379),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_841),
.B(n_695),
.Y(n_1030)
);

NOR2xp67_ASAP7_75t_L g1031 ( 
.A(n_760),
.B(n_311),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_847),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_770),
.B(n_818),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_845),
.B(n_720),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_839),
.B(n_663),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_770),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_793),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_778),
.B(n_601),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_778),
.B(n_601),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_866),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_874),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_833),
.A2(n_720),
.B(n_716),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_778),
.B(n_601),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_845),
.B(n_695),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_876),
.B(n_680),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_779),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_876),
.B(n_680),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_SL g1048 ( 
.A1(n_878),
.A2(n_379),
.B1(n_362),
.B2(n_356),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_772),
.B(n_806),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_815),
.B(n_405),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_747),
.A2(n_704),
.B1(n_716),
.B2(n_713),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_762),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_747),
.A2(n_835),
.B1(n_869),
.B2(n_871),
.Y(n_1053)
);

NOR2xp67_ASAP7_75t_L g1054 ( 
.A(n_791),
.B(n_796),
.Y(n_1054)
);

NOR2x1p5_ASAP7_75t_L g1055 ( 
.A(n_847),
.B(n_352),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_891),
.B(n_713),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_833),
.A2(n_716),
.B(n_713),
.C(n_366),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_870),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_835),
.A2(n_869),
.B1(n_871),
.B2(n_882),
.Y(n_1059)
);

NOR2xp67_ASAP7_75t_L g1060 ( 
.A(n_800),
.B(n_312),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_736),
.A2(n_356),
.B1(n_585),
.B2(n_590),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_773),
.B(n_226),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_772),
.B(n_680),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_825),
.B(n_233),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_891),
.B(n_585),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_793),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_763),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_899),
.B(n_792),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_902),
.B(n_752),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_922),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_997),
.B(n_848),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_982),
.B(n_780),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_983),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_990),
.B(n_867),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_R g1075 ( 
.A(n_948),
.B(n_840),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_927),
.A2(n_889),
.B(n_837),
.Y(n_1076)
);

NOR2xp67_ASAP7_75t_L g1077 ( 
.A(n_970),
.B(n_877),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_911),
.A2(n_903),
.B1(n_1049),
.B2(n_946),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1022),
.B(n_824),
.Y(n_1079)
);

CKINVDCx8_ASAP7_75t_R g1080 ( 
.A(n_975),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_927),
.A2(n_797),
.B(n_765),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_960),
.A2(n_830),
.B(n_768),
.C(n_777),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_972),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_960),
.A2(n_860),
.B(n_859),
.C(n_882),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1045),
.A2(n_853),
.B(n_851),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_977),
.A2(n_860),
.B(n_859),
.C(n_883),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1045),
.A2(n_888),
.B(n_875),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1047),
.A2(n_680),
.B(n_711),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_963),
.Y(n_1089)
);

BUFx12f_ASAP7_75t_L g1090 ( 
.A(n_896),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_974),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_977),
.A2(n_590),
.B(n_522),
.C(n_885),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_SL g1093 ( 
.A1(n_935),
.A2(n_590),
.B(n_522),
.C(n_849),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1047),
.A2(n_711),
.B(n_708),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_924),
.A2(n_711),
.B(n_708),
.Y(n_1095)
);

AND2x6_ASAP7_75t_L g1096 ( 
.A(n_898),
.B(n_906),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1024),
.B(n_243),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1011),
.B(n_687),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1040),
.B(n_243),
.Y(n_1099)
);

OR2x6_ASAP7_75t_L g1100 ( 
.A(n_975),
.B(n_885),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_911),
.A2(n_244),
.B1(n_245),
.B2(n_402),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1041),
.B(n_244),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_987),
.B(n_245),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1021),
.B(n_342),
.Y(n_1104)
);

BUFx4f_ASAP7_75t_L g1105 ( 
.A(n_975),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_978),
.B(n_342),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_SL g1107 ( 
.A(n_1048),
.B(n_349),
.C(n_402),
.Y(n_1107)
);

INVxp33_ASAP7_75t_SL g1108 ( 
.A(n_926),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_985),
.A2(n_314),
.B1(n_319),
.B2(n_321),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_901),
.A2(n_935),
.B(n_1017),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_L g1111 ( 
.A(n_910),
.B(n_926),
.C(n_923),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_941),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_906),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_903),
.A2(n_377),
.B1(n_400),
.B2(n_387),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_923),
.B(n_852),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_901),
.A2(n_711),
.B(n_708),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_963),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_978),
.B(n_343),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_SL g1119 ( 
.A(n_1064),
.B(n_370),
.C(n_387),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1019),
.A2(n_708),
.B(n_687),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_921),
.B(n_992),
.Y(n_1121)
);

INVx5_ASAP7_75t_L g1122 ( 
.A(n_906),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_996),
.B(n_343),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_SL g1124 ( 
.A1(n_1050),
.A2(n_370),
.B1(n_400),
.B2(n_377),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_970),
.B(n_324),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1006),
.Y(n_1126)
);

NAND3xp33_ASAP7_75t_SL g1127 ( 
.A(n_1064),
.B(n_346),
.C(n_349),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_938),
.B(n_346),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_976),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_897),
.Y(n_1130)
);

NOR3xp33_ASAP7_75t_L g1131 ( 
.A(n_1050),
.B(n_373),
.C(n_375),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_SL g1132 ( 
.A1(n_1010),
.A2(n_522),
.B(n_704),
.C(n_336),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_946),
.A2(n_373),
.B1(n_375),
.B2(n_340),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1036),
.B(n_687),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_920),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_1032),
.Y(n_1136)
);

O2A1O1Ixp5_ASAP7_75t_SL g1137 ( 
.A1(n_940),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_915),
.B(n_3),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_995),
.A2(n_4),
.B(n_6),
.C(n_9),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1036),
.B(n_530),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_998),
.B(n_518),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1012),
.B(n_530),
.Y(n_1142)
);

OR2x6_ASAP7_75t_L g1143 ( 
.A(n_998),
.B(n_1028),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1012),
.B(n_530),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1046),
.B(n_10),
.Y(n_1145)
);

OA22x2_ASAP7_75t_L g1146 ( 
.A1(n_944),
.A2(n_993),
.B1(n_994),
.B2(n_981),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_912),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_918),
.A2(n_10),
.B1(n_14),
.B2(n_18),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_906),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1007),
.B(n_530),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1038),
.A2(n_93),
.B(n_199),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_979),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_995),
.A2(n_19),
.B(n_23),
.C(n_28),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1046),
.B(n_23),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1039),
.A2(n_98),
.B(n_193),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1054),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1057),
.A2(n_101),
.B(n_189),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_964),
.B(n_32),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_919),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1039),
.A2(n_1043),
.B(n_1004),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_998),
.B(n_70),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1015),
.B(n_108),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_993),
.A2(n_33),
.B(n_36),
.C(n_40),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1043),
.A2(n_200),
.B(n_185),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_979),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_914),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1028),
.B(n_181),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_959),
.B(n_36),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_918),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1055),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_893),
.B(n_42),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1052),
.B(n_43),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1014),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_928),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_929),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1004),
.A2(n_961),
.B(n_941),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_941),
.B(n_68),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_894),
.B(n_149),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_941),
.A2(n_169),
.B(n_166),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_994),
.A2(n_45),
.B(n_49),
.C(n_50),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_919),
.Y(n_1181)
);

BUFx10_ASAP7_75t_L g1182 ( 
.A(n_894),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_955),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1062),
.A2(n_52),
.B(n_54),
.C(n_55),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_939),
.A2(n_126),
.B1(n_152),
.B2(n_150),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_933),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_981),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_933),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_943),
.B(n_63),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1009),
.B(n_116),
.Y(n_1190)
);

AND2x2_ASAP7_75t_SL g1191 ( 
.A(n_917),
.B(n_128),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_930),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_919),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_958),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_929),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1016),
.B(n_129),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_965),
.B(n_1066),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1053),
.A2(n_1059),
.B(n_1010),
.C(n_907),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1067),
.B(n_900),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_945),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_947),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_949),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_968),
.B(n_952),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_965),
.B(n_1066),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1066),
.B(n_1035),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_936),
.B(n_904),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_905),
.B(n_908),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1066),
.B(n_1035),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1033),
.B(n_1025),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_937),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_984),
.A2(n_989),
.B(n_1002),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1061),
.A2(n_1025),
.B1(n_1029),
.B2(n_942),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_950),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1000),
.A2(n_937),
.B(n_907),
.C(n_973),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_895),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_954),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_895),
.B(n_951),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_1129),
.Y(n_1218)
);

CKINVDCx11_ASAP7_75t_R g1219 ( 
.A(n_1090),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1198),
.A2(n_1003),
.B(n_953),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1143),
.B(n_1023),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1078),
.A2(n_1001),
.A3(n_1063),
.B(n_1034),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1110),
.A2(n_1042),
.B(n_986),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1199),
.B(n_1026),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1078),
.A2(n_971),
.B(n_962),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1143),
.B(n_951),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1082),
.A2(n_1060),
.B(n_1031),
.C(n_909),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1126),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1108),
.B(n_932),
.Y(n_1229)
);

INVxp67_ASAP7_75t_SL g1230 ( 
.A(n_1152),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1070),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1081),
.A2(n_1065),
.B(n_1044),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1111),
.B(n_1029),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1074),
.B(n_1008),
.Y(n_1234)
);

NAND2x1p5_ASAP7_75t_L g1235 ( 
.A(n_1122),
.B(n_971),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1076),
.A2(n_962),
.B(n_991),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1214),
.A2(n_999),
.B(n_1030),
.Y(n_1237)
);

AOI21xp33_ASAP7_75t_L g1238 ( 
.A1(n_1212),
.A2(n_1020),
.B(n_1037),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1068),
.B(n_1058),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1079),
.B(n_1206),
.Y(n_1240)
);

OAI22x1_ASAP7_75t_L g1241 ( 
.A1(n_1209),
.A2(n_1008),
.B1(n_969),
.B2(n_931),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1121),
.B(n_969),
.Y(n_1242)
);

INVxp67_ASAP7_75t_SL g1243 ( 
.A(n_1165),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_SL g1244 ( 
.A1(n_1186),
.A2(n_1051),
.B(n_967),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1116),
.A2(n_934),
.B(n_916),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1189),
.B(n_942),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1215),
.B(n_956),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1085),
.A2(n_1087),
.B(n_1211),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1091),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_SL g1250 ( 
.A1(n_1186),
.A2(n_980),
.B(n_957),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1212),
.A2(n_1037),
.B1(n_919),
.B2(n_991),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1187),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1083),
.Y(n_1253)
);

INVx5_ASAP7_75t_L g1254 ( 
.A(n_1112),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1136),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1160),
.A2(n_991),
.B(n_1013),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1188),
.A2(n_1148),
.A3(n_1169),
.B(n_1176),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1157),
.A2(n_988),
.B(n_1027),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1120),
.A2(n_913),
.B(n_925),
.Y(n_1259)
);

OAI21xp33_ASAP7_75t_L g1260 ( 
.A1(n_1124),
.A2(n_962),
.B(n_966),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1188),
.A2(n_988),
.A3(n_1027),
.B(n_913),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1084),
.A2(n_1086),
.B(n_1131),
.C(n_1203),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1095),
.A2(n_988),
.B(n_1027),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1201),
.Y(n_1264)
);

AOI21x1_ASAP7_75t_SL g1265 ( 
.A1(n_1106),
.A2(n_1056),
.B(n_1018),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1207),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1135),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1075),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1148),
.A2(n_1169),
.A3(n_1138),
.B(n_1171),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1217),
.Y(n_1270)
);

NOR3xp33_ASAP7_75t_L g1271 ( 
.A(n_1119),
.B(n_1056),
.C(n_1013),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1205),
.A2(n_1013),
.B(n_1208),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1073),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1118),
.A2(n_1112),
.B(n_1072),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1191),
.B(n_1145),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1151),
.A2(n_1155),
.B(n_1164),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1137),
.A2(n_1172),
.B(n_1069),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_L g1278 ( 
.A(n_1128),
.B(n_1156),
.C(n_1153),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1077),
.B(n_1115),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1179),
.A2(n_1150),
.B(n_1092),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1089),
.B(n_1117),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1127),
.A2(n_1184),
.B(n_1154),
.C(n_1168),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1197),
.A2(n_1204),
.B(n_1132),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1122),
.A2(n_1144),
.B(n_1142),
.Y(n_1284)
);

INVxp67_ASAP7_75t_SL g1285 ( 
.A(n_1113),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1196),
.A2(n_1139),
.B(n_1158),
.C(n_1103),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1122),
.A2(n_1093),
.B(n_1167),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1096),
.A2(n_1185),
.B(n_1146),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_SL g1289 ( 
.A1(n_1177),
.A2(n_1143),
.B(n_1161),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1122),
.A2(n_1162),
.B(n_1140),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1097),
.B(n_1104),
.Y(n_1291)
);

NOR2xp67_ASAP7_75t_L g1292 ( 
.A(n_1099),
.B(n_1102),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1130),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1096),
.A2(n_1146),
.B(n_1216),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1173),
.Y(n_1295)
);

NOR2xp67_ASAP7_75t_L g1296 ( 
.A(n_1175),
.B(n_1213),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1080),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1147),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1194),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1166),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_1113),
.Y(n_1301)
);

INVx4_ASAP7_75t_L g1302 ( 
.A(n_1113),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1174),
.B(n_1202),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1114),
.A2(n_1183),
.B1(n_1101),
.B2(n_1161),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1210),
.B(n_1195),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1163),
.A2(n_1180),
.B(n_1190),
.C(n_1125),
.Y(n_1306)
);

AO21x1_ASAP7_75t_L g1307 ( 
.A1(n_1101),
.A2(n_1114),
.B(n_1134),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1195),
.A2(n_1071),
.B1(n_1178),
.B2(n_1109),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1192),
.A2(n_1200),
.A3(n_1123),
.B(n_1096),
.Y(n_1309)
);

AND2x2_ASAP7_75t_SL g1310 ( 
.A(n_1105),
.B(n_1178),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1096),
.A2(n_1133),
.B(n_1098),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_SL g1312 ( 
.A(n_1107),
.B(n_1161),
.C(n_1182),
.Y(n_1312)
);

AOI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1098),
.A2(n_1141),
.B(n_1071),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1149),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1182),
.B(n_1105),
.Y(n_1315)
);

BUFx8_ASAP7_75t_L g1316 ( 
.A(n_1170),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1141),
.B(n_1100),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1159),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1149),
.A2(n_1181),
.B(n_1141),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1193),
.B(n_1181),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1181),
.A2(n_1198),
.B(n_1110),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1198),
.A2(n_1005),
.B(n_1081),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1113),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1198),
.A2(n_1005),
.B(n_1081),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1199),
.B(n_899),
.Y(n_1325)
);

O2A1O1Ixp5_ASAP7_75t_L g1326 ( 
.A1(n_1198),
.A2(n_813),
.B(n_899),
.C(n_1212),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1083),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1198),
.A2(n_1110),
.B(n_1157),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1088),
.A2(n_1094),
.B(n_1116),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1199),
.B(n_899),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1199),
.B(n_899),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1198),
.A2(n_1081),
.B(n_1005),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1070),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_SL g1334 ( 
.A(n_1212),
.B(n_911),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1082),
.A2(n_855),
.B(n_838),
.C(n_1198),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1198),
.A2(n_1110),
.B(n_1078),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1083),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1198),
.A2(n_1005),
.B(n_1081),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1198),
.A2(n_1078),
.A3(n_1057),
.B(n_1110),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1143),
.B(n_975),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1129),
.Y(n_1341)
);

O2A1O1Ixp5_ASAP7_75t_SL g1342 ( 
.A1(n_1148),
.A2(n_1169),
.B(n_1188),
.C(n_1186),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1198),
.A2(n_1078),
.A3(n_1057),
.B(n_1110),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1074),
.B(n_902),
.Y(n_1344)
);

INVx1_ASAP7_75t_SL g1345 ( 
.A(n_1129),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1143),
.B(n_1215),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1113),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1129),
.B(n_990),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1082),
.A2(n_855),
.B(n_838),
.C(n_1198),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1108),
.B(n_421),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1070),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_R g1352 ( 
.A(n_1083),
.B(n_879),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1199),
.B(n_899),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1173),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1199),
.B(n_899),
.Y(n_1355)
);

O2A1O1Ixp5_ASAP7_75t_L g1356 ( 
.A1(n_1198),
.A2(n_813),
.B(n_899),
.C(n_1212),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1199),
.B(n_899),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1111),
.B(n_902),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1091),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1088),
.A2(n_1094),
.B(n_1116),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1082),
.A2(n_855),
.B(n_838),
.C(n_1198),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1088),
.A2(n_1094),
.B(n_1116),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1325),
.B(n_1330),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1219),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1234),
.B(n_1233),
.Y(n_1365)
);

NOR2x1_ASAP7_75t_L g1366 ( 
.A(n_1240),
.B(n_1296),
.Y(n_1366)
);

OR2x6_ASAP7_75t_L g1367 ( 
.A(n_1289),
.B(n_1225),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_1255),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1218),
.Y(n_1369)
);

AOI221xp5_ASAP7_75t_L g1370 ( 
.A1(n_1304),
.A2(n_1356),
.B1(n_1326),
.B2(n_1334),
.C(n_1278),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1348),
.B(n_1270),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1334),
.A2(n_1304),
.B1(n_1331),
.B2(n_1325),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1359),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1344),
.B(n_1275),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1232),
.A2(n_1259),
.B(n_1329),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1330),
.A2(n_1353),
.B1(n_1355),
.B2(n_1357),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1254),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1221),
.B(n_1340),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_1352),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1270),
.B(n_1218),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1262),
.A2(n_1286),
.B(n_1361),
.C(n_1335),
.Y(n_1381)
);

NOR2xp67_ASAP7_75t_L g1382 ( 
.A(n_1228),
.B(n_1267),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1349),
.A2(n_1227),
.B(n_1258),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1268),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1322),
.A2(n_1338),
.B(n_1324),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1360),
.A2(n_1362),
.B(n_1245),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1307),
.A2(n_1241),
.A3(n_1220),
.B(n_1251),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1345),
.B(n_1341),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1220),
.A2(n_1251),
.A3(n_1283),
.B(n_1256),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1248),
.A2(n_1258),
.B(n_1328),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1263),
.A2(n_1236),
.B(n_1321),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1336),
.A2(n_1321),
.B(n_1277),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1277),
.A2(n_1237),
.B(n_1238),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1246),
.A2(n_1358),
.B1(n_1288),
.B2(n_1355),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_SL g1395 ( 
.A1(n_1282),
.A2(n_1306),
.B(n_1353),
.C(n_1331),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1276),
.A2(n_1265),
.B(n_1280),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1298),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1292),
.B(n_1288),
.C(n_1291),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1357),
.B(n_1345),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1314),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1302),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1300),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1346),
.B(n_1317),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1354),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1237),
.A2(n_1238),
.B(n_1244),
.Y(n_1405)
);

AO21x2_ASAP7_75t_L g1406 ( 
.A1(n_1287),
.A2(n_1311),
.B(n_1294),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1274),
.A2(n_1223),
.B(n_1313),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1254),
.B(n_1310),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1247),
.B(n_1305),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1346),
.B(n_1308),
.Y(n_1410)
);

A2O1A1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1260),
.A2(n_1240),
.B(n_1311),
.C(n_1266),
.Y(n_1411)
);

NAND2x1_ASAP7_75t_L g1412 ( 
.A(n_1319),
.B(n_1250),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1279),
.A2(n_1312),
.B1(n_1271),
.B2(n_1229),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1223),
.A2(n_1272),
.B(n_1290),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1242),
.A2(n_1239),
.B(n_1224),
.Y(n_1415)
);

AND2x2_ASAP7_75t_SL g1416 ( 
.A(n_1315),
.B(n_1350),
.Y(n_1416)
);

OAI21xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1342),
.A2(n_1224),
.B(n_1239),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1242),
.A2(n_1284),
.B(n_1264),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1333),
.A2(n_1351),
.B(n_1303),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1273),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1281),
.A2(n_1293),
.B(n_1303),
.C(n_1318),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1253),
.A2(n_1327),
.B1(n_1337),
.B2(n_1249),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1297),
.Y(n_1423)
);

OAI211xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1230),
.A2(n_1243),
.B(n_1252),
.C(n_1281),
.Y(n_1424)
);

OAI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1299),
.A2(n_1295),
.B1(n_1269),
.B2(n_1320),
.C(n_1285),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1320),
.B(n_1269),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1301),
.B(n_1302),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1301),
.B(n_1314),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1254),
.A2(n_1235),
.B(n_1343),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1222),
.A2(n_1343),
.B(n_1339),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1222),
.A2(n_1339),
.B(n_1235),
.Y(n_1431)
);

INVx5_ASAP7_75t_L g1432 ( 
.A(n_1347),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1323),
.Y(n_1433)
);

NAND2x1p5_ASAP7_75t_L g1434 ( 
.A(n_1323),
.B(n_1347),
.Y(n_1434)
);

BUFx8_ASAP7_75t_SL g1435 ( 
.A(n_1323),
.Y(n_1435)
);

CKINVDCx8_ASAP7_75t_R g1436 ( 
.A(n_1316),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1309),
.A2(n_1222),
.B(n_1261),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1309),
.A2(n_1257),
.B(n_1261),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1316),
.A2(n_1232),
.B(n_1259),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1231),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1334),
.A2(n_1212),
.B1(n_1233),
.B2(n_1234),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1234),
.A2(n_911),
.B1(n_1212),
.B2(n_1188),
.Y(n_1442)
);

AND2x2_ASAP7_75t_SL g1443 ( 
.A(n_1334),
.B(n_911),
.Y(n_1443)
);

NOR2xp67_ASAP7_75t_L g1444 ( 
.A(n_1228),
.B(n_879),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1255),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1234),
.A2(n_926),
.B1(n_1111),
.B2(n_1108),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1234),
.A2(n_911),
.B1(n_1212),
.B2(n_1188),
.Y(n_1447)
);

AO21x1_ASAP7_75t_L g1448 ( 
.A1(n_1334),
.A2(n_1188),
.B(n_1186),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1289),
.B(n_1225),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1334),
.A2(n_1212),
.B1(n_1233),
.B2(n_1234),
.Y(n_1450)
);

O2A1O1Ixp33_ASAP7_75t_SL g1451 ( 
.A1(n_1262),
.A2(n_1286),
.B(n_1349),
.C(n_1335),
.Y(n_1451)
);

AO31x2_ASAP7_75t_L g1452 ( 
.A1(n_1335),
.A2(n_1198),
.A3(n_1361),
.B(n_1349),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1352),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1322),
.A2(n_1198),
.B(n_1324),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1231),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1283),
.A2(n_1232),
.B(n_1332),
.Y(n_1456)
);

AOI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1283),
.A2(n_1232),
.B(n_1332),
.Y(n_1457)
);

CKINVDCx6p67_ASAP7_75t_R g1458 ( 
.A(n_1219),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1334),
.A2(n_1212),
.B1(n_1233),
.B2(n_1234),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1218),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1348),
.B(n_1270),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1326),
.A2(n_1356),
.B(n_1349),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1359),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1234),
.B(n_1108),
.Y(n_1464)
);

O2A1O1Ixp33_ASAP7_75t_SL g1465 ( 
.A1(n_1262),
.A2(n_1286),
.B(n_1349),
.C(n_1335),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1226),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1275),
.B(n_1108),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1322),
.A2(n_1198),
.B(n_1324),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1232),
.A2(n_1259),
.B(n_1329),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1326),
.A2(n_1356),
.B(n_1349),
.Y(n_1470)
);

O2A1O1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1233),
.A2(n_1262),
.B(n_1282),
.C(n_1335),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1325),
.B(n_1330),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1231),
.Y(n_1473)
);

BUFx2_ASAP7_75t_R g1474 ( 
.A(n_1228),
.Y(n_1474)
);

AOI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1234),
.A2(n_1212),
.B1(n_1233),
.B2(n_1111),
.C(n_960),
.Y(n_1475)
);

NAND3x1_ASAP7_75t_L g1476 ( 
.A(n_1234),
.B(n_1111),
.C(n_1115),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1254),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1231),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1232),
.A2(n_1259),
.B(n_1329),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1234),
.B(n_1108),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1325),
.B(n_1330),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1334),
.A2(n_1212),
.B1(n_1234),
.B2(n_911),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1326),
.A2(n_1356),
.B(n_1349),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1334),
.A2(n_1212),
.B1(n_1233),
.B2(n_1234),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1218),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1321),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1464),
.A2(n_1480),
.B1(n_1365),
.B2(n_1482),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1369),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1464),
.B(n_1480),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1419),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1482),
.A2(n_1459),
.B1(n_1441),
.B2(n_1450),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1363),
.B(n_1472),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1374),
.B(n_1409),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1419),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1369),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1441),
.A2(n_1484),
.B1(n_1450),
.B2(n_1459),
.Y(n_1496)
);

AND2x2_ASAP7_75t_SL g1497 ( 
.A(n_1443),
.B(n_1484),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1365),
.A2(n_1442),
.B1(n_1447),
.B2(n_1475),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1371),
.B(n_1461),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1367),
.A2(n_1449),
.B(n_1381),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1388),
.B(n_1380),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1481),
.B(n_1399),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1462),
.A2(n_1483),
.B(n_1470),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_SL g1504 ( 
.A1(n_1367),
.A2(n_1449),
.B(n_1411),
.Y(n_1504)
);

CKINVDCx16_ASAP7_75t_R g1505 ( 
.A(n_1368),
.Y(n_1505)
);

NAND2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1439),
.B(n_1412),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1426),
.B(n_1460),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1462),
.A2(n_1483),
.B(n_1470),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1364),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1463),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1485),
.B(n_1394),
.Y(n_1511)
);

AND2x6_ASAP7_75t_L g1512 ( 
.A(n_1366),
.B(n_1410),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1376),
.B(n_1475),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1440),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1376),
.B(n_1394),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1435),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1442),
.A2(n_1447),
.B1(n_1446),
.B2(n_1476),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1395),
.B(n_1398),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1400),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1372),
.B(n_1486),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1370),
.A2(n_1372),
.B1(n_1471),
.B2(n_1413),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1471),
.B(n_1455),
.Y(n_1522)
);

CKINVDCx14_ASAP7_75t_R g1523 ( 
.A(n_1458),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1445),
.Y(n_1524)
);

O2A1O1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1451),
.A2(n_1465),
.B(n_1413),
.C(n_1424),
.Y(n_1525)
);

AOI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1370),
.A2(n_1448),
.B1(n_1383),
.B2(n_1425),
.C(n_1417),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1404),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1390),
.A2(n_1430),
.B(n_1431),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1467),
.A2(n_1425),
.B(n_1429),
.C(n_1424),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1373),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1473),
.B(n_1478),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1420),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1422),
.B(n_1415),
.Y(n_1533)
);

BUFx2_ASAP7_75t_SL g1534 ( 
.A(n_1382),
.Y(n_1534)
);

OR2x6_ASAP7_75t_L g1535 ( 
.A(n_1408),
.B(n_1407),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1408),
.A2(n_1421),
.B(n_1477),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1437),
.A2(n_1414),
.B(n_1396),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1400),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1416),
.B(n_1402),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1418),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1397),
.B(n_1466),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1433),
.Y(n_1542)
);

AND2x6_ASAP7_75t_L g1543 ( 
.A(n_1378),
.B(n_1401),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1384),
.B(n_1423),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1438),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1379),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1452),
.B(n_1378),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1436),
.A2(n_1453),
.B1(n_1392),
.B2(n_1474),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1392),
.A2(n_1444),
.B1(n_1432),
.B2(n_1427),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1452),
.B(n_1393),
.Y(n_1550)
);

OA21x2_ASAP7_75t_L g1551 ( 
.A1(n_1391),
.A2(n_1375),
.B(n_1479),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1428),
.B(n_1427),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1406),
.B(n_1405),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1387),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1387),
.B(n_1406),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1405),
.B(n_1389),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1400),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1428),
.B(n_1389),
.Y(n_1558)
);

OAI31xp33_ASAP7_75t_L g1559 ( 
.A1(n_1434),
.A2(n_1456),
.A3(n_1457),
.B(n_1377),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1386),
.B(n_1469),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1367),
.A2(n_1198),
.B(n_1335),
.Y(n_1561)
);

INVx6_ASAP7_75t_L g1562 ( 
.A(n_1463),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1363),
.B(n_1472),
.Y(n_1563)
);

O2A1O1Ixp5_ASAP7_75t_L g1564 ( 
.A1(n_1448),
.A2(n_1381),
.B(n_1233),
.C(n_1356),
.Y(n_1564)
);

NOR2xp67_ASAP7_75t_L g1565 ( 
.A(n_1444),
.B(n_1453),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1462),
.A2(n_1483),
.B(n_1470),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1369),
.Y(n_1567)
);

O2A1O1Ixp5_ASAP7_75t_L g1568 ( 
.A1(n_1448),
.A2(n_1381),
.B(n_1233),
.C(n_1356),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1385),
.A2(n_1468),
.B(n_1454),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1419),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_SL g1571 ( 
.A1(n_1367),
.A2(n_1198),
.B(n_1335),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1364),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1367),
.A2(n_1198),
.B(n_1335),
.Y(n_1573)
);

O2A1O1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1365),
.A2(n_1233),
.B(n_1262),
.C(n_1234),
.Y(n_1574)
);

O2A1O1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1365),
.A2(n_1233),
.B(n_1262),
.C(n_1234),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1374),
.B(n_1409),
.Y(n_1576)
);

AND2x2_ASAP7_75t_SL g1577 ( 
.A(n_1443),
.B(n_1441),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1364),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_R g1579 ( 
.A(n_1368),
.B(n_879),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1385),
.A2(n_1468),
.B(n_1454),
.Y(n_1580)
);

O2A1O1Ixp5_ASAP7_75t_L g1581 ( 
.A1(n_1448),
.A2(n_1381),
.B(n_1233),
.C(n_1356),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1403),
.Y(n_1582)
);

NOR2xp67_ASAP7_75t_L g1583 ( 
.A(n_1444),
.B(n_1453),
.Y(n_1583)
);

O2A1O1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1365),
.A2(n_1233),
.B(n_1262),
.C(n_1234),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1513),
.B(n_1502),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1507),
.B(n_1492),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1533),
.B(n_1555),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1560),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1535),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1490),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1563),
.B(n_1515),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1494),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1503),
.B(n_1508),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1528),
.B(n_1503),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1570),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1535),
.Y(n_1596)
);

AO21x2_ASAP7_75t_L g1597 ( 
.A1(n_1569),
.A2(n_1580),
.B(n_1540),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1545),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1566),
.B(n_1554),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1489),
.B(n_1505),
.Y(n_1600)
);

INVx4_ASAP7_75t_L g1601 ( 
.A(n_1543),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1550),
.B(n_1553),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1560),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1566),
.B(n_1558),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1514),
.B(n_1498),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1537),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1520),
.B(n_1547),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_1524),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1537),
.Y(n_1609)
);

OR2x6_ASAP7_75t_L g1610 ( 
.A(n_1504),
.B(n_1500),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1574),
.A2(n_1584),
.B(n_1575),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1551),
.Y(n_1612)
);

OR2x6_ASAP7_75t_L g1613 ( 
.A(n_1506),
.B(n_1561),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1488),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1526),
.A2(n_1556),
.B(n_1564),
.Y(n_1615)
);

AO21x2_ASAP7_75t_L g1616 ( 
.A1(n_1549),
.A2(n_1529),
.B(n_1521),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1514),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1498),
.B(n_1495),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1532),
.B(n_1571),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1531),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1567),
.B(n_1521),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1522),
.B(n_1511),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1501),
.B(n_1499),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1541),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1512),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1568),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1518),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1581),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1573),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1517),
.A2(n_1491),
.B(n_1496),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1525),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1539),
.B(n_1517),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1559),
.B(n_1576),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1512),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1496),
.A2(n_1491),
.B(n_1577),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1594),
.B(n_1559),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1589),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1598),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1594),
.B(n_1497),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1586),
.B(n_1552),
.Y(n_1640)
);

NOR2x1_ASAP7_75t_L g1641 ( 
.A(n_1616),
.B(n_1613),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1611),
.A2(n_1487),
.B(n_1523),
.Y(n_1642)
);

INVx4_ASAP7_75t_L g1643 ( 
.A(n_1601),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1594),
.B(n_1493),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1596),
.Y(n_1645)
);

INVxp33_ASAP7_75t_L g1646 ( 
.A(n_1600),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1613),
.B(n_1536),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1586),
.B(n_1487),
.Y(n_1648)
);

OR2x2_ASAP7_75t_SL g1649 ( 
.A(n_1615),
.B(n_1562),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1590),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1617),
.B(n_1542),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1604),
.B(n_1538),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1604),
.B(n_1538),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1612),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1617),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1592),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1587),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1602),
.B(n_1582),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1596),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1593),
.B(n_1599),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1599),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1592),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1595),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1588),
.B(n_1603),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1597),
.B(n_1510),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1642),
.A2(n_1630),
.B1(n_1635),
.B2(n_1611),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1657),
.B(n_1602),
.Y(n_1667)
);

AO21x2_ASAP7_75t_L g1668 ( 
.A1(n_1654),
.A2(n_1606),
.B(n_1609),
.Y(n_1668)
);

OAI221xp5_ASAP7_75t_SL g1669 ( 
.A1(n_1642),
.A2(n_1632),
.B1(n_1618),
.B2(n_1631),
.C(n_1605),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1656),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1642),
.A2(n_1630),
.B1(n_1635),
.B2(n_1610),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1649),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1648),
.A2(n_1631),
.B1(n_1610),
.B2(n_1548),
.Y(n_1673)
);

AOI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1648),
.A2(n_1621),
.B1(n_1627),
.B2(n_1618),
.C(n_1630),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1651),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1647),
.A2(n_1630),
.B1(n_1610),
.B2(n_1616),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1656),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1656),
.Y(n_1678)
);

AOI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1665),
.A2(n_1621),
.B1(n_1627),
.B2(n_1591),
.C(n_1605),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1647),
.A2(n_1610),
.B1(n_1616),
.B2(n_1629),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1665),
.A2(n_1591),
.B1(n_1585),
.B2(n_1622),
.C(n_1614),
.Y(n_1681)
);

OAI33xp33_ASAP7_75t_L g1682 ( 
.A1(n_1651),
.A2(n_1585),
.A3(n_1622),
.B1(n_1614),
.B2(n_1632),
.B3(n_1620),
.Y(n_1682)
);

AOI33xp33_ASAP7_75t_L g1683 ( 
.A1(n_1665),
.A2(n_1628),
.A3(n_1626),
.B1(n_1633),
.B2(n_1624),
.B3(n_1620),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1649),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1647),
.A2(n_1610),
.B1(n_1616),
.B2(n_1629),
.Y(n_1685)
);

OAI31xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1641),
.A2(n_1629),
.A3(n_1633),
.B(n_1619),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1662),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1664),
.Y(n_1688)
);

AND3x1_ASAP7_75t_L g1689 ( 
.A(n_1639),
.B(n_1544),
.C(n_1633),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1655),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1639),
.A2(n_1610),
.B1(n_1548),
.B2(n_1615),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1644),
.B(n_1607),
.Y(n_1692)
);

OR2x2_ASAP7_75t_SL g1693 ( 
.A(n_1640),
.B(n_1615),
.Y(n_1693)
);

OAI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1641),
.A2(n_1613),
.B1(n_1534),
.B2(n_1623),
.C(n_1619),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1637),
.B(n_1589),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1662),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1655),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1650),
.Y(n_1698)
);

OAI21xp33_ASAP7_75t_L g1699 ( 
.A1(n_1641),
.A2(n_1619),
.B(n_1607),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1640),
.B(n_1623),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_1647),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1644),
.B(n_1603),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_R g1703 ( 
.A(n_1643),
.B(n_1509),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1638),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1660),
.B(n_1603),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1647),
.A2(n_1613),
.B1(n_1634),
.B2(n_1625),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1646),
.A2(n_1626),
.B(n_1628),
.C(n_1634),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1662),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1663),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1649),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1670),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1677),
.Y(n_1712)
);

CKINVDCx6p67_ASAP7_75t_R g1713 ( 
.A(n_1672),
.Y(n_1713)
);

CKINVDCx14_ASAP7_75t_R g1714 ( 
.A(n_1703),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1681),
.B(n_1657),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1701),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1672),
.B(n_1660),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1678),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1668),
.Y(n_1719)
);

INVx4_ASAP7_75t_SL g1720 ( 
.A(n_1701),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1687),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1696),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1668),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1708),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1709),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1690),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1704),
.Y(n_1727)
);

INVx4_ASAP7_75t_SL g1728 ( 
.A(n_1701),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1704),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1697),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1701),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1679),
.B(n_1661),
.Y(n_1732)
);

INVx4_ASAP7_75t_L g1733 ( 
.A(n_1701),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1674),
.B(n_1661),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1684),
.B(n_1636),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1710),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1667),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1698),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1707),
.A2(n_1682),
.B(n_1686),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1667),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1669),
.B(n_1646),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1705),
.B(n_1636),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1705),
.B(n_1636),
.Y(n_1743)
);

OR2x6_ASAP7_75t_L g1744 ( 
.A(n_1706),
.B(n_1647),
.Y(n_1744)
);

NOR2x1_ASAP7_75t_L g1745 ( 
.A(n_1741),
.B(n_1707),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1736),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1720),
.B(n_1728),
.Y(n_1747)
);

OR2x6_ASAP7_75t_L g1748 ( 
.A(n_1739),
.B(n_1647),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1720),
.B(n_1688),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1739),
.B(n_1666),
.C(n_1741),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1715),
.A2(n_1671),
.B1(n_1691),
.B2(n_1673),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1711),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1734),
.B(n_1676),
.C(n_1683),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1713),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1736),
.Y(n_1755)
);

AOI222xp33_ASAP7_75t_L g1756 ( 
.A1(n_1715),
.A2(n_1699),
.B1(n_1639),
.B2(n_1694),
.C1(n_1626),
.C2(n_1700),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1734),
.B(n_1693),
.Y(n_1757)
);

INVxp33_ASAP7_75t_L g1758 ( 
.A(n_1737),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1720),
.B(n_1688),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1736),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1720),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1737),
.B(n_1693),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1720),
.B(n_1728),
.Y(n_1763)
);

NOR3xp33_ASAP7_75t_SL g1764 ( 
.A(n_1732),
.B(n_1578),
.C(n_1572),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1730),
.Y(n_1765)
);

BUFx3_ASAP7_75t_L g1766 ( 
.A(n_1713),
.Y(n_1766)
);

NAND2x1_ASAP7_75t_L g1767 ( 
.A(n_1733),
.B(n_1695),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1720),
.B(n_1692),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1713),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1711),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1728),
.B(n_1692),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1735),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1738),
.Y(n_1773)
);

OAI33xp33_ASAP7_75t_L g1774 ( 
.A1(n_1732),
.A2(n_1675),
.A3(n_1652),
.B1(n_1653),
.B2(n_1658),
.B3(n_1663),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1728),
.B(n_1702),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1712),
.Y(n_1776)
);

NAND2x1p5_ASAP7_75t_L g1777 ( 
.A(n_1733),
.B(n_1643),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1712),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1726),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1718),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1718),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1721),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1740),
.B(n_1683),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1728),
.B(n_1702),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1721),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1735),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1722),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1728),
.B(n_1695),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1722),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1740),
.B(n_1675),
.Y(n_1790)
);

OAI211xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1714),
.A2(n_1685),
.B(n_1680),
.C(n_1527),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1755),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1747),
.B(n_1735),
.Y(n_1793)
);

AOI311xp33_ASAP7_75t_L g1794 ( 
.A1(n_1783),
.A2(n_1725),
.A3(n_1724),
.B(n_1729),
.C(n_1727),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1772),
.B(n_1730),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1747),
.B(n_1731),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1747),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1755),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1760),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1763),
.B(n_1731),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1763),
.B(n_1731),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1760),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1763),
.B(n_1731),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1750),
.B(n_1714),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1751),
.B(n_1742),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1745),
.B(n_1742),
.Y(n_1806)
);

NOR2xp67_ASAP7_75t_L g1807 ( 
.A(n_1761),
.B(n_1733),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1767),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1752),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1786),
.B(n_1765),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1779),
.B(n_1726),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1746),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1770),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1766),
.B(n_1733),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1754),
.B(n_1742),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1776),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1762),
.B(n_1743),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1778),
.Y(n_1818)
);

NAND2xp67_ASAP7_75t_SL g1819 ( 
.A(n_1749),
.B(n_1717),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1780),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1790),
.B(n_1743),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1768),
.B(n_1743),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1781),
.Y(n_1823)
);

NAND2x1p5_ASAP7_75t_L g1824 ( 
.A(n_1766),
.B(n_1733),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1753),
.A2(n_1744),
.B1(n_1716),
.B2(n_1647),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1782),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1768),
.B(n_1717),
.Y(n_1827)
);

NOR3x1_ASAP7_75t_L g1828 ( 
.A(n_1761),
.B(n_1659),
.C(n_1645),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1792),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1793),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_SL g1831 ( 
.A1(n_1804),
.A2(n_1748),
.B1(n_1769),
.B2(n_1757),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1807),
.B(n_1769),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1792),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1811),
.B(n_1757),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1797),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1806),
.B(n_1756),
.Y(n_1836)
);

OA21x2_ASAP7_75t_L g1837 ( 
.A1(n_1799),
.A2(n_1723),
.B(n_1719),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1793),
.B(n_1788),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1797),
.B(n_1788),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1817),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1805),
.B(n_1774),
.Y(n_1841)
);

NOR2x1_ASAP7_75t_L g1842 ( 
.A(n_1799),
.B(n_1767),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1798),
.B(n_1758),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1802),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1814),
.B(n_1689),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1797),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1827),
.B(n_1822),
.Y(n_1847)
);

NOR2x1_ASAP7_75t_L g1848 ( 
.A(n_1802),
.B(n_1748),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1811),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1827),
.B(n_1788),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1809),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1822),
.B(n_1771),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1809),
.Y(n_1853)
);

AOI222xp33_ASAP7_75t_L g1854 ( 
.A1(n_1825),
.A2(n_1791),
.B1(n_1758),
.B2(n_1771),
.C1(n_1639),
.C2(n_1784),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1812),
.B(n_1748),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1820),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1839),
.B(n_1796),
.Y(n_1857)
);

AOI21xp33_ASAP7_75t_SL g1858 ( 
.A1(n_1841),
.A2(n_1824),
.B(n_1810),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1843),
.B(n_1821),
.Y(n_1859)
);

INVx1_ASAP7_75t_SL g1860 ( 
.A(n_1839),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1830),
.B(n_1812),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1839),
.B(n_1796),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1831),
.A2(n_1748),
.B1(n_1794),
.B2(n_1824),
.C(n_1815),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1844),
.Y(n_1864)
);

AOI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1836),
.A2(n_1800),
.B1(n_1803),
.B2(n_1801),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1838),
.B(n_1800),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1849),
.B(n_1814),
.Y(n_1867)
);

OAI21xp33_ASAP7_75t_SL g1868 ( 
.A1(n_1848),
.A2(n_1808),
.B(n_1803),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1838),
.B(n_1801),
.Y(n_1869)
);

AOI221xp5_ASAP7_75t_L g1870 ( 
.A1(n_1849),
.A2(n_1823),
.B1(n_1820),
.B2(n_1813),
.C(n_1816),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1829),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1847),
.B(n_1814),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1829),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1829),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1845),
.A2(n_1784),
.B1(n_1775),
.B2(n_1824),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1855),
.B(n_1810),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1835),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1877),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1860),
.B(n_1847),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1877),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1864),
.B(n_1833),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1865),
.B(n_1835),
.Y(n_1882)
);

INVxp67_ASAP7_75t_L g1883 ( 
.A(n_1857),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1858),
.B(n_1832),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1866),
.B(n_1869),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1861),
.B(n_1834),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1876),
.B(n_1846),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1867),
.B(n_1834),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1871),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1872),
.B(n_1840),
.Y(n_1890)
);

AOI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1884),
.A2(n_1875),
.B1(n_1857),
.B2(n_1862),
.Y(n_1891)
);

OAI21xp33_ASAP7_75t_L g1892 ( 
.A1(n_1879),
.A2(n_1859),
.B(n_1868),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1883),
.B(n_1862),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1887),
.B(n_1863),
.Y(n_1894)
);

A2O1A1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1878),
.A2(n_1848),
.B(n_1880),
.C(n_1882),
.Y(n_1895)
);

NAND5xp2_ASAP7_75t_L g1896 ( 
.A(n_1885),
.B(n_1870),
.C(n_1854),
.D(n_1873),
.E(n_1874),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1886),
.A2(n_1846),
.B(n_1832),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1881),
.A2(n_1832),
.B(n_1842),
.Y(n_1898)
);

AOI211xp5_ASAP7_75t_L g1899 ( 
.A1(n_1888),
.A2(n_1832),
.B(n_1833),
.C(n_1839),
.Y(n_1899)
);

NOR2x1_ASAP7_75t_L g1900 ( 
.A(n_1881),
.B(n_1833),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1890),
.A2(n_1850),
.B1(n_1840),
.B2(n_1852),
.Y(n_1901)
);

NAND4xp25_ASAP7_75t_L g1902 ( 
.A(n_1889),
.B(n_1842),
.C(n_1840),
.D(n_1850),
.Y(n_1902)
);

OAI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1882),
.A2(n_1808),
.B1(n_1764),
.B2(n_1777),
.C(n_1762),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1900),
.Y(n_1904)
);

XNOR2xp5_ASAP7_75t_L g1905 ( 
.A(n_1891),
.B(n_1565),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1895),
.A2(n_1853),
.B(n_1851),
.Y(n_1906)
);

INVx4_ASAP7_75t_L g1907 ( 
.A(n_1893),
.Y(n_1907)
);

INVx1_ASAP7_75t_SL g1908 ( 
.A(n_1897),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1899),
.B(n_1795),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1894),
.A2(n_1852),
.B1(n_1826),
.B2(n_1818),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1901),
.B(n_1516),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1908),
.B(n_1892),
.Y(n_1912)
);

NOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1904),
.B(n_1902),
.Y(n_1913)
);

INVxp67_ASAP7_75t_L g1914 ( 
.A(n_1909),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_L g1915 ( 
.A(n_1906),
.B(n_1898),
.C(n_1903),
.Y(n_1915)
);

NOR3xp33_ASAP7_75t_L g1916 ( 
.A(n_1907),
.B(n_1896),
.C(n_1853),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1911),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1910),
.Y(n_1918)
);

INVx2_ASAP7_75t_SL g1919 ( 
.A(n_1913),
.Y(n_1919)
);

OAI32xp33_ASAP7_75t_L g1920 ( 
.A1(n_1916),
.A2(n_1856),
.A3(n_1851),
.B1(n_1777),
.B2(n_1817),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1912),
.Y(n_1921)
);

NAND3xp33_ASAP7_75t_L g1922 ( 
.A(n_1915),
.B(n_1905),
.C(n_1856),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1914),
.B(n_1608),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1917),
.B(n_1823),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1919),
.B(n_1918),
.Y(n_1925)
);

NAND4xp25_ASAP7_75t_SL g1926 ( 
.A(n_1922),
.B(n_1795),
.C(n_1749),
.D(n_1759),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1921),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1925),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1928),
.Y(n_1929)
);

OAI22x1_ASAP7_75t_L g1930 ( 
.A1(n_1929),
.A2(n_1927),
.B1(n_1923),
.B2(n_1926),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1929),
.A2(n_1924),
.B(n_1920),
.Y(n_1931)
);

XNOR2xp5_ASAP7_75t_L g1932 ( 
.A(n_1930),
.B(n_1583),
.Y(n_1932)
);

OAI332xp33_ASAP7_75t_L g1933 ( 
.A1(n_1931),
.A2(n_1819),
.A3(n_1579),
.B1(n_1828),
.B2(n_1785),
.B3(n_1787),
.C1(n_1789),
.C2(n_1773),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_SL g1934 ( 
.A1(n_1932),
.A2(n_1562),
.B1(n_1546),
.B2(n_1530),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1933),
.A2(n_1837),
.B1(n_1773),
.B2(n_1777),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1934),
.Y(n_1936)
);

OR2x2_ASAP7_75t_SL g1937 ( 
.A(n_1936),
.B(n_1935),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1937),
.B(n_1837),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_SL g1939 ( 
.A1(n_1938),
.A2(n_1759),
.B(n_1775),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1939),
.A2(n_1837),
.B1(n_1716),
.B2(n_1819),
.Y(n_1940)
);

AOI211xp5_ASAP7_75t_L g1941 ( 
.A1(n_1940),
.A2(n_1716),
.B(n_1519),
.C(n_1557),
.Y(n_1941)
);


endmodule