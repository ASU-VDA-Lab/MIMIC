module fake_jpeg_20599_n_397 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_397);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_397;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_8),
.B(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_47),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_48),
.B(n_59),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_60),
.Y(n_93)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g120 ( 
.A(n_53),
.Y(n_120)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_35),
.Y(n_55)
);

AO22x1_ASAP7_75t_L g129 ( 
.A1(n_55),
.A2(n_74),
.B1(n_87),
.B2(n_34),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_14),
.B(n_13),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_26),
.B(n_40),
.C(n_18),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_20),
.B(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_12),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_66),
.B(n_71),
.Y(n_135)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_70),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_33),
.B(n_0),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_33),
.B(n_10),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_73),
.B(n_0),
.Y(n_136)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_83),
.Y(n_97)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_34),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_24),
.Y(n_109)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_90),
.B(n_118),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_43),
.B1(n_23),
.B2(n_41),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_92),
.A2(n_121),
.B1(n_127),
.B2(n_134),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_R g180 ( 
.A(n_98),
.B(n_10),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_64),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_100),
.A2(n_107),
.B1(n_122),
.B2(n_57),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_23),
.B1(n_27),
.B2(n_39),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_110),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_29),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_45),
.B(n_17),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_81),
.A2(n_87),
.B1(n_55),
.B2(n_53),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_51),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_22),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_124),
.B(n_128),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_24),
.B1(n_39),
.B2(n_29),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_46),
.B(n_16),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_25),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_133),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_25),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_77),
.A2(n_16),
.B1(n_38),
.B2(n_30),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_136),
.B(n_2),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_84),
.B(n_38),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_22),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_93),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_142),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_97),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_69),
.C(n_84),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_179),
.C(n_126),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_17),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_165),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_91),
.B(n_30),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_28),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_102),
.A2(n_78),
.B1(n_18),
.B2(n_40),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_108),
.B1(n_130),
.B2(n_112),
.Y(n_193)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_88),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_161),
.Y(n_199)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx6_ASAP7_75t_SL g207 ( 
.A(n_157),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_98),
.A2(n_28),
.B(n_40),
.C(n_18),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_82),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_159),
.B(n_178),
.Y(n_188)
);

NAND2x1_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_121),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_160),
.A2(n_162),
.B(n_108),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_22),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_19),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_166),
.B(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_95),
.B(n_61),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_0),
.B(n_1),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_96),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_168),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_121),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_123),
.A2(n_1),
.B(n_2),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_173),
.Y(n_212)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_172),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_101),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_50),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_138),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_119),
.A2(n_2),
.B(n_3),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_102),
.A2(n_49),
.B1(n_3),
.B2(n_4),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_117),
.C(n_47),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_5),
.Y(n_192)
);

CKINVDCx6p67_ASAP7_75t_R g181 ( 
.A(n_105),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_182),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_117),
.B(n_4),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_183),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_219),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_149),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_191),
.B(n_205),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_192),
.A2(n_209),
.B(n_175),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_193),
.A2(n_141),
.B1(n_179),
.B2(n_154),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_204),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_114),
.B1(n_112),
.B2(n_104),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_198),
.A2(n_200),
.B1(n_120),
.B2(n_173),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_111),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_111),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_139),
.B(n_104),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_178),
.B(n_99),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_211),
.B(n_215),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_139),
.A2(n_115),
.B1(n_125),
.B2(n_120),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_162),
.B1(n_172),
.B2(n_115),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_145),
.B(n_106),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_165),
.B(n_113),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_216),
.B(n_217),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_158),
.B(n_144),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_146),
.B(n_120),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_218),
.B(n_220),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_99),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_185),
.A2(n_159),
.B1(n_180),
.B2(n_162),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_224),
.A2(n_231),
.B(n_240),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_225),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_206),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_228),
.Y(n_279)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_230),
.Y(n_259)
);

NAND2x1_ASAP7_75t_SL g231 ( 
.A(n_191),
.B(n_156),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_237),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_140),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_217),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_186),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_160),
.B1(n_141),
.B2(n_174),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_243),
.A2(n_204),
.B1(n_205),
.B2(n_186),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_187),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_244),
.Y(n_272)
);

BUFx12_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_254),
.B(n_190),
.Y(n_271)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_202),
.A2(n_160),
.B(n_142),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_252),
.B1(n_253),
.B2(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_251),
.B1(n_189),
.B2(n_220),
.Y(n_278)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_221),
.A2(n_169),
.B1(n_167),
.B2(n_163),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_255),
.A2(n_277),
.B1(n_248),
.B2(n_231),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_184),
.C(n_221),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_262),
.C(n_264),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_282),
.B1(n_232),
.B2(n_226),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_216),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_215),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_275),
.C(n_281),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_208),
.A3(n_188),
.B1(n_196),
.B2(n_199),
.C1(n_200),
.C2(n_147),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_273),
.B(n_276),
.Y(n_297)
);

A2O1A1O1Ixp25_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_194),
.B(n_200),
.C(n_188),
.D(n_209),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_177),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_222),
.B(n_223),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_252),
.A2(n_200),
.B1(n_198),
.B2(n_196),
.Y(n_277)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_224),
.A2(n_192),
.B(n_213),
.Y(n_280)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_280),
.A2(n_211),
.B(n_143),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_213),
.C(n_197),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_243),
.A2(n_198),
.B1(n_193),
.B2(n_189),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_284),
.A2(n_285),
.B1(n_277),
.B2(n_255),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_250),
.B1(n_227),
.B2(n_254),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_290),
.Y(n_309)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_257),
.A2(n_237),
.B1(n_246),
.B2(n_248),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_305),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_265),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_248),
.B(n_238),
.C(n_231),
.Y(n_291)
);

AOI22x1_ASAP7_75t_L g328 ( 
.A1(n_291),
.A2(n_245),
.B1(n_126),
.B2(n_207),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_249),
.Y(n_292)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_293),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_226),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_298),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_230),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_273),
.B1(n_257),
.B2(n_259),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_229),
.C(n_247),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_264),
.C(n_266),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_270),
.Y(n_301)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_301),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_251),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_197),
.Y(n_303)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_303),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_271),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_306),
.Y(n_315)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_262),
.B(n_198),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_299),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_312),
.A2(n_318),
.B1(n_287),
.B2(n_295),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_316),
.C(n_292),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_281),
.C(n_276),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_317),
.A2(n_289),
.B1(n_297),
.B2(n_285),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_287),
.A2(n_280),
.B1(n_259),
.B2(n_272),
.Y(n_318)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_323),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_275),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_296),
.Y(n_334)
);

OAI32xp33_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_198),
.A3(n_241),
.B1(n_245),
.B2(n_89),
.Y(n_323)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_263),
.Y(n_327)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_328),
.A2(n_323),
.B1(n_304),
.B2(n_286),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_309),
.Y(n_329)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_329),
.Y(n_350)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_309),
.Y(n_333)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_333),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_338),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_335),
.B(n_345),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_344),
.Y(n_347)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_341),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_296),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_316),
.A2(n_295),
.B(n_300),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_340),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_297),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_284),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_343),
.C(n_312),
.Y(n_352)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_326),
.A2(n_291),
.B(n_298),
.C(n_305),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_290),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_305),
.B(n_291),
.C(n_288),
.D(n_183),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_346),
.A2(n_328),
.B1(n_291),
.B2(n_325),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_332),
.A2(n_315),
.B1(n_317),
.B2(n_327),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_349),
.A2(n_356),
.B1(n_342),
.B2(n_336),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_351),
.B(n_352),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_344),
.A2(n_315),
.B(n_328),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_360),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_330),
.A2(n_311),
.B1(n_291),
.B2(n_324),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_346),
.A2(n_308),
.B(n_311),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_357),
.A2(n_5),
.B(n_6),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_320),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_365),
.Y(n_378)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_357),
.B(n_340),
.CI(n_343),
.CON(n_362),
.SN(n_362)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_359),
.Y(n_377)
);

MAJx2_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_334),
.C(n_338),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_364),
.A2(n_370),
.B(n_371),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_347),
.A2(n_324),
.B1(n_320),
.B2(n_321),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_349),
.A2(n_319),
.B1(n_201),
.B2(n_163),
.Y(n_366)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_239),
.C(n_171),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_354),
.C(n_350),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_369),
.B(n_365),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_347),
.A2(n_181),
.B(n_157),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_353),
.A2(n_348),
.B(n_358),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_367),
.A2(n_352),
.B1(n_355),
.B2(n_350),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_372),
.A2(n_377),
.B1(n_361),
.B2(n_366),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_374),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_362),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_368),
.A2(n_355),
.B(n_360),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_380),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_363),
.A2(n_356),
.B(n_181),
.Y(n_380)
);

NOR2xp67_ASAP7_75t_SL g387 ( 
.A(n_381),
.B(n_372),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_383),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_378),
.B(n_362),
.Y(n_384)
);

AOI322xp5_ASAP7_75t_L g388 ( 
.A1(n_384),
.A2(n_385),
.A3(n_375),
.B1(n_377),
.B2(n_373),
.C1(n_364),
.C2(n_181),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_153),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_388),
.C(n_390),
.Y(n_391)
);

NOR2x1_ASAP7_75t_SL g390 ( 
.A(n_382),
.B(n_120),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_389),
.B(n_386),
.C(n_382),
.Y(n_392)
);

AOI321xp33_ASAP7_75t_L g394 ( 
.A1(n_392),
.A2(n_393),
.A3(n_153),
.B1(n_105),
.B2(n_89),
.C(n_113),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_381),
.C(n_153),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_394),
.A2(n_395),
.B(n_7),
.Y(n_396)
);

AOI321xp33_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_116),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_7),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_396),
.B(n_8),
.Y(n_397)
);


endmodule