module fake_netlist_5_1039_n_830 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_830);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_830;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_629;
wire n_590;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_804;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_647;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_826;
wire n_335;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_185;
wire n_243;
wire n_183;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_673;
wire n_631;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_680;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_813;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_772;
wire n_691;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_781;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_332;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_795;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_754;
wire n_712;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_348;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_74),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_11),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_67),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_120),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_5),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_76),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_42),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_59),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_64),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_8),
.Y(n_190)
);

INVx4_ASAP7_75t_R g191 ( 
.A(n_146),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_109),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_48),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_73),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_116),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_103),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_53),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_164),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_1),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_66),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_128),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_37),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_19),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_161),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_56),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_27),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_33),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_16),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_40),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_85),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_30),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_47),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_99),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_90),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_131),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_35),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_95),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_14),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_162),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_68),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_113),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_117),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_51),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_122),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_93),
.Y(n_239)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_190),
.A2(n_0),
.B(n_1),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

BUFx8_ASAP7_75t_SL g242 ( 
.A(n_179),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_198),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_0),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_206),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_230),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_179),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_177),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

AND2x4_ASAP7_75t_L g262 ( 
.A(n_197),
.B(n_18),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_178),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_184),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_5),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_188),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_196),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_182),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_207),
.B(n_6),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

OAI22x1_ASAP7_75t_L g271 ( 
.A1(n_200),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_202),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_215),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_216),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

OA22x2_ASAP7_75t_SL g277 ( 
.A1(n_239),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_195),
.B(n_9),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_10),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_229),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_193),
.B(n_12),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

AND2x4_ASAP7_75t_L g284 ( 
.A(n_237),
.B(n_20),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_176),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_180),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_241),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_241),
.Y(n_289)
);

AND3x2_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_191),
.C(n_193),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_243),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_244),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_247),
.Y(n_294)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_265),
.C(n_282),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_261),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_181),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_246),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_12),
.Y(n_307)
);

NOR3xp33_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_185),
.C(n_183),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_246),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

BUFx6f_ASAP7_75t_SL g312 ( 
.A(n_249),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_248),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_253),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_261),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_253),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_254),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_249),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_260),
.B(n_187),
.Y(n_322)
);

AOI21x1_ASAP7_75t_L g323 ( 
.A1(n_254),
.A2(n_238),
.B(n_235),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_SL g324 ( 
.A(n_271),
.B(n_186),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_258),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_242),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_258),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_258),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_260),
.B(n_189),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_284),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_269),
.B(n_192),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_245),
.A2(n_233),
.B1(n_232),
.B2(n_228),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_255),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_259),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_259),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_266),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_286),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_306),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_285),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_262),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_262),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_286),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_329),
.Y(n_345)
);

AND2x2_ASAP7_75t_SL g346 ( 
.A(n_308),
.B(n_262),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_292),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_286),
.Y(n_348)
);

A2O1A1Ixp33_ASAP7_75t_L g349 ( 
.A1(n_311),
.A2(n_279),
.B(n_263),
.C(n_281),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_297),
.B(n_261),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_286),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_261),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_330),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_322),
.Y(n_359)
);

BUFx12f_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_320),
.B(n_264),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_322),
.A2(n_255),
.B1(n_252),
.B2(n_203),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_272),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_290),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_273),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_298),
.B(n_194),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_318),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_274),
.Y(n_368)
);

NAND2xp33_ASAP7_75t_L g369 ( 
.A(n_305),
.B(n_201),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_321),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_316),
.B(n_205),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_323),
.A2(n_277),
.B1(n_209),
.B2(n_211),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_291),
.B(n_266),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_324),
.A2(n_240),
.B1(n_267),
.B2(n_270),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_324),
.B(n_208),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_312),
.A2(n_213),
.B1(n_214),
.B2(n_217),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_335),
.A2(n_240),
.B1(n_267),
.B2(n_270),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_293),
.B(n_275),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_302),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_302),
.Y(n_381)
);

BUFx6f_ASAP7_75t_SL g382 ( 
.A(n_294),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_296),
.B(n_272),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_303),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_300),
.B(n_272),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_334),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_L g387 ( 
.A(n_305),
.B(n_222),
.Y(n_387)
);

INVx8_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_301),
.B(n_276),
.Y(n_389)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_303),
.B(n_275),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g391 ( 
.A(n_337),
.B(n_283),
.C(n_280),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_336),
.A2(n_256),
.B1(n_240),
.B2(n_268),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_334),
.A2(n_227),
.B1(n_225),
.B2(n_223),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_276),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_305),
.B(n_336),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_325),
.B(n_276),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_287),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_288),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_304),
.B(n_276),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_304),
.B(n_280),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_314),
.B(n_280),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_SL g402 ( 
.A(n_287),
.B(n_280),
.Y(n_402)
);

NOR2x1p5_ASAP7_75t_L g403 ( 
.A(n_314),
.B(n_242),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_325),
.B(n_283),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_315),
.A2(n_283),
.B1(n_268),
.B2(n_15),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_367),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_359),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_358),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_354),
.A2(n_295),
.B(n_287),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_345),
.A2(n_283),
.B1(n_315),
.B2(n_319),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_340),
.B(n_326),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_341),
.B(n_317),
.Y(n_413)
);

O2A1O1Ixp33_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_319),
.B(n_317),
.C(n_289),
.Y(n_414)
);

AO21x2_ASAP7_75t_L g415 ( 
.A1(n_338),
.A2(n_289),
.B(n_288),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_341),
.A2(n_295),
.B(n_287),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_344),
.B(n_327),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_365),
.B(n_13),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_343),
.B(n_327),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_343),
.B(n_328),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_378),
.A2(n_328),
.B(n_295),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_342),
.A2(n_346),
.B1(n_375),
.B2(n_348),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_363),
.A2(n_361),
.B(n_353),
.Y(n_423)
);

AND2x2_ASAP7_75t_SL g424 ( 
.A(n_405),
.B(n_362),
.Y(n_424)
);

NAND2xp33_ASAP7_75t_L g425 ( 
.A(n_390),
.B(n_349),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_351),
.B(n_295),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_368),
.B(n_21),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_339),
.B(n_22),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_373),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_388),
.B(n_13),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_394),
.A2(n_92),
.B(n_173),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_23),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_395),
.B(n_24),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_374),
.B(n_14),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_388),
.B(n_15),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_376),
.B(n_16),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_379),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_347),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_355),
.B(n_380),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_350),
.B(n_17),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_403),
.Y(n_442)
);

O2A1O1Ixp33_ASAP7_75t_L g443 ( 
.A1(n_392),
.A2(n_17),
.B(n_25),
.C(n_26),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_388),
.B(n_28),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_R g446 ( 
.A(n_360),
.B(n_29),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_384),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_383),
.A2(n_31),
.B(n_32),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_386),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_352),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_372),
.Y(n_452)
);

AND2x2_ASAP7_75t_SL g453 ( 
.A(n_377),
.B(n_34),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_393),
.B(n_36),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_356),
.B(n_357),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_399),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_370),
.B(n_38),
.Y(n_457)
);

OAI21xp33_ASAP7_75t_L g458 ( 
.A1(n_366),
.A2(n_39),
.B(n_41),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_390),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_399),
.B(n_43),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_400),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_400),
.B(n_401),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_401),
.Y(n_463)
);

NOR3xp33_ASAP7_75t_L g464 ( 
.A(n_371),
.B(n_44),
.C(n_45),
.Y(n_464)
);

OAI21xp33_ASAP7_75t_L g465 ( 
.A1(n_369),
.A2(n_46),
.B(n_49),
.Y(n_465)
);

NOR3xp33_ASAP7_75t_L g466 ( 
.A(n_391),
.B(n_50),
.C(n_52),
.Y(n_466)
);

OAI21xp33_ASAP7_75t_L g467 ( 
.A1(n_387),
.A2(n_54),
.B(n_55),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_385),
.B(n_57),
.Y(n_468)
);

AOI21xp33_ASAP7_75t_L g469 ( 
.A1(n_389),
.A2(n_58),
.B(n_60),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_390),
.B(n_61),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_396),
.A2(n_62),
.B(n_63),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_382),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_390),
.B(n_71),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_382),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

AO21x2_ASAP7_75t_L g476 ( 
.A1(n_422),
.A2(n_79),
.B(n_80),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_448),
.Y(n_477)
);

OAI21x1_ASAP7_75t_SL g478 ( 
.A1(n_443),
.A2(n_81),
.B(n_82),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_423),
.A2(n_397),
.B(n_402),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_439),
.Y(n_480)
);

AO31x2_ASAP7_75t_L g481 ( 
.A1(n_418),
.A2(n_83),
.A3(n_84),
.B(n_86),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_R g482 ( 
.A(n_412),
.B(n_87),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_440),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_409),
.B(n_397),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_440),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_463),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_413),
.A2(n_88),
.B(n_89),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_407),
.B(n_91),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_456),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_462),
.A2(n_94),
.B(n_96),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_421),
.A2(n_175),
.B(n_98),
.Y(n_492)
);

OAI21xp33_ASAP7_75t_SL g493 ( 
.A1(n_424),
.A2(n_172),
.B(n_100),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

AO31x2_ASAP7_75t_L g495 ( 
.A1(n_437),
.A2(n_97),
.A3(n_102),
.B(n_104),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_406),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_408),
.B(n_110),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_417),
.B(n_111),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_413),
.B(n_112),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_115),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_419),
.A2(n_121),
.B(n_123),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_438),
.B(n_124),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_452),
.Y(n_503)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_435),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_420),
.B(n_411),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_434),
.A2(n_125),
.B(n_126),
.Y(n_506)
);

AO31x2_ASAP7_75t_L g507 ( 
.A1(n_434),
.A2(n_129),
.A3(n_130),
.B(n_132),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_425),
.A2(n_133),
.B(n_134),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_416),
.A2(n_171),
.B(n_137),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_136),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_455),
.B(n_138),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_447),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_460),
.A2(n_426),
.B(n_468),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_450),
.B(n_139),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_410),
.A2(n_141),
.B(n_142),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_415),
.A2(n_143),
.B(n_144),
.Y(n_516)
);

OAI22x1_ASAP7_75t_L g517 ( 
.A1(n_442),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_517)
);

AO21x1_ASAP7_75t_L g518 ( 
.A1(n_454),
.A2(n_150),
.B(n_151),
.Y(n_518)
);

OAI21x1_ASAP7_75t_SL g519 ( 
.A1(n_429),
.A2(n_457),
.B(n_471),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_427),
.Y(n_520)
);

OAI22x1_ASAP7_75t_L g521 ( 
.A1(n_441),
.A2(n_474),
.B1(n_436),
.B2(n_431),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_428),
.A2(n_153),
.B(n_157),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_451),
.B(n_158),
.Y(n_524)
);

OAI21xp33_ASAP7_75t_L g525 ( 
.A1(n_453),
.A2(n_159),
.B(n_163),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_430),
.B(n_165),
.Y(n_526)
);

BUFx4_ASAP7_75t_SL g527 ( 
.A(n_459),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_430),
.A2(n_166),
.B(n_167),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_415),
.A2(n_168),
.B(n_433),
.Y(n_529)
);

OAI22x1_ASAP7_75t_L g530 ( 
.A1(n_445),
.A2(n_446),
.B1(n_473),
.B2(n_470),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_414),
.B(n_458),
.Y(n_531)
);

AO31x2_ASAP7_75t_L g532 ( 
.A1(n_470),
.A2(n_473),
.A3(n_433),
.B(n_472),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_465),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_503),
.B(n_464),
.Y(n_534)
);

NOR2xp67_ASAP7_75t_L g535 ( 
.A(n_530),
.B(n_432),
.Y(n_535)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_500),
.A2(n_467),
.B(n_469),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_469),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_522),
.B(n_449),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_477),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_526),
.A2(n_466),
.B(n_513),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_504),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_524),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_522),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_499),
.A2(n_531),
.B(n_505),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_520),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_490),
.B(n_487),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g547 ( 
.A1(n_519),
.A2(n_498),
.B(n_501),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_528),
.A2(n_509),
.B(n_515),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_493),
.A2(n_485),
.B(n_483),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_510),
.Y(n_550)
);

AO21x2_ASAP7_75t_L g551 ( 
.A1(n_506),
.A2(n_491),
.B(n_516),
.Y(n_551)
);

AO21x2_ASAP7_75t_L g552 ( 
.A1(n_478),
.A2(n_497),
.B(n_511),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_527),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_494),
.B(n_480),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_502),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_486),
.Y(n_556)
);

AO21x2_ASAP7_75t_L g557 ( 
.A1(n_476),
.A2(n_508),
.B(n_514),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_523),
.Y(n_558)
);

CKINVDCx16_ASAP7_75t_R g559 ( 
.A(n_482),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_533),
.A2(n_490),
.B(n_486),
.Y(n_560)
);

OR2x6_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_525),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_487),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_533),
.A2(n_488),
.B(n_512),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_484),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_518),
.A2(n_496),
.B(n_489),
.Y(n_565)
);

OAI21x1_ASAP7_75t_SL g566 ( 
.A1(n_517),
.A2(n_495),
.B(n_507),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_532),
.B(n_495),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_532),
.A2(n_507),
.B(n_495),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_481),
.B(n_365),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_481),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g571 ( 
.A1(n_479),
.A2(n_423),
.B(n_492),
.Y(n_571)
);

CKINVDCx11_ASAP7_75t_R g572 ( 
.A(n_477),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_503),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_479),
.A2(n_423),
.B(n_492),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_486),
.Y(n_575)
);

OAI21x1_ASAP7_75t_SL g576 ( 
.A1(n_518),
.A2(n_506),
.B(n_491),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_503),
.Y(n_578)
);

AO21x2_ASAP7_75t_L g579 ( 
.A1(n_529),
.A2(n_519),
.B(n_513),
.Y(n_579)
);

NAND3xp33_ASAP7_75t_L g580 ( 
.A(n_503),
.B(n_418),
.C(n_437),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_486),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_486),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_562),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_577),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_581),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_581),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_561),
.B(n_577),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_556),
.Y(n_588)
);

NAND2x1p5_ASAP7_75t_L g589 ( 
.A(n_563),
.B(n_550),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_543),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_561),
.A2(n_537),
.B1(n_580),
.B2(n_534),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_543),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_546),
.B(n_542),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_561),
.B(n_569),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_539),
.Y(n_595)
);

BUFx4f_ASAP7_75t_SL g596 ( 
.A(n_539),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_575),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_582),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_554),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_546),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_548),
.A2(n_571),
.B(n_574),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_543),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_578),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_560),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_560),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_554),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_549),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_549),
.Y(n_608)
);

INVxp67_ASAP7_75t_SL g609 ( 
.A(n_578),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_567),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_568),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_567),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_566),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_538),
.Y(n_614)
);

BUFx4f_ASAP7_75t_SL g615 ( 
.A(n_541),
.Y(n_615)
);

AO21x2_ASAP7_75t_L g616 ( 
.A1(n_576),
.A2(n_544),
.B(n_551),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_558),
.Y(n_617)
);

OA21x2_ASAP7_75t_L g618 ( 
.A1(n_540),
.A2(n_565),
.B(n_535),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_572),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_555),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_538),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_558),
.Y(n_622)
);

AO21x1_ASAP7_75t_SL g623 ( 
.A1(n_564),
.A2(n_551),
.B(n_570),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_536),
.A2(n_580),
.B(n_579),
.Y(n_624)
);

NOR2x1_ASAP7_75t_L g625 ( 
.A(n_593),
.B(n_545),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_599),
.B(n_559),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_587),
.B(n_550),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_587),
.B(n_550),
.Y(n_628)
);

AO21x2_ASAP7_75t_L g629 ( 
.A1(n_624),
.A2(n_601),
.B(n_605),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_594),
.B(n_555),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_583),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_596),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_599),
.B(n_534),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_604),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_591),
.B(n_573),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_584),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_594),
.B(n_555),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_604),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_591),
.A2(n_595),
.B(n_607),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_600),
.B(n_570),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_621),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_600),
.B(n_570),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_588),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_603),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_588),
.B(n_545),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_592),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_620),
.B(n_541),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_603),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_606),
.B(n_573),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_597),
.Y(n_650)
);

CKINVDCx16_ASAP7_75t_R g651 ( 
.A(n_619),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_597),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_609),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_605),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_598),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_595),
.A2(n_536),
.B1(n_547),
.B2(n_552),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_585),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_598),
.B(n_552),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_585),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_620),
.B(n_547),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_586),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_586),
.Y(n_662)
);

BUFx2_ASAP7_75t_SL g663 ( 
.A(n_592),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_611),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_613),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_611),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_617),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_620),
.B(n_579),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_606),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_615),
.B(n_572),
.Y(n_670)
);

INVxp67_ASAP7_75t_R g671 ( 
.A(n_624),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_613),
.Y(n_672)
);

CKINVDCx11_ASAP7_75t_R g673 ( 
.A(n_619),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_607),
.B(n_557),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_627),
.B(n_608),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_661),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_661),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_657),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_657),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_653),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_662),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_626),
.B(n_541),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_625),
.B(n_608),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_648),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_630),
.B(n_616),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_665),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_630),
.B(n_616),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_662),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_659),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_637),
.B(n_616),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_637),
.B(n_623),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_632),
.B(n_553),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_627),
.B(n_628),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_628),
.B(n_623),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_635),
.B(n_602),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_672),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_643),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_633),
.A2(n_673),
.B1(n_614),
.B2(n_669),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_674),
.B(n_612),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_644),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_651),
.A2(n_614),
.B1(n_672),
.B2(n_645),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_650),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_645),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_658),
.B(n_612),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_674),
.B(n_610),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_649),
.B(n_602),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_SL g707 ( 
.A1(n_651),
.A2(n_621),
.B1(n_663),
.B2(n_640),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_650),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_639),
.B(n_610),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_652),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_652),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_655),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_655),
.B(n_602),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_665),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_685),
.B(n_658),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_685),
.B(n_687),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_686),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_686),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_687),
.B(n_668),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_714),
.B(n_668),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_690),
.B(n_660),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_678),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_675),
.B(n_642),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_690),
.B(n_660),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_684),
.B(n_642),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_679),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_695),
.B(n_640),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_694),
.B(n_664),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_680),
.B(n_634),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_680),
.B(n_634),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_689),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_704),
.B(n_671),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_704),
.B(n_671),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_694),
.B(n_629),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_691),
.B(n_681),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_700),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_691),
.B(n_693),
.Y(n_737)
);

NOR3xp33_ASAP7_75t_L g738 ( 
.A(n_683),
.B(n_656),
.C(n_670),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_689),
.Y(n_739)
);

OAI221xp5_ASAP7_75t_SL g740 ( 
.A1(n_698),
.A2(n_654),
.B1(n_638),
.B2(n_667),
.C(n_590),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_699),
.B(n_654),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_696),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_706),
.B(n_638),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_699),
.B(n_666),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_742),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_725),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_719),
.B(n_703),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_716),
.B(n_696),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_734),
.B(n_629),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_736),
.B(n_709),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_718),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_734),
.B(n_629),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_719),
.B(n_701),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_718),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_715),
.B(n_724),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_717),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_722),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_726),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_742),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_731),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_724),
.B(n_705),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_731),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_735),
.B(n_677),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_739),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_739),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_727),
.B(n_723),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_756),
.Y(n_767)
);

INVxp33_ASAP7_75t_L g768 ( 
.A(n_766),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_748),
.B(n_761),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_745),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_750),
.A2(n_738),
.B1(n_735),
.B2(n_683),
.Y(n_771)
);

AOI32xp33_ASAP7_75t_L g772 ( 
.A1(n_753),
.A2(n_735),
.A3(n_733),
.B1(n_732),
.B2(n_737),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_746),
.B(n_755),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_760),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_760),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_763),
.A2(n_682),
.B1(n_707),
.B2(n_709),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_751),
.Y(n_777)
);

AOI32xp33_ASAP7_75t_L g778 ( 
.A1(n_749),
.A2(n_733),
.A3(n_732),
.B1(n_715),
.B2(n_721),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_759),
.A2(n_740),
.B(n_743),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_757),
.A2(n_729),
.B1(n_730),
.B2(n_741),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_777),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_768),
.A2(n_763),
.B1(n_749),
.B2(n_752),
.Y(n_782)
);

OAI221xp5_ASAP7_75t_SL g783 ( 
.A1(n_771),
.A2(n_759),
.B1(n_752),
.B2(n_758),
.C(n_745),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_L g784 ( 
.A(n_779),
.B(n_765),
.C(n_764),
.Y(n_784)
);

OAI21xp33_ASAP7_75t_SL g785 ( 
.A1(n_772),
.A2(n_755),
.B(n_747),
.Y(n_785)
);

AOI222xp33_ASAP7_75t_L g786 ( 
.A1(n_780),
.A2(n_720),
.B1(n_763),
.B2(n_692),
.C1(n_721),
.C2(n_754),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_781),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_784),
.A2(n_776),
.B1(n_773),
.B2(n_767),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_783),
.A2(n_776),
.B(n_770),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_782),
.B(n_769),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_785),
.A2(n_778),
.B1(n_721),
.B2(n_728),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_786),
.B(n_775),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_792),
.B(n_647),
.C(n_713),
.Y(n_793)
);

OAI321xp33_ASAP7_75t_L g794 ( 
.A1(n_789),
.A2(n_762),
.A3(n_676),
.B1(n_774),
.B2(n_744),
.C(n_697),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_788),
.B(n_728),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_787),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_791),
.B(n_728),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_793),
.B(n_790),
.Y(n_798)
);

AOI211xp5_ASAP7_75t_L g799 ( 
.A1(n_794),
.A2(n_647),
.B(n_712),
.C(n_702),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_798),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_799),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_798),
.A2(n_795),
.B1(n_796),
.B2(n_797),
.Y(n_802)
);

NAND4xp75_ASAP7_75t_L g803 ( 
.A(n_800),
.B(n_646),
.C(n_618),
.D(n_688),
.Y(n_803)
);

XNOR2xp5_ASAP7_75t_L g804 ( 
.A(n_802),
.B(n_801),
.Y(n_804)
);

XOR2x1_ASAP7_75t_L g805 ( 
.A(n_800),
.B(n_647),
.Y(n_805)
);

NAND4xp75_ASAP7_75t_L g806 ( 
.A(n_800),
.B(n_646),
.C(n_618),
.D(n_708),
.Y(n_806)
);

NOR2x1_ASAP7_75t_L g807 ( 
.A(n_801),
.B(n_590),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_804),
.B(n_807),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_SL g809 ( 
.A(n_805),
.B(n_803),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_806),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_807),
.Y(n_811)
);

XNOR2x1_ASAP7_75t_L g812 ( 
.A(n_804),
.B(n_590),
.Y(n_812)
);

NOR2x1_ASAP7_75t_L g813 ( 
.A(n_807),
.B(n_602),
.Y(n_813)
);

NOR2xp67_ASAP7_75t_L g814 ( 
.A(n_811),
.B(n_592),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_SL g815 ( 
.A1(n_808),
.A2(n_663),
.B1(n_592),
.B2(n_589),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_812),
.A2(n_720),
.B1(n_705),
.B2(n_711),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_810),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_817),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_814),
.Y(n_819)
);

AOI21xp33_ASAP7_75t_L g820 ( 
.A1(n_815),
.A2(n_816),
.B(n_813),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_814),
.Y(n_821)
);

OAI22x1_ASAP7_75t_L g822 ( 
.A1(n_818),
.A2(n_809),
.B1(n_720),
.B2(n_589),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_819),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_821),
.A2(n_592),
.B1(n_641),
.B2(n_667),
.Y(n_824)
);

AOI22x1_ASAP7_75t_L g825 ( 
.A1(n_822),
.A2(n_820),
.B1(n_589),
.B2(n_617),
.Y(n_825)
);

AO21x1_ASAP7_75t_L g826 ( 
.A1(n_823),
.A2(n_631),
.B(n_636),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_825),
.A2(n_826),
.B(n_824),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_827),
.A2(n_621),
.B(n_710),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_828),
.B(n_622),
.Y(n_829)
);

AOI21xp33_ASAP7_75t_SL g830 ( 
.A1(n_829),
.A2(n_557),
.B(n_618),
.Y(n_830)
);


endmodule