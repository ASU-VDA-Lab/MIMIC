module fake_jpeg_19100_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_60),
.Y(n_97)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_48),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_76),
.B1(n_91),
.B2(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_99),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_43),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_50),
.B1(n_44),
.B2(n_33),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_76),
.B1(n_91),
.B2(n_95),
.Y(n_118)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_83),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_87),
.Y(n_115)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_18),
.B1(n_21),
.B2(n_28),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_101),
.B1(n_16),
.B2(n_34),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_49),
.B1(n_28),
.B2(n_21),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_37),
.B(n_35),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_28),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_45),
.C(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_18),
.B1(n_17),
.B2(n_19),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_122),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_35),
.A3(n_41),
.B1(n_16),
.B2(n_30),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_124),
.B(n_94),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_125),
.B1(n_94),
.B2(n_87),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_34),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_32),
.B1(n_30),
.B2(n_25),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_32),
.B1(n_25),
.B2(n_20),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_75),
.B1(n_71),
.B2(n_70),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_146),
.B1(n_155),
.B2(n_126),
.Y(n_161)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_117),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_72),
.B(n_95),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_136),
.B(n_141),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_76),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_103),
.B(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_128),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_24),
.B(n_77),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_142),
.B(n_151),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_78),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_149),
.B(n_156),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_102),
.C(n_96),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_153),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_118),
.A2(n_78),
.B1(n_80),
.B2(n_75),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_150),
.B1(n_119),
.B2(n_116),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_102),
.B1(n_31),
.B2(n_29),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_27),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_125),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_82),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_112),
.A2(n_31),
.B(n_29),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_20),
.B1(n_29),
.B2(n_27),
.Y(n_155)
);

AOI22x1_ASAP7_75t_SL g156 ( 
.A1(n_109),
.A2(n_20),
.B1(n_29),
.B2(n_27),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_112),
.B1(n_125),
.B2(n_104),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_158),
.B1(n_164),
.B2(n_155),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_104),
.B1(n_107),
.B2(n_129),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_156),
.B(n_153),
.C(n_149),
.D(n_135),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_159),
.A2(n_174),
.B(n_143),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_167),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_163),
.B1(n_176),
.B2(n_180),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_122),
.B1(n_129),
.B2(n_107),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_117),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_168),
.B(n_169),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_144),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_139),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_178),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_128),
.C(n_123),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_173),
.B(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_119),
.B1(n_116),
.B2(n_113),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_179),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_183),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_132),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_187),
.A2(n_199),
.B1(n_200),
.B2(n_209),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_173),
.B(n_171),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_191),
.A2(n_195),
.B1(n_202),
.B2(n_166),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_197),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_149),
.B1(n_137),
.B2(n_145),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_186),
.A3(n_175),
.B1(n_170),
.B2(n_159),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_31),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_177),
.B1(n_179),
.B2(n_182),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_145),
.B1(n_150),
.B2(n_148),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_172),
.C(n_170),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_207),
.C(n_211),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_145),
.B1(n_132),
.B2(n_148),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_206),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_172),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_148),
.C(n_110),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_148),
.B1(n_131),
.B2(n_113),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_160),
.B(n_110),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_210),
.B(n_114),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_106),
.C(n_123),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_114),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_212),
.B(n_183),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_225),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_218),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_176),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_226),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_224),
.B1(n_200),
.B2(n_187),
.Y(n_242)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_194),
.A2(n_166),
.B1(n_165),
.B2(n_164),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_165),
.B(n_106),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_114),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_230),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_188),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_232),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_197),
.B(n_183),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_198),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_203),
.B(n_31),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_27),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_208),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_203),
.B(n_192),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_225),
.B1(n_217),
.B2(n_223),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_247),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_219),
.A2(n_191),
.B1(n_193),
.B2(n_207),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_249),
.B1(n_0),
.B2(n_2),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_246),
.B1(n_205),
.B2(n_231),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_211),
.C(n_195),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_251),
.C(n_213),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_199),
.B1(n_209),
.B2(n_196),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_219),
.A2(n_202),
.B1(n_205),
.B2(n_208),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_253),
.B(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_213),
.C(n_218),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_255),
.C(n_258),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_230),
.C(n_215),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_259),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_215),
.C(n_233),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_251),
.C(n_247),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_263),
.B1(n_240),
.B2(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

OAI31xp33_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_0),
.A3(n_1),
.B(n_2),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_265),
.A2(n_239),
.B1(n_237),
.B2(n_6),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_0),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_266),
.A2(n_267),
.B1(n_6),
.B2(n_7),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_271),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_235),
.B1(n_239),
.B2(n_242),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_267),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_244),
.B1(n_246),
.B2(n_6),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_7),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_4),
.C(n_5),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_278),
.C(n_266),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_261),
.A2(n_4),
.B(n_5),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_7),
.B(n_8),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_4),
.C(n_5),
.Y(n_278)
);

XOR2x1_ASAP7_75t_SL g279 ( 
.A(n_256),
.B(n_6),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_279),
.B(n_265),
.CI(n_264),
.CON(n_284),
.SN(n_284)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_288)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_283),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_258),
.C(n_261),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_286),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_259),
.C(n_8),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_274),
.C(n_276),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_288),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_273),
.B(n_271),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_269),
.B(n_10),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_290),
.A2(n_279),
.B(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_294),
.B(n_297),
.CI(n_293),
.CON(n_303),
.SN(n_303)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_269),
.C(n_10),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_286),
.B1(n_289),
.B2(n_281),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_285),
.B1(n_284),
.B2(n_12),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_303),
.A2(n_298),
.B(n_284),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_300),
.Y(n_308)
);

A2O1A1O1Ixp25_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_298),
.B(n_11),
.C(n_12),
.D(n_13),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_305),
.B(n_303),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_307),
.C(n_11),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_8),
.B(n_11),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_12),
.B(n_13),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_13),
.Y(n_313)
);


endmodule