module fake_jpeg_1662_n_19 (n_3, n_2, n_1, n_0, n_4, n_19);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_19;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_18;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g5 ( 
.A(n_3),
.Y(n_5)
);

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_0),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

AOI22xp5_ASAP7_75t_L g9 ( 
.A1(n_8),
.A2(n_6),
.B1(n_5),
.B2(n_7),
.Y(n_9)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_9),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_7),
.B(n_8),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_0),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_2),
.B1(n_9),
.B2(n_13),
.Y(n_16)
);

A2O1A1Ixp33_ASAP7_75t_SL g18 ( 
.A1(n_16),
.A2(n_17),
.B(n_15),
.C(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_18),
.Y(n_19)
);


endmodule