module fake_jpeg_16346_n_243 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_45),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

OR2x4_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_23),
.A2(n_3),
.B(n_5),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_60),
.C(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_11),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_5),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_22),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_22),
.A2(n_6),
.B(n_7),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_15),
.B(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_6),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_62),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_58),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_30),
.C(n_17),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_7),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_16),
.B(n_8),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_16),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_17),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_21),
.B1(n_34),
.B2(n_25),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_72),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_25),
.B1(n_37),
.B2(n_35),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_39),
.A2(n_37),
.B1(n_35),
.B2(n_33),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_63),
.B1(n_62),
.B2(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_83),
.Y(n_112)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_87),
.B(n_91),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_28),
.B1(n_33),
.B2(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_103),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_29),
.B1(n_32),
.B2(n_20),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_93),
.A2(n_81),
.B1(n_80),
.B2(n_94),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_41),
.B(n_9),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_56),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_102),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_41),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_29),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_36),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_32),
.B1(n_10),
.B2(n_27),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_27),
.B1(n_36),
.B2(n_10),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_46),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_116),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_72),
.A2(n_59),
.B(n_46),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_135),
.B(n_100),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_59),
.B(n_46),
.C(n_57),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_124),
.B(n_75),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_44),
.Y(n_113)
);

BUFx24_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_47),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_54),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_133),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_54),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_36),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_36),
.Y(n_128)
);

AO21x1_ASAP7_75t_SL g137 ( 
.A1(n_129),
.A2(n_116),
.B(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_130),
.B(n_89),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_68),
.B(n_69),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_90),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_134),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_121),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_122),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_107),
.B(n_89),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_140),
.B(n_161),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_145),
.B(n_124),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_96),
.B1(n_80),
.B2(n_88),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_120),
.B1(n_104),
.B2(n_106),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_152),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_129),
.B1(n_125),
.B2(n_109),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_133),
.B1(n_108),
.B2(n_111),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_69),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_100),
.Y(n_173)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_126),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_119),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_78),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_112),
.B(n_94),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_97),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_145),
.A2(n_110),
.B1(n_118),
.B2(n_124),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_165),
.B(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_97),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_180),
.C(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_174),
.B(n_176),
.Y(n_200)
);

NOR4xp25_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_114),
.C(n_95),
.D(n_78),
.Y(n_175)
);

NOR4xp25_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_162),
.C(n_158),
.D(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_84),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_84),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_181),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_140),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_141),
.A2(n_114),
.B(n_121),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_136),
.B(n_146),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_185),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_143),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_150),
.B(n_157),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_198),
.B(n_204),
.C(n_168),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_142),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_194),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_159),
.C(n_144),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_197),
.C(n_171),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_137),
.B1(n_148),
.B2(n_159),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_194),
.B1(n_203),
.B2(n_199),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_185),
.B1(n_179),
.B2(n_184),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_160),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_143),
.B(n_149),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_203),
.B(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_142),
.B(n_185),
.Y(n_203)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_202),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_210),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_188),
.B(n_183),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_209),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_207),
.A2(n_208),
.B(n_198),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_187),
.B(n_171),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_183),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_211),
.B(n_213),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_216),
.B1(n_195),
.B2(n_197),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_166),
.C(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_217),
.A2(n_196),
.B(n_186),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_192),
.B(n_191),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_219),
.A2(n_222),
.B(n_224),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_214),
.C(n_210),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_217),
.A2(n_192),
.B(n_191),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_212),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_228),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_208),
.A3(n_217),
.B1(n_215),
.B2(n_197),
.C1(n_200),
.C2(n_201),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_230),
.B(n_231),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_226),
.A2(n_201),
.A3(n_200),
.B1(n_190),
.B2(n_193),
.C1(n_181),
.C2(n_174),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_193),
.C(n_204),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_218),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_237),
.C(n_167),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_223),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_204),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_225),
.C(n_219),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_240),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_234),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_242),
.Y(n_243)
);


endmodule