module fake_aes_10528_n_574 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_574);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_574;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_73;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_67;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g67 ( .A(n_33), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_41), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_29), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_60), .Y(n_70) );
BUFx6f_ASAP7_75t_L g71 ( .A(n_5), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_28), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_59), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_40), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_16), .Y(n_75) );
BUFx6f_ASAP7_75t_L g76 ( .A(n_7), .Y(n_76) );
CKINVDCx16_ASAP7_75t_R g77 ( .A(n_24), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_0), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_46), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_10), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_39), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_14), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_52), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_0), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_25), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_56), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_55), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_37), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_20), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_44), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_18), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_27), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_34), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_49), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_35), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_62), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_36), .Y(n_97) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_53), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_8), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_14), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_17), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_65), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_48), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_43), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_63), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_64), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_47), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_7), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_50), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_57), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_89), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_89), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_98), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_98), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_86), .Y(n_115) );
CKINVDCx8_ASAP7_75t_R g116 ( .A(n_67), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_77), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_108), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_79), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_98), .Y(n_120) );
AND2x6_ASAP7_75t_L g121 ( .A(n_109), .B(n_23), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_71), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_109), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_95), .B(n_1), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_78), .Y(n_125) );
NOR2x1_ASAP7_75t_L g126 ( .A(n_68), .B(n_1), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_108), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_80), .B(n_2), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx4_ASAP7_75t_L g130 ( .A(n_98), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_104), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_104), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_75), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_106), .B(n_2), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_69), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_96), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_106), .B(n_3), .Y(n_138) );
INVx4_ASAP7_75t_L g139 ( .A(n_106), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_70), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_78), .Y(n_141) );
BUFx2_ASAP7_75t_L g142 ( .A(n_101), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_106), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_100), .B(n_3), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_100), .Y(n_145) );
BUFx12f_ASAP7_75t_L g146 ( .A(n_71), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_82), .B(n_4), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_106), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_122), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_118), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_122), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_118), .B(n_83), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_142), .B(n_110), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_111), .B(n_75), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_113), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
OR2x2_ASAP7_75t_SL g157 ( .A(n_134), .B(n_99), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_146), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_127), .B(n_88), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
INVx5_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_121), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_115), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_142), .B(n_87), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_111), .B(n_84), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_127), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_113), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
NOR2xp33_ASAP7_75t_SL g174 ( .A(n_116), .B(n_105), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_117), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_121), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
NAND2x1p5_ASAP7_75t_L g179 ( .A(n_144), .B(n_90), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_112), .B(n_71), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_112), .B(n_81), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_117), .B(n_137), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_133), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_123), .B(n_71), .Y(n_186) );
NAND3xp33_ASAP7_75t_L g187 ( .A(n_124), .B(n_71), .C(n_76), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_144), .B(n_92), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_139), .Y(n_189) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_123), .B(n_72), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_133), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_148), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_139), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_137), .B(n_116), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_121), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_148), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_139), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_148), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_136), .B(n_140), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_113), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_166), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_175), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_179), .B(n_140), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_168), .B(n_126), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_196), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_199), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_180), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_199), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_150), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_193), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_179), .B(n_136), .Y(n_212) );
CKINVDCx6p67_ASAP7_75t_R g213 ( .A(n_166), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_179), .B(n_147), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_180), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_196), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_152), .B(n_128), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_193), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_197), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_153), .B(n_145), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_190), .A2(n_103), .B1(n_105), .B2(n_79), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_168), .B(n_121), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_190), .A2(n_103), .B1(n_91), .B2(n_121), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_186), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_197), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_165), .B(n_145), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_186), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_180), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_190), .B(n_141), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_180), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_160), .B(n_141), .Y(n_231) );
INVx2_ASAP7_75t_SL g232 ( .A(n_188), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_154), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_161), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_154), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_154), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_154), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_161), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_164), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_164), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_168), .B(n_121), .Y(n_241) );
INVx4_ASAP7_75t_L g242 ( .A(n_158), .Y(n_242) );
INVx3_ASAP7_75t_SL g243 ( .A(n_188), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_170), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_170), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_168), .B(n_126), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_171), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_177), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_177), .Y(n_249) );
AND3x1_ASAP7_75t_L g250 ( .A(n_174), .B(n_119), .C(n_125), .Y(n_250) );
AND2x6_ASAP7_75t_SL g251 ( .A(n_184), .B(n_125), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_188), .A2(n_76), .B1(n_138), .B2(n_135), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_178), .Y(n_253) );
BUFx5_ASAP7_75t_L g254 ( .A(n_188), .Y(n_254) );
INVx5_ASAP7_75t_L g255 ( .A(n_188), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_188), .B(n_73), .Y(n_256) );
NAND2x1_ASAP7_75t_L g257 ( .A(n_233), .B(n_176), .Y(n_257) );
AOI21xp33_ASAP7_75t_L g258 ( .A1(n_232), .A2(n_195), .B(n_175), .Y(n_258) );
AOI22xp33_ASAP7_75t_SL g259 ( .A1(n_203), .A2(n_188), .B1(n_91), .B2(n_163), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_231), .A2(n_200), .B(n_192), .C(n_178), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_214), .B(n_157), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_243), .Y(n_262) );
CKINVDCx11_ASAP7_75t_R g263 ( .A(n_210), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g264 ( .A(n_255), .B(n_158), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_210), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_203), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_223), .A2(n_157), .B1(n_163), .B2(n_176), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_253), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_243), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_217), .B(n_182), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_213), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_213), .Y(n_272) );
INVxp67_ASAP7_75t_SL g273 ( .A(n_233), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_255), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_233), .Y(n_275) );
NOR2x1_ASAP7_75t_SL g276 ( .A(n_255), .B(n_176), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_214), .B(n_158), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_237), .A2(n_163), .B1(n_176), .B2(n_162), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_237), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_229), .A2(n_181), .B1(n_192), .B2(n_185), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_247), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_255), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_237), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_255), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_206), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_206), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_229), .A2(n_181), .B1(n_185), .B2(n_162), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_235), .A2(n_162), .B1(n_198), .B2(n_167), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_205), .A2(n_162), .B1(n_183), .B2(n_194), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_205), .A2(n_162), .B1(n_76), .B2(n_187), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_236), .A2(n_162), .B1(n_198), .B2(n_167), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_206), .Y(n_292) );
INVx4_ASAP7_75t_L g293 ( .A(n_242), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_242), .B(n_76), .Y(n_294) );
INVx2_ASAP7_75t_SL g295 ( .A(n_202), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_205), .B(n_167), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_253), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_253), .Y(n_298) );
OA21x2_ASAP7_75t_L g299 ( .A1(n_260), .A2(n_241), .B(n_222), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_281), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_261), .A2(n_250), .B1(n_220), .B2(n_226), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_270), .B(n_204), .Y(n_302) );
OAI211xp5_ASAP7_75t_SL g303 ( .A1(n_263), .A2(n_221), .B(n_246), .C(n_252), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_262), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_280), .A2(n_212), .B1(n_256), .B2(n_232), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_265), .B(n_224), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_268), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_263), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_262), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_261), .B(n_227), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_266), .B(n_251), .Y(n_311) );
CKINVDCx11_ASAP7_75t_R g312 ( .A(n_271), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_268), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_280), .A2(n_256), .B1(n_234), .B2(n_249), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_260), .B(n_256), .C(n_249), .Y(n_315) );
AOI221xp5_ASAP7_75t_SL g316 ( .A1(n_267), .A2(n_245), .B1(n_240), .B2(n_234), .C(n_239), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_277), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_259), .B(n_242), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_297), .A2(n_240), .B(n_245), .C(n_238), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_290), .B(n_120), .C(n_114), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_275), .A2(n_254), .B1(n_208), .B2(n_230), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_298), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_298), .Y(n_323) );
AOI21xp33_ASAP7_75t_L g324 ( .A1(n_295), .A2(n_202), .B(n_230), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_302), .B(n_244), .Y(n_325) );
OAI21xp33_ASAP7_75t_L g326 ( .A1(n_301), .A2(n_294), .B(n_287), .Y(n_326) );
OAI22xp33_ASAP7_75t_L g327 ( .A1(n_301), .A2(n_272), .B1(n_262), .B2(n_269), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_303), .A2(n_258), .B1(n_254), .B2(n_279), .Y(n_328) );
AOI222xp33_ASAP7_75t_L g329 ( .A1(n_310), .A2(n_283), .B1(n_296), .B2(n_273), .C1(n_215), .C2(n_208), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_300), .A2(n_254), .B1(n_215), .B2(n_293), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_309), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_317), .B(n_244), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_307), .B(n_248), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_300), .A2(n_254), .B1(n_293), .B2(n_228), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_307), .B(n_248), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_306), .B(n_211), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_311), .A2(n_254), .B1(n_269), .B2(n_294), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_306), .A2(n_254), .B1(n_262), .B2(n_282), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_314), .A2(n_254), .B1(n_211), .B2(n_218), .Y(n_340) );
AOI222xp33_ASAP7_75t_L g341 ( .A1(n_308), .A2(n_76), .B1(n_93), .B2(n_74), .C1(n_102), .C2(n_97), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_315), .A2(n_290), .B1(n_225), .B2(n_219), .C(n_218), .Y(n_342) );
AOI22xp33_ASAP7_75t_SL g343 ( .A1(n_318), .A2(n_254), .B1(n_276), .B2(n_264), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_313), .B(n_219), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_309), .Y(n_345) );
OAI211xp5_ASAP7_75t_L g346 ( .A1(n_312), .A2(n_85), .B(n_94), .C(n_289), .Y(n_346) );
AOI21xp33_ASAP7_75t_L g347 ( .A1(n_316), .A2(n_282), .B(n_274), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_313), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_336), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_325), .B(n_313), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_346), .A2(n_315), .B1(n_316), .B2(n_305), .C(n_324), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_336), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g353 ( .A1(n_326), .A2(n_321), .B1(n_319), .B2(n_320), .C(n_299), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_337), .A2(n_320), .B1(n_323), .B2(n_322), .C(n_107), .Y(n_354) );
INVx5_ASAP7_75t_L g355 ( .A(n_331), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_326), .A2(n_323), .B(n_322), .Y(n_356) );
OAI31xp33_ASAP7_75t_L g357 ( .A1(n_327), .A2(n_264), .A3(n_322), .B(n_323), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_325), .B(n_299), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g359 ( .A1(n_341), .A2(n_299), .B1(n_304), .B2(n_309), .C(n_288), .Y(n_359) );
NAND4xp25_ASAP7_75t_L g360 ( .A(n_341), .B(n_4), .C(n_5), .D(n_6), .Y(n_360) );
OAI31xp33_ASAP7_75t_L g361 ( .A1(n_332), .A2(n_278), .A3(n_291), .B(n_304), .Y(n_361) );
OA21x2_ASAP7_75t_L g362 ( .A1(n_347), .A2(n_225), .B(n_299), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_329), .A2(n_304), .B1(n_274), .B2(n_284), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_344), .B(n_304), .Y(n_364) );
AOI21xp5_ASAP7_75t_SL g365 ( .A1(n_340), .A2(n_292), .B(n_286), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_344), .B(n_6), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_332), .B(n_8), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_329), .A2(n_292), .B1(n_286), .B2(n_285), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_348), .Y(n_369) );
OAI22xp5_ASAP7_75t_SL g370 ( .A1(n_343), .A2(n_284), .B1(n_286), .B2(n_285), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g371 ( .A1(n_333), .A2(n_292), .B1(n_286), .B2(n_285), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_328), .A2(n_292), .B1(n_285), .B2(n_216), .Y(n_372) );
OAI21xp33_ASAP7_75t_L g373 ( .A1(n_333), .A2(n_113), .B(n_143), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_335), .B(n_348), .Y(n_374) );
AOI33xp33_ASAP7_75t_L g375 ( .A1(n_330), .A2(n_159), .A3(n_149), .B1(n_151), .B2(n_156), .B3(n_183), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_335), .B(n_9), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_331), .B(n_9), .Y(n_377) );
OR2x6_ASAP7_75t_L g378 ( .A(n_331), .B(n_257), .Y(n_378) );
OA21x2_ASAP7_75t_L g379 ( .A1(n_340), .A2(n_209), .B(n_207), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_331), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_367), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_367), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_374), .B(n_345), .Y(n_385) );
NAND4xp25_ASAP7_75t_SL g386 ( .A(n_368), .B(n_338), .C(n_334), .D(n_339), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_349), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_358), .B(n_345), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_350), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_374), .B(n_345), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_373), .A2(n_342), .B(n_345), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_349), .Y(n_393) );
OAI31xp33_ASAP7_75t_L g394 ( .A1(n_360), .A2(n_207), .A3(n_209), .B(n_156), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_358), .Y(n_395) );
OAI21xp33_ASAP7_75t_SL g396 ( .A1(n_368), .A2(n_345), .B(n_331), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_357), .B(n_113), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_366), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_352), .B(n_10), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_352), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_352), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_369), .B(n_11), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_366), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_360), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_355), .B(n_61), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_369), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_376), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_376), .B(n_12), .Y(n_408) );
AND3x1_ASAP7_75t_L g409 ( .A(n_357), .B(n_13), .C(n_15), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_351), .A2(n_359), .B1(n_363), .B2(n_377), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_364), .B(n_15), .Y(n_411) );
NAND2xp33_ASAP7_75t_SL g412 ( .A(n_370), .B(n_16), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_356), .B(n_114), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_380), .B(n_114), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_356), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_361), .A2(n_114), .B1(n_143), .B2(n_131), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_356), .B(n_143), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_355), .B(n_120), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_375), .B(n_143), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_355), .B(n_19), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_356), .B(n_120), .Y(n_421) );
OAI31xp33_ASAP7_75t_L g422 ( .A1(n_353), .A2(n_361), .A3(n_373), .B(n_372), .Y(n_422) );
INVx4_ASAP7_75t_L g423 ( .A(n_355), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_362), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_407), .B(n_355), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_423), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_384), .B(n_362), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_389), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_385), .B(n_362), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_399), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_385), .B(n_362), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_398), .B(n_354), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_412), .A2(n_365), .B1(n_371), .B2(n_378), .C(n_379), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_390), .B(n_379), .Y(n_436) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_409), .B(n_131), .C(n_143), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_399), .Y(n_438) );
AOI222xp33_ASAP7_75t_L g439 ( .A1(n_404), .A2(n_131), .B1(n_120), .B2(n_365), .C1(n_151), .C2(n_149), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_395), .B(n_379), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_391), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_403), .B(n_379), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_390), .B(n_378), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_395), .B(n_378), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_402), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_408), .B(n_378), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_388), .B(n_378), .Y(n_447) );
OR2x6_ASAP7_75t_L g448 ( .A(n_423), .B(n_131), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_411), .B(n_131), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_383), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_402), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_411), .B(n_120), .Y(n_452) );
NAND3xp33_ASAP7_75t_SL g453 ( .A(n_394), .B(n_21), .C(n_22), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_387), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_388), .B(n_26), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_391), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_412), .B(n_201), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g458 ( .A(n_410), .B(n_159), .C(n_194), .D(n_191), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_391), .B(n_30), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_393), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
OAI33xp33_ASAP7_75t_L g462 ( .A1(n_419), .A2(n_31), .A3(n_32), .B1(n_38), .B2(n_42), .B3(n_45), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_400), .B(n_51), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_423), .B(n_54), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_401), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_406), .B(n_58), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_405), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_386), .B(n_189), .C(n_169), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_406), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_422), .B(n_66), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_425), .B(n_414), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_430), .B(n_396), .Y(n_472) );
XOR2x2_ASAP7_75t_L g473 ( .A(n_457), .B(n_405), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_426), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_437), .A2(n_457), .B1(n_428), .B2(n_448), .Y(n_475) );
OAI31xp33_ASAP7_75t_L g476 ( .A1(n_435), .A2(n_397), .A3(n_420), .B(n_405), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g477 ( .A(n_470), .B(n_416), .C(n_414), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_443), .B(n_424), .Y(n_478) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_460), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_432), .B(n_424), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_447), .B(n_415), .Y(n_481) );
OAI21xp33_ASAP7_75t_L g482 ( .A1(n_429), .A2(n_420), .B(n_418), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_431), .B(n_433), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_438), .B(n_415), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_441), .B(n_420), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_446), .B(n_392), .Y(n_486) );
OR2x6_ASAP7_75t_L g487 ( .A(n_448), .B(n_441), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_447), .B(n_427), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_448), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_446), .A2(n_413), .B1(n_421), .B2(n_417), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_450), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_447), .B(n_413), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_444), .B(n_436), .Y(n_493) );
OAI31xp33_ASAP7_75t_L g494 ( .A1(n_456), .A2(n_421), .A3(n_417), .B(n_198), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_460), .B(n_155), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_454), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_469), .B(n_155), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_461), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_445), .B(n_155), .Y(n_499) );
XNOR2xp5_ASAP7_75t_L g500 ( .A(n_449), .B(n_189), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_465), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_451), .B(n_155), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_467), .B(n_155), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_469), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_452), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_464), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_440), .B(n_172), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_454), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_453), .A2(n_169), .B(n_173), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_475), .A2(n_453), .B(n_434), .C(n_452), .Y(n_510) );
XNOR2x1_ASAP7_75t_L g511 ( .A(n_473), .B(n_455), .Y(n_511) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_476), .B(n_439), .C(n_442), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_486), .B(n_459), .Y(n_513) );
XNOR2x1_ASAP7_75t_L g514 ( .A(n_473), .B(n_466), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_504), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_489), .A2(n_468), .B(n_458), .C(n_463), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_487), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_SL g518 ( .A1(n_486), .A2(n_468), .B(n_462), .C(n_191), .Y(n_518) );
XNOR2xp5_ASAP7_75t_L g519 ( .A(n_488), .B(n_173), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_483), .B(n_172), .Y(n_520) );
INVx3_ASAP7_75t_L g521 ( .A(n_487), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_477), .B(n_172), .C(n_201), .Y(n_522) );
OAI21xp5_ASAP7_75t_SL g523 ( .A1(n_485), .A2(n_201), .B(n_216), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_472), .Y(n_524) );
OAI21xp33_ASAP7_75t_SL g525 ( .A1(n_485), .A2(n_206), .B(n_216), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_480), .B(n_484), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_493), .B(n_479), .Y(n_527) );
XOR2x2_ASAP7_75t_L g528 ( .A(n_500), .B(n_478), .Y(n_528) );
AOI211xp5_ASAP7_75t_L g529 ( .A1(n_505), .A2(n_479), .B(n_494), .C(n_482), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_505), .A2(n_471), .B1(n_509), .B2(n_501), .C(n_498), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_493), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_502), .B(n_508), .C(n_493), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_481), .Y(n_533) );
XNOR2xp5_ASAP7_75t_L g534 ( .A(n_492), .B(n_481), .Y(n_534) );
AOI211xp5_ASAP7_75t_L g535 ( .A1(n_481), .A2(n_490), .B(n_499), .C(n_503), .Y(n_535) );
OAI221xp5_ASAP7_75t_SL g536 ( .A1(n_495), .A2(n_497), .B1(n_507), .B2(n_491), .C(n_496), .Y(n_536) );
NAND2xp33_ASAP7_75t_SL g537 ( .A(n_489), .B(n_428), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_506), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_476), .B(n_486), .C(n_472), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_486), .B(n_425), .Y(n_540) );
XNOR2x1_ASAP7_75t_L g541 ( .A(n_473), .B(n_308), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_476), .A2(n_489), .B(n_412), .C(n_475), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_474), .Y(n_543) );
BUFx2_ASAP7_75t_L g544 ( .A(n_487), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_475), .A2(n_437), .B(n_457), .Y(n_545) );
NAND5xp2_ASAP7_75t_L g546 ( .A(n_542), .B(n_510), .C(n_545), .D(n_516), .E(n_523), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_540), .Y(n_547) );
AOI21xp33_ASAP7_75t_SL g548 ( .A1(n_541), .A2(n_542), .B(n_539), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_524), .A2(n_537), .B1(n_512), .B2(n_511), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_515), .Y(n_550) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_544), .A2(n_521), .B1(n_517), .B2(n_527), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_538), .B(n_531), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_517), .B(n_521), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_514), .A2(n_513), .B1(n_528), .B2(n_535), .Y(n_554) );
NOR3xp33_ASAP7_75t_SL g555 ( .A(n_530), .B(n_523), .C(n_536), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_533), .A2(n_529), .B1(n_532), .B2(n_520), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_526), .Y(n_557) );
AOI211xp5_ASAP7_75t_L g558 ( .A1(n_548), .A2(n_519), .B(n_525), .C(n_522), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_550), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_546), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_549), .A2(n_534), .B1(n_515), .B2(n_526), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_557), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_547), .B(n_543), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_563), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_562), .B(n_555), .Y(n_565) );
AOI211xp5_ASAP7_75t_L g566 ( .A1(n_560), .A2(n_546), .B(n_551), .C(n_554), .Y(n_566) );
XOR2x2_ASAP7_75t_L g567 ( .A(n_566), .B(n_561), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_565), .A2(n_559), .B1(n_553), .B2(n_556), .Y(n_568) );
BUFx3_ASAP7_75t_L g569 ( .A(n_567), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_568), .B(n_564), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_569), .B(n_558), .Y(n_571) );
XOR2xp5_ASAP7_75t_L g572 ( .A(n_571), .B(n_570), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_572), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_573), .A2(n_552), .B(n_518), .Y(n_574) );
endmodule