module fake_jpeg_1506_n_159 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_19),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_58),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_38),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_65),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_50),
.Y(n_65)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_59),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_80),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_55),
.B1(n_61),
.B2(n_59),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_67),
.B1(n_69),
.B2(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_60),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_55),
.B1(n_45),
.B2(n_38),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_53),
.B1(n_46),
.B2(n_42),
.Y(n_95)
);

AO22x2_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_51),
.B1(n_44),
.B2(n_39),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_42),
.B1(n_69),
.B2(n_44),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_50),
.B(n_39),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_47),
.B(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_48),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_94),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_66),
.B(n_85),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_90),
.C(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_62),
.B(n_48),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_68),
.B1(n_67),
.B2(n_46),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_93),
.B1(n_95),
.B2(n_81),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_98),
.B1(n_16),
.B2(n_36),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_49),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_100),
.Y(n_107)
);

AOI22x1_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_47),
.B1(n_49),
.B2(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_0),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_29),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_119),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_74),
.B1(n_2),
.B2(n_4),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

AOI22x1_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_37),
.B1(n_34),
.B2(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_117),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_28),
.C(n_27),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_23),
.C(n_9),
.Y(n_124)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_26),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_1),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_10),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_5),
.B(n_6),
.Y(n_121)
);

AOI221xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_14),
.B1(n_15),
.B2(n_114),
.C(n_128),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_124),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_25),
.C(n_24),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_126),
.C(n_128),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_127),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_7),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_12),
.C(n_13),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_103),
.A2(n_13),
.B(n_14),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_119),
.B1(n_117),
.B2(n_111),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_140),
.A2(n_132),
.B1(n_131),
.B2(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_121),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_145),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_137),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_135),
.B1(n_140),
.B2(n_136),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_150),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_152),
.A2(n_146),
.B(n_151),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_153),
.C(n_145),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_153),
.B(n_144),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_157),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_138),
.B(n_124),
.Y(n_159)
);


endmodule