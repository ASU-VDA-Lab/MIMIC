module fake_jpeg_23028_n_28 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_28);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_28;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_26;
wire n_17;
wire n_25;
wire n_15;

INVx5_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp33_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_12),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_0),
.C(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_2),
.Y(n_20)
);

AO22x1_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

AND2x6_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_10),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_22),
.C(n_15),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_26),
.A2(n_23),
.B(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);


endmodule