module real_aes_10563_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_1806, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_1806;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_1797;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1768;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_1712;
wire n_991;
wire n_667;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_1740;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_1404;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1699;
wire n_419;
wire n_730;
wire n_1023;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_1749;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_1772;
wire n_831;
wire n_487;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_1790;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_719;
wire n_1343;
wire n_465;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_1691;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1777;
wire n_444;
wire n_1200;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_1352;
wire n_729;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1272 ( .A(n_0), .Y(n_1272) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_1), .A2(n_153), .B1(n_457), .B2(n_698), .C(n_699), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g754 ( .A1(n_1), .A2(n_308), .B1(n_755), .B2(n_756), .C(n_758), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g1475 ( .A1(n_2), .A2(n_299), .B1(n_1449), .B2(n_1457), .Y(n_1475) );
INVx1_ASAP7_75t_L g785 ( .A(n_3), .Y(n_785) );
INVx1_ASAP7_75t_L g919 ( .A(n_4), .Y(n_919) );
OAI221xp5_ASAP7_75t_L g1253 ( .A1(n_5), .A2(n_274), .B1(n_712), .B2(n_934), .C(n_936), .Y(n_1253) );
OAI22xp33_ASAP7_75t_SL g1283 ( .A1(n_5), .A2(n_274), .B1(n_1284), .B2(n_1285), .Y(n_1283) );
INVxp33_ASAP7_75t_L g1249 ( .A(n_6), .Y(n_1249) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_6), .A2(n_93), .B1(n_424), .B2(n_999), .C(n_1278), .Y(n_1277) );
AOI22xp33_ASAP7_75t_SL g1126 ( .A1(n_7), .A2(n_136), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_7), .A2(n_55), .B1(n_996), .B2(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1270 ( .A(n_8), .Y(n_1270) );
AOI221xp5_ASAP7_75t_L g1309 ( .A1(n_9), .A2(n_232), .B1(n_1310), .B2(n_1311), .C(n_1312), .Y(n_1309) );
INVx1_ASAP7_75t_L g1343 ( .A(n_9), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_10), .A2(n_61), .B1(n_599), .B2(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g674 ( .A(n_10), .Y(n_674) );
XNOR2x2_ASAP7_75t_L g1119 ( .A(n_11), .B(n_1120), .Y(n_1119) );
OAI22xp33_ASAP7_75t_L g1700 ( .A1(n_12), .A2(n_67), .B1(n_1701), .B2(n_1703), .Y(n_1700) );
OAI22xp33_ASAP7_75t_L g1711 ( .A1(n_12), .A2(n_164), .B1(n_327), .B2(n_1712), .Y(n_1711) );
AOI22xp5_ASAP7_75t_L g1476 ( .A1(n_13), .A2(n_248), .B1(n_1465), .B2(n_1471), .Y(n_1476) );
AOI22xp33_ASAP7_75t_SL g1130 ( .A1(n_14), .A2(n_55), .B1(n_1108), .B2(n_1131), .Y(n_1130) );
AOI21xp33_ASAP7_75t_L g1153 ( .A1(n_14), .A2(n_578), .B(n_820), .Y(n_1153) );
CKINVDCx5p33_ASAP7_75t_R g1081 ( .A(n_15), .Y(n_1081) );
INVxp67_ASAP7_75t_L g1034 ( .A(n_16), .Y(n_1034) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_16), .A2(n_58), .B1(n_389), .B2(n_416), .C(n_914), .Y(n_1061) );
CKINVDCx16_ASAP7_75t_R g1503 ( .A(n_17), .Y(n_1503) );
INVxp33_ASAP7_75t_L g795 ( .A(n_18), .Y(n_795) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_18), .A2(n_72), .B1(n_858), .B2(n_860), .C(n_861), .Y(n_857) );
INVx1_ASAP7_75t_L g1143 ( .A(n_19), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_19), .A2(n_257), .B1(n_820), .B2(n_996), .Y(n_1155) );
INVx1_ASAP7_75t_L g1695 ( .A(n_20), .Y(n_1695) );
OAI222xp33_ASAP7_75t_L g1707 ( .A1(n_20), .A2(n_205), .B1(n_280), .B2(n_943), .C1(n_1708), .C2(n_1710), .Y(n_1707) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_21), .A2(n_300), .B1(n_568), .B2(n_616), .C(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g657 ( .A(n_21), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g1190 ( .A(n_22), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_23), .A2(n_296), .B1(n_374), .B2(n_379), .Y(n_373) );
INVxp67_ASAP7_75t_SL g516 ( .A(n_23), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g1306 ( .A1(n_24), .A2(n_310), .B1(n_910), .B2(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1330 ( .A(n_24), .Y(n_1330) );
INVx1_ASAP7_75t_L g971 ( .A(n_25), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_25), .A2(n_52), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
OAI221xp5_ASAP7_75t_L g1030 ( .A1(n_26), .A2(n_109), .B1(n_934), .B2(n_935), .C(n_1031), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_26), .A2(n_109), .B1(n_910), .B2(n_1059), .Y(n_1058) );
INVxp67_ASAP7_75t_SL g1361 ( .A(n_27), .Y(n_1361) );
AOI221xp5_ASAP7_75t_L g1379 ( .A1(n_27), .A2(n_288), .B1(n_645), .B2(n_755), .C(n_914), .Y(n_1379) );
INVxp33_ASAP7_75t_L g963 ( .A(n_28), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_28), .A2(n_74), .B1(n_995), .B2(n_996), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_29), .A2(n_293), .B1(n_771), .B2(n_824), .Y(n_823) );
INVxp67_ASAP7_75t_SL g875 ( .A(n_29), .Y(n_875) );
XNOR2xp5_ASAP7_75t_L g1753 ( .A(n_30), .B(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g318 ( .A(n_31), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g1697 ( .A1(n_32), .A2(n_98), .B1(n_1698), .B2(n_1699), .Y(n_1697) );
AOI22xp33_ASAP7_75t_SL g1729 ( .A1(n_32), .A2(n_98), .B1(n_1728), .B2(n_1730), .Y(n_1729) );
INVx1_ASAP7_75t_L g1319 ( .A(n_33), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g1338 ( .A1(n_33), .A2(n_270), .B1(n_486), .B2(n_858), .Y(n_1338) );
CKINVDCx5p33_ASAP7_75t_R g1225 ( .A(n_34), .Y(n_1225) );
AOI22xp5_ASAP7_75t_L g1448 ( .A1(n_35), .A2(n_142), .B1(n_1449), .B2(n_1457), .Y(n_1448) );
OAI221xp5_ASAP7_75t_L g968 ( .A1(n_36), .A2(n_169), .B1(n_705), .B2(n_711), .C(n_715), .Y(n_968) );
OAI33xp33_ASAP7_75t_L g1001 ( .A1(n_36), .A2(n_169), .A3(n_430), .B1(n_750), .B2(n_1002), .B3(n_1806), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_37), .A2(n_195), .B1(n_1461), .B2(n_1490), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_38), .A2(n_59), .B1(n_379), .B2(n_910), .Y(n_909) );
OAI221xp5_ASAP7_75t_L g933 ( .A1(n_38), .A2(n_59), .B1(n_934), .B2(n_935), .C(n_936), .Y(n_933) );
AOI21xp33_ASAP7_75t_L g1088 ( .A1(n_39), .A2(n_624), .B(n_1009), .Y(n_1088) );
AOI221xp5_ASAP7_75t_L g1112 ( .A1(n_39), .A2(n_83), .B1(n_459), .B2(n_490), .C(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g397 ( .A(n_40), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_40), .A2(n_251), .B1(n_447), .B2(n_457), .C(n_464), .Y(n_446) );
INVx1_ASAP7_75t_L g805 ( .A(n_41), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_42), .A2(n_291), .B1(n_450), .B2(n_563), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_42), .A2(n_213), .B1(n_599), .B2(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g1718 ( .A(n_43), .Y(n_1718) );
AOI22xp33_ASAP7_75t_L g1738 ( .A1(n_43), .A2(n_203), .B1(n_917), .B2(n_1739), .Y(n_1738) );
INVx1_ASAP7_75t_L g1325 ( .A(n_44), .Y(n_1325) );
AOI22xp33_ASAP7_75t_L g1335 ( .A1(n_44), .A2(n_279), .B1(n_493), .B2(n_1336), .Y(n_1335) );
OAI222xp33_ASAP7_75t_L g1767 ( .A1(n_45), .A2(n_156), .B1(n_234), .B2(n_1768), .C1(n_1770), .C2(n_1771), .Y(n_1767) );
AOI221xp5_ASAP7_75t_L g1793 ( .A1(n_45), .A2(n_156), .B1(n_1794), .B2(n_1796), .C(n_1797), .Y(n_1793) );
AO221x2_ASAP7_75t_L g1477 ( .A1(n_46), .A2(n_215), .B1(n_1465), .B2(n_1471), .C(n_1478), .Y(n_1477) );
AOI22x1_ASAP7_75t_SL g1685 ( .A1(n_46), .A2(n_1686), .B1(n_1740), .B2(n_1741), .Y(n_1685) );
INVx1_ASAP7_75t_L g1740 ( .A(n_46), .Y(n_1740) );
AOI22xp33_ASAP7_75t_L g1748 ( .A1(n_46), .A2(n_1749), .B1(n_1752), .B2(n_1799), .Y(n_1748) );
AOI22xp5_ASAP7_75t_L g1469 ( .A1(n_47), .A2(n_113), .B1(n_1449), .B2(n_1457), .Y(n_1469) );
CKINVDCx16_ASAP7_75t_R g339 ( .A(n_48), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g1124 ( .A(n_49), .Y(n_1124) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_50), .Y(n_637) );
AOI22xp5_ASAP7_75t_SL g1507 ( .A1(n_51), .A2(n_209), .B1(n_1461), .B2(n_1465), .Y(n_1507) );
INVx1_ASAP7_75t_L g976 ( .A(n_52), .Y(n_976) );
INVxp67_ASAP7_75t_SL g1360 ( .A(n_53), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g1380 ( .A1(n_53), .A2(n_186), .B1(n_907), .B2(n_1292), .Y(n_1380) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_54), .A2(n_102), .B1(n_705), .B2(n_710), .C(n_715), .Y(n_704) );
OAI221xp5_ASAP7_75t_SL g747 ( .A1(n_54), .A2(n_102), .B1(n_748), .B2(n_749), .C(n_751), .Y(n_747) );
INVx1_ASAP7_75t_L g981 ( .A(n_56), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_57), .A2(n_174), .B1(n_830), .B2(n_831), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_57), .A2(n_174), .B1(n_890), .B2(n_892), .Y(n_889) );
INVxp33_ASAP7_75t_L g1040 ( .A(n_58), .Y(n_1040) );
INVx1_ASAP7_75t_L g543 ( .A(n_60), .Y(n_543) );
INVx1_ASAP7_75t_L g676 ( .A(n_61), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_62), .A2(n_135), .B1(n_549), .B2(n_552), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g566 ( .A1(n_62), .A2(n_188), .B1(n_567), .B2(n_568), .C(n_571), .Y(n_566) );
CKINVDCx14_ASAP7_75t_R g1551 ( .A(n_63), .Y(n_1551) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_64), .A2(n_179), .B1(n_384), .B2(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_64), .A2(n_179), .B1(n_486), .B2(n_488), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g1082 ( .A1(n_65), .A2(n_125), .B1(n_604), .B2(n_1002), .C(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1117 ( .A(n_65), .Y(n_1117) );
INVx1_ASAP7_75t_L g958 ( .A(n_66), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g1731 ( .A1(n_67), .A2(n_123), .B1(n_486), .B2(n_1333), .Y(n_1731) );
AOI21xp33_ASAP7_75t_L g1400 ( .A1(n_68), .A2(n_904), .B(n_1315), .Y(n_1400) );
INVxp33_ASAP7_75t_L g1421 ( .A(n_68), .Y(n_1421) );
XOR2x2_ASAP7_75t_L g780 ( .A(n_69), .B(n_781), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g1487 ( .A1(n_70), .A2(n_183), .B1(n_1449), .B2(n_1488), .Y(n_1487) );
INVxp33_ASAP7_75t_L g966 ( .A(n_71), .Y(n_966) );
AOI21xp33_ASAP7_75t_L g998 ( .A1(n_71), .A2(n_591), .B(n_999), .Y(n_998) );
INVxp33_ASAP7_75t_L g799 ( .A(n_72), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g1726 ( .A1(n_73), .A2(n_132), .B1(n_1110), .B2(n_1333), .Y(n_1726) );
AOI22xp33_ASAP7_75t_L g1735 ( .A1(n_73), .A2(n_132), .B1(n_755), .B2(n_916), .Y(n_1735) );
INVxp33_ASAP7_75t_L g967 ( .A(n_74), .Y(n_967) );
XNOR2x2_ASAP7_75t_L g612 ( .A(n_75), .B(n_613), .Y(n_612) );
INVxp33_ASAP7_75t_L g1247 ( .A(n_76), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_76), .A2(n_236), .B1(n_1281), .B2(n_1282), .Y(n_1280) );
INVx1_ASAP7_75t_L g530 ( .A(n_77), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g1395 ( .A(n_78), .Y(n_1395) );
CKINVDCx5p33_ASAP7_75t_R g1141 ( .A(n_79), .Y(n_1141) );
AOI221xp5_ASAP7_75t_L g901 ( .A1(n_80), .A2(n_298), .B1(n_902), .B2(n_903), .C(n_904), .Y(n_901) );
INVxp33_ASAP7_75t_L g929 ( .A(n_80), .Y(n_929) );
INVxp33_ASAP7_75t_L g1029 ( .A(n_81), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_81), .A2(n_311), .B1(n_907), .B2(n_1057), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_82), .A2(n_158), .B1(n_490), .B2(n_1133), .Y(n_1132) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_82), .A2(n_158), .B1(n_581), .B2(n_1164), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_83), .A2(n_207), .B1(n_570), .B2(n_996), .Y(n_1087) );
INVxp33_ASAP7_75t_SL g435 ( .A(n_84), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_84), .A2(n_294), .B1(n_488), .B2(n_492), .Y(n_496) );
CKINVDCx14_ASAP7_75t_R g1479 ( .A(n_85), .Y(n_1479) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_86), .A2(n_252), .B1(n_916), .B2(n_917), .Y(n_915) );
INVxp67_ASAP7_75t_SL g949 ( .A(n_86), .Y(n_949) );
INVx1_ASAP7_75t_L g1385 ( .A(n_87), .Y(n_1385) );
AOI22xp33_ASAP7_75t_SL g905 ( .A1(n_88), .A2(n_198), .B1(n_906), .B2(n_907), .Y(n_905) );
INVxp33_ASAP7_75t_SL g932 ( .A(n_88), .Y(n_932) );
OR2x2_ASAP7_75t_L g345 ( .A(n_89), .B(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g349 ( .A(n_89), .Y(n_349) );
BUFx2_ASAP7_75t_L g444 ( .A(n_89), .Y(n_444) );
INVx1_ASAP7_75t_L g454 ( .A(n_89), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g1727 ( .A1(n_90), .A2(n_210), .B1(n_493), .B2(n_1728), .Y(n_1727) );
AOI22xp33_ASAP7_75t_L g1733 ( .A1(n_90), .A2(n_210), .B1(n_1282), .B2(n_1734), .Y(n_1733) );
AOI221xp5_ASAP7_75t_L g1222 ( .A1(n_91), .A2(n_255), .B1(n_450), .B2(n_536), .C(n_1128), .Y(n_1222) );
INVx1_ASAP7_75t_L g1235 ( .A(n_91), .Y(n_1235) );
AOI22xp33_ASAP7_75t_SL g1134 ( .A1(n_92), .A2(n_101), .B1(n_1127), .B2(n_1128), .Y(n_1134) );
INVx1_ASAP7_75t_L g1162 ( .A(n_92), .Y(n_1162) );
INVxp33_ASAP7_75t_L g1251 ( .A(n_93), .Y(n_1251) );
CKINVDCx5p33_ASAP7_75t_R g1392 ( .A(n_94), .Y(n_1392) );
AOI221xp5_ASAP7_75t_L g1403 ( .A1(n_95), .A2(n_202), .B1(n_1404), .B2(n_1406), .C(n_1409), .Y(n_1403) );
INVxp67_ASAP7_75t_SL g1431 ( .A(n_95), .Y(n_1431) );
INVx1_ASAP7_75t_L g731 ( .A(n_96), .Y(n_731) );
XOR2x2_ASAP7_75t_L g1074 ( .A(n_97), .B(n_1075), .Y(n_1074) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_99), .Y(n_1226) );
INVxp67_ASAP7_75t_SL g977 ( .A(n_100), .Y(n_977) );
AOI221xp5_ASAP7_75t_L g1006 ( .A1(n_100), .A2(n_259), .B1(n_1007), .B2(n_1008), .C(n_1009), .Y(n_1006) );
NOR2xp33_ASAP7_75t_L g1146 ( .A(n_101), .B(n_434), .Y(n_1146) );
CKINVDCx5p33_ASAP7_75t_R g743 ( .A(n_103), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_104), .A2(n_227), .B1(n_627), .B2(n_820), .Y(n_1093) );
OAI211xp5_ASAP7_75t_L g1095 ( .A1(n_104), .A2(n_1096), .B(n_1098), .C(n_1100), .Y(n_1095) );
INVx1_ASAP7_75t_L g1185 ( .A(n_105), .Y(n_1185) );
AOI221xp5_ASAP7_75t_L g1213 ( .A1(n_105), .A2(n_118), .B1(n_459), .B2(n_1131), .C(n_1214), .Y(n_1213) );
OAI22xp33_ASAP7_75t_SL g643 ( .A1(n_106), .A2(n_134), .B1(n_572), .B2(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g681 ( .A(n_106), .Y(n_681) );
INVx1_ASAP7_75t_L g1267 ( .A(n_107), .Y(n_1267) );
XNOR2x1_ASAP7_75t_L g1020 ( .A(n_108), .B(n_1021), .Y(n_1020) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_110), .Y(n_630) );
INVx1_ASAP7_75t_L g596 ( .A(n_111), .Y(n_596) );
OAI222xp33_ASAP7_75t_L g1772 ( .A1(n_112), .A2(n_171), .B1(n_289), .B2(n_1160), .C1(n_1285), .C2(n_1773), .Y(n_1772) );
INVx1_ASAP7_75t_L g1783 ( .A(n_112), .Y(n_1783) );
OAI22xp33_ASAP7_75t_L g1079 ( .A1(n_114), .A2(n_266), .B1(n_385), .B2(n_604), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_114), .A2(n_163), .B1(n_859), .B2(n_1110), .Y(n_1109) );
AOI221xp5_ASAP7_75t_L g1320 ( .A1(n_115), .A2(n_262), .B1(n_578), .B2(n_638), .C(n_1281), .Y(n_1320) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_115), .A2(n_193), .B1(n_493), .B2(n_952), .Y(n_1334) );
AOI21xp5_ASAP7_75t_L g1094 ( .A1(n_116), .A2(n_591), .B(n_999), .Y(n_1094) );
INVx1_ASAP7_75t_L g1101 ( .A(n_116), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_117), .A2(n_163), .B1(n_599), .B2(n_644), .Y(n_1078) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_117), .A2(n_266), .B1(n_468), .B2(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1205 ( .A(n_118), .Y(n_1205) );
OAI221xp5_ASAP7_75t_L g1357 ( .A1(n_119), .A2(n_155), .B1(n_712), .B2(n_934), .C(n_1031), .Y(n_1357) );
OAI22xp33_ASAP7_75t_L g1384 ( .A1(n_119), .A2(n_155), .B1(n_1284), .B2(n_1285), .Y(n_1384) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_120), .A2(n_260), .B1(n_389), .B2(n_415), .C(n_419), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_120), .A2(n_260), .B1(n_492), .B2(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g533 ( .A(n_121), .Y(n_533) );
XNOR2xp5_ASAP7_75t_L g1242 ( .A(n_122), .B(n_1243), .Y(n_1242) );
INVx1_ASAP7_75t_L g1690 ( .A(n_123), .Y(n_1690) );
CKINVDCx5p33_ASAP7_75t_R g1085 ( .A(n_124), .Y(n_1085) );
INVx1_ASAP7_75t_L g1099 ( .A(n_125), .Y(n_1099) );
AOI22xp5_ASAP7_75t_SL g1506 ( .A1(n_126), .A2(n_147), .B1(n_1449), .B2(n_1457), .Y(n_1506) );
AOI221xp5_ASAP7_75t_L g1760 ( .A1(n_127), .A2(n_258), .B1(n_416), .B2(n_578), .C(n_1761), .Y(n_1760) );
INVx1_ASAP7_75t_L g1792 ( .A(n_127), .Y(n_1792) );
INVx1_ASAP7_75t_L g694 ( .A(n_128), .Y(n_694) );
INVxp33_ASAP7_75t_SL g432 ( .A(n_129), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_129), .A2(n_244), .B1(n_486), .B2(n_494), .Y(n_497) );
INVx1_ASAP7_75t_L g1045 ( .A(n_130), .Y(n_1045) );
INVx1_ASAP7_75t_L g1453 ( .A(n_131), .Y(n_1453) );
CKINVDCx5p33_ASAP7_75t_R g989 ( .A(n_133), .Y(n_989) );
INVx1_ASAP7_75t_L g671 ( .A(n_134), .Y(n_671) );
INVx1_ASAP7_75t_L g574 ( .A(n_135), .Y(n_574) );
INVx1_ASAP7_75t_L g1149 ( .A(n_136), .Y(n_1149) );
INVx1_ASAP7_75t_L g964 ( .A(n_137), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_137), .B(n_399), .Y(n_1000) );
INVx1_ASAP7_75t_L g734 ( .A(n_138), .Y(n_734) );
CKINVDCx16_ASAP7_75t_R g1500 ( .A(n_139), .Y(n_1500) );
INVx1_ASAP7_75t_L g811 ( .A(n_140), .Y(n_811) );
INVxp67_ASAP7_75t_L g1265 ( .A(n_141), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_141), .A2(n_176), .B1(n_384), .B2(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1047 ( .A(n_143), .Y(n_1047) );
INVx1_ASAP7_75t_L g1454 ( .A(n_144), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_144), .B(n_1452), .Y(n_1459) );
AOI22xp33_ASAP7_75t_SL g818 ( .A1(n_145), .A2(n_168), .B1(n_819), .B2(n_821), .Y(n_818) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_145), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g1321 ( .A1(n_146), .A2(n_193), .B1(n_756), .B2(n_1322), .Y(n_1321) );
AOI22xp33_ASAP7_75t_SL g1332 ( .A1(n_146), .A2(n_262), .B1(n_1110), .B2(n_1333), .Y(n_1332) );
AOI21xp5_ASAP7_75t_L g1314 ( .A1(n_148), .A2(n_404), .B(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1342 ( .A(n_148), .Y(n_1342) );
INVx1_ASAP7_75t_L g1273 ( .A(n_149), .Y(n_1273) );
INVx2_ASAP7_75t_L g330 ( .A(n_150), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g1181 ( .A(n_151), .Y(n_1181) );
AOI221xp5_ASAP7_75t_L g912 ( .A1(n_152), .A2(n_281), .B1(n_368), .B2(n_913), .C(n_914), .Y(n_912) );
INVxp33_ASAP7_75t_SL g942 ( .A(n_152), .Y(n_942) );
INVx1_ASAP7_75t_L g753 ( .A(n_153), .Y(n_753) );
BUFx3_ASAP7_75t_L g358 ( .A(n_154), .Y(n_358) );
INVx1_ASAP7_75t_L g388 ( .A(n_154), .Y(n_388) );
INVx1_ASAP7_75t_L g790 ( .A(n_157), .Y(n_790) );
INVx1_ASAP7_75t_L g983 ( .A(n_159), .Y(n_983) );
INVxp33_ASAP7_75t_L g1355 ( .A(n_160), .Y(n_1355) );
AOI221xp5_ASAP7_75t_L g1382 ( .A1(n_160), .A2(n_199), .B1(n_416), .B2(n_591), .C(n_999), .Y(n_1382) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_161), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_162), .A2(n_269), .B1(n_673), .B2(n_1108), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_162), .A2(n_269), .B1(n_626), .B2(n_819), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1736 ( .A1(n_164), .A2(n_205), .B1(n_416), .B2(n_1737), .Y(n_1736) );
INVxp67_ASAP7_75t_L g719 ( .A(n_165), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_165), .A2(n_278), .B1(n_423), .B2(n_771), .Y(n_770) );
OAI221xp5_ASAP7_75t_SL g1396 ( .A1(n_166), .A2(n_297), .B1(n_379), .B2(n_1284), .C(n_1397), .Y(n_1396) );
OAI221xp5_ASAP7_75t_L g1423 ( .A1(n_166), .A2(n_297), .B1(n_705), .B2(n_712), .C(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g701 ( .A(n_167), .Y(n_701) );
INVxp67_ASAP7_75t_SL g881 ( .A(n_168), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g839 ( .A(n_170), .Y(n_839) );
INVx1_ASAP7_75t_L g1777 ( .A(n_171), .Y(n_1777) );
INVxp33_ASAP7_75t_SL g524 ( .A(n_172), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_172), .A2(n_216), .B1(n_567), .B2(n_580), .C(n_583), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g1759 ( .A1(n_173), .A2(n_250), .B1(n_830), .B2(n_1322), .Y(n_1759) );
INVx1_ASAP7_75t_L g1782 ( .A(n_173), .Y(n_1782) );
INVxp67_ASAP7_75t_L g1038 ( .A(n_175), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_175), .A2(n_226), .B1(n_903), .B2(n_907), .Y(n_1062) );
INVxp33_ASAP7_75t_L g1259 ( .A(n_176), .Y(n_1259) );
INVx1_ASAP7_75t_L g1414 ( .A(n_177), .Y(n_1414) );
INVx1_ASAP7_75t_L g353 ( .A(n_178), .Y(n_353) );
INVx1_ASAP7_75t_L g406 ( .A(n_178), .Y(n_406) );
INVxp33_ASAP7_75t_SL g1352 ( .A(n_180), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_180), .A2(n_187), .B1(n_389), .B2(n_601), .Y(n_1383) );
INVx1_ASAP7_75t_L g1194 ( .A(n_181), .Y(n_1194) );
OAI221xp5_ASAP7_75t_L g1217 ( .A1(n_181), .A2(n_206), .B1(n_867), .B2(n_1218), .C(n_1220), .Y(n_1217) );
INVx1_ASAP7_75t_L g980 ( .A(n_182), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g1549 ( .A(n_184), .Y(n_1549) );
INVx1_ASAP7_75t_L g908 ( .A(n_185), .Y(n_908) );
INVx1_ASAP7_75t_L g1364 ( .A(n_186), .Y(n_1364) );
INVxp33_ASAP7_75t_SL g1356 ( .A(n_187), .Y(n_1356) );
INVx1_ASAP7_75t_L g547 ( .A(n_188), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_189), .Y(n_1090) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_190), .A2(n_267), .B1(n_624), .B2(n_626), .C(n_628), .Y(n_623) );
INVx1_ASAP7_75t_L g686 ( .A(n_190), .Y(n_686) );
INVx1_ASAP7_75t_L g1042 ( .A(n_191), .Y(n_1042) );
AOI22xp33_ASAP7_75t_SL g826 ( .A1(n_192), .A2(n_241), .B1(n_821), .B2(n_827), .Y(n_826) );
OAI211xp5_ASAP7_75t_SL g849 ( .A1(n_192), .A2(n_850), .B(n_854), .C(n_863), .Y(n_849) );
INVx1_ASAP7_75t_L g1345 ( .A(n_194), .Y(n_1345) );
AOI221xp5_ASAP7_75t_L g1758 ( .A1(n_196), .A2(n_264), .B1(n_424), .B2(n_904), .C(n_1691), .Y(n_1758) );
INVx1_ASAP7_75t_L g1780 ( .A(n_196), .Y(n_1780) );
CKINVDCx14_ASAP7_75t_R g1481 ( .A(n_197), .Y(n_1481) );
INVxp33_ASAP7_75t_L g927 ( .A(n_198), .Y(n_927) );
INVxp33_ASAP7_75t_L g1353 ( .A(n_199), .Y(n_1353) );
INVx1_ASAP7_75t_L g1050 ( .A(n_200), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g1123 ( .A(n_201), .Y(n_1123) );
INVx1_ASAP7_75t_L g1429 ( .A(n_202), .Y(n_1429) );
INVx1_ASAP7_75t_L g1720 ( .A(n_203), .Y(n_1720) );
AOI22xp33_ASAP7_75t_L g1410 ( .A1(n_204), .A2(n_254), .B1(n_616), .B2(n_1411), .Y(n_1410) );
INVx1_ASAP7_75t_L g1428 ( .A(n_204), .Y(n_1428) );
INVx1_ASAP7_75t_L g1199 ( .A(n_206), .Y(n_1199) );
INVx1_ASAP7_75t_L g1114 ( .A(n_207), .Y(n_1114) );
INVxp67_ASAP7_75t_L g1262 ( .A(n_208), .Y(n_1262) );
AOI221xp5_ASAP7_75t_L g1289 ( .A1(n_208), .A2(n_303), .B1(n_755), .B2(n_914), .C(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1144 ( .A(n_211), .Y(n_1144) );
OAI211xp5_ASAP7_75t_L g1159 ( .A1(n_211), .A2(n_1160), .B(n_1161), .C(n_1165), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_212), .A2(n_222), .B1(n_582), .B2(n_627), .Y(n_1399) );
INVxp33_ASAP7_75t_L g1422 ( .A(n_212), .Y(n_1422) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_213), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g1052 ( .A(n_214), .Y(n_1052) );
INVxp33_ASAP7_75t_SL g528 ( .A(n_216), .Y(n_528) );
INVx1_ASAP7_75t_L g732 ( .A(n_217), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g1497 ( .A(n_218), .Y(n_1497) );
BUFx3_ASAP7_75t_L g360 ( .A(n_219), .Y(n_360) );
INVx1_ASAP7_75t_L g370 ( .A(n_219), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_220), .Y(n_620) );
AO221x2_ASAP7_75t_L g1546 ( .A1(n_221), .A2(n_283), .B1(n_1490), .B2(n_1547), .C(n_1548), .Y(n_1546) );
INVxp33_ASAP7_75t_L g1419 ( .A(n_222), .Y(n_1419) );
AOI22xp5_ASAP7_75t_L g1470 ( .A1(n_223), .A2(n_224), .B1(n_1465), .B2(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1439 ( .A(n_224), .Y(n_1439) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_225), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_225), .B(n_286), .Y(n_346) );
AND2x2_ASAP7_75t_L g455 ( .A(n_225), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g505 ( .A(n_225), .Y(n_505) );
INVxp67_ASAP7_75t_L g1036 ( .A(n_226), .Y(n_1036) );
INVx1_ASAP7_75t_L g1103 ( .A(n_227), .Y(n_1103) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_228), .A2(n_399), .B(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g472 ( .A(n_228), .Y(n_472) );
INVx1_ASAP7_75t_L g921 ( .A(n_229), .Y(n_921) );
INVx1_ASAP7_75t_L g595 ( .A(n_230), .Y(n_595) );
INVx2_ASAP7_75t_L g355 ( .A(n_231), .Y(n_355) );
OR2x2_ASAP7_75t_L g372 ( .A(n_231), .B(n_353), .Y(n_372) );
INVx1_ASAP7_75t_L g1340 ( .A(n_232), .Y(n_1340) );
INVxp67_ASAP7_75t_L g724 ( .A(n_233), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_233), .A2(n_277), .B1(n_764), .B2(n_765), .C(n_769), .Y(n_763) );
INVx1_ASAP7_75t_L g1798 ( .A(n_234), .Y(n_1798) );
INVx1_ASAP7_75t_L g1367 ( .A(n_235), .Y(n_1367) );
INVxp33_ASAP7_75t_SL g1252 ( .A(n_236), .Y(n_1252) );
INVx1_ASAP7_75t_L g1326 ( .A(n_237), .Y(n_1326) );
INVx1_ASAP7_75t_L g922 ( .A(n_238), .Y(n_922) );
INVx1_ASAP7_75t_L g1229 ( .A(n_239), .Y(n_1229) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_239), .A2(n_263), .B1(n_819), .B2(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1402 ( .A(n_240), .Y(n_1402) );
OAI221xp5_ASAP7_75t_L g868 ( .A1(n_241), .A2(n_869), .B1(n_871), .B2(n_878), .C(n_888), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g1762 ( .A1(n_242), .A2(n_261), .B1(n_907), .B2(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g1790 ( .A(n_242), .Y(n_1790) );
AOI22xp5_ASAP7_75t_SL g1460 ( .A1(n_243), .A2(n_247), .B1(n_1461), .B2(n_1465), .Y(n_1460) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_244), .Y(n_413) );
INVx1_ASAP7_75t_L g737 ( .A(n_245), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_246), .A2(n_251), .B1(n_384), .B2(n_389), .C(n_390), .Y(n_383) );
INVxp33_ASAP7_75t_L g465 ( .A(n_246), .Y(n_465) );
XNOR2xp5_ASAP7_75t_L g1171 ( .A(n_247), .B(n_1172), .Y(n_1171) );
INVx1_ASAP7_75t_L g956 ( .A(n_248), .Y(n_956) );
INVx1_ASAP7_75t_L g1137 ( .A(n_249), .Y(n_1137) );
AOI21xp5_ASAP7_75t_L g1156 ( .A1(n_249), .A2(n_570), .B(n_632), .Y(n_1156) );
INVx1_ASAP7_75t_L g1779 ( .A(n_250), .Y(n_1779) );
INVxp33_ASAP7_75t_L g939 ( .A(n_252), .Y(n_939) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_253), .Y(n_619) );
INVx1_ASAP7_75t_L g1434 ( .A(n_254), .Y(n_1434) );
INVx1_ASAP7_75t_L g1236 ( .A(n_255), .Y(n_1236) );
INVx1_ASAP7_75t_L g985 ( .A(n_256), .Y(n_985) );
INVx1_ASAP7_75t_L g1140 ( .A(n_257), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1786 ( .A1(n_258), .A2(n_261), .B1(n_1728), .B2(n_1787), .C(n_1789), .Y(n_1786) );
INVxp33_ASAP7_75t_L g972 ( .A(n_259), .Y(n_972) );
INVx1_ASAP7_75t_L g1228 ( .A(n_263), .Y(n_1228) );
INVx1_ASAP7_75t_L g1785 ( .A(n_264), .Y(n_1785) );
CKINVDCx5p33_ASAP7_75t_R g1766 ( .A(n_265), .Y(n_1766) );
INVx1_ASAP7_75t_L g688 ( .A(n_267), .Y(n_688) );
INVx1_ASAP7_75t_L g923 ( .A(n_268), .Y(n_923) );
INVx1_ASAP7_75t_L g1324 ( .A(n_270), .Y(n_1324) );
INVx1_ASAP7_75t_L g1398 ( .A(n_271), .Y(n_1398) );
INVx1_ASAP7_75t_L g1347 ( .A(n_272), .Y(n_1347) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_273), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_273), .B(n_318), .Y(n_1456) );
AND3x2_ASAP7_75t_L g1464 ( .A(n_273), .B(n_318), .C(n_1453), .Y(n_1464) );
INVx2_ASAP7_75t_L g331 ( .A(n_275), .Y(n_331) );
XNOR2x2_ASAP7_75t_L g520 ( .A(n_276), .B(n_521), .Y(n_520) );
INVxp67_ASAP7_75t_SL g728 ( .A(n_277), .Y(n_728) );
INVxp33_ASAP7_75t_SL g721 ( .A(n_278), .Y(n_721) );
INVx1_ASAP7_75t_L g1305 ( .A(n_279), .Y(n_1305) );
CKINVDCx5p33_ASAP7_75t_R g1694 ( .A(n_280), .Y(n_1694) );
INVxp67_ASAP7_75t_SL g945 ( .A(n_281), .Y(n_945) );
INVx1_ASAP7_75t_L g526 ( .A(n_282), .Y(n_526) );
INVx1_ASAP7_75t_L g1370 ( .A(n_284), .Y(n_1370) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_285), .Y(n_652) );
INVx1_ASAP7_75t_L g333 ( .A(n_286), .Y(n_333) );
INVx2_ASAP7_75t_L g456 ( .A(n_286), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_287), .Y(n_650) );
INVxp67_ASAP7_75t_SL g1363 ( .A(n_288), .Y(n_1363) );
INVx1_ASAP7_75t_L g1776 ( .A(n_289), .Y(n_1776) );
INVxp33_ASAP7_75t_L g1028 ( .A(n_290), .Y(n_1028) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_290), .A2(n_292), .B1(n_424), .B2(n_902), .C(n_904), .Y(n_1055) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_291), .A2(n_304), .B1(n_603), .B2(n_604), .Y(n_602) );
INVxp33_ASAP7_75t_L g1026 ( .A(n_292), .Y(n_1026) );
INVxp67_ASAP7_75t_SL g887 ( .A(n_293), .Y(n_887) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_294), .Y(n_364) );
INVx1_ASAP7_75t_L g1368 ( .A(n_295), .Y(n_1368) );
INVxp67_ASAP7_75t_SL g511 ( .A(n_296), .Y(n_511) );
INVxp33_ASAP7_75t_L g931 ( .A(n_298), .Y(n_931) );
INVx1_ASAP7_75t_L g669 ( .A(n_300), .Y(n_669) );
INVx1_ASAP7_75t_L g1295 ( .A(n_301), .Y(n_1295) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_302), .Y(n_361) );
INVxp33_ASAP7_75t_L g1260 ( .A(n_303), .Y(n_1260) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_304), .Y(n_559) );
INVx1_ASAP7_75t_L g1202 ( .A(n_305), .Y(n_1202) );
AOI21xp5_ASAP7_75t_L g1216 ( .A1(n_305), .A2(n_861), .B(n_1127), .Y(n_1216) );
INVx1_ASAP7_75t_L g1413 ( .A(n_306), .Y(n_1413) );
INVx1_ASAP7_75t_L g1371 ( .A(n_307), .Y(n_1371) );
INVxp33_ASAP7_75t_SL g700 ( .A(n_308), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g1313 ( .A(n_309), .Y(n_1313) );
INVx1_ASAP7_75t_L g1329 ( .A(n_310), .Y(n_1329) );
INVxp33_ASAP7_75t_L g1025 ( .A(n_311), .Y(n_1025) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_334), .B(n_1441), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_321), .Y(n_315) );
AND2x4_ASAP7_75t_L g1747 ( .A(n_316), .B(n_322), .Y(n_1747) );
NOR2xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_SL g1751 ( .A(n_317), .Y(n_1751) );
NAND2xp5_ASAP7_75t_L g1804 ( .A(n_317), .B(n_319), .Y(n_1804) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_319), .B(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x6_ASAP7_75t_L g1724 ( .A(n_324), .B(n_349), .Y(n_1724) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g484 ( .A(n_325), .B(n_333), .Y(n_484) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g536 ( .A(n_326), .B(n_537), .Y(n_536) );
OR2x6_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .Y(n_327) );
OR2x2_ASAP7_75t_L g344 ( .A(n_328), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g659 ( .A(n_328), .Y(n_659) );
INVx2_ASAP7_75t_SL g874 ( .A(n_328), .Y(n_874) );
BUFx6f_ASAP7_75t_L g941 ( .A(n_328), .Y(n_941) );
INVx2_ASAP7_75t_SL g975 ( .A(n_328), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_328), .A2(n_679), .B1(n_1085), .B2(n_1114), .Y(n_1113) );
OR2x6_ASAP7_75t_L g1712 ( .A(n_328), .B(n_1713), .Y(n_1712) );
BUFx2_ASAP7_75t_L g1791 ( .A(n_328), .Y(n_1791) );
OAI22xp33_ASAP7_75t_L g1797 ( .A1(n_328), .A2(n_679), .B1(n_1766), .B2(n_1798), .Y(n_1797) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
AND2x2_ASAP7_75t_L g452 ( .A(n_330), .B(n_331), .Y(n_452) );
INVx2_ASAP7_75t_L g461 ( .A(n_330), .Y(n_461) );
AND2x4_ASAP7_75t_L g470 ( .A(n_330), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g477 ( .A(n_330), .Y(n_477) );
INVx1_ASAP7_75t_L g515 ( .A(n_330), .Y(n_515) );
INVx1_ASAP7_75t_L g463 ( .A(n_331), .Y(n_463) );
INVx2_ASAP7_75t_L g471 ( .A(n_331), .Y(n_471) );
INVx1_ASAP7_75t_L g509 ( .A(n_331), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_331), .B(n_461), .Y(n_542) );
INVx1_ASAP7_75t_L g664 ( .A(n_331), .Y(n_664) );
AND2x4_ASAP7_75t_L g1709 ( .A(n_332), .B(n_509), .Y(n_1709) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g1710 ( .A(n_333), .B(n_514), .Y(n_1710) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_1068), .B1(n_1069), .B2(n_1440), .Y(n_334) );
INVx3_ASAP7_75t_L g1440 ( .A(n_335), .Y(n_1440) );
AO22x2_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_777), .B1(n_1066), .B2(n_1067), .Y(n_335) );
INVx1_ASAP7_75t_L g1067 ( .A(n_336), .Y(n_1067) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_692), .B1(n_693), .B2(n_776), .Y(n_336) );
INVx2_ASAP7_75t_L g776 ( .A(n_337), .Y(n_776) );
AO22x2_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_518), .B1(n_519), .B2(n_691), .Y(n_337) );
INVx2_ASAP7_75t_SL g691 ( .A(n_338), .Y(n_691) );
XNOR2x1_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_339), .A2(n_1491), .B1(n_1502), .B2(n_1503), .Y(n_1501) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_445), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_361), .B(n_362), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g1372 ( .A1(n_342), .A2(n_440), .B1(n_1373), .B2(n_1385), .Y(n_1372) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx5_ASAP7_75t_L g742 ( .A(n_343), .Y(n_742) );
INVx1_ASAP7_75t_L g988 ( .A(n_343), .Y(n_988) );
INVx2_ASAP7_75t_L g1296 ( .A(n_343), .Y(n_1296) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_347), .Y(n_343) );
INVx2_ASAP7_75t_L g531 ( .A(n_344), .Y(n_531) );
INVx3_ASAP7_75t_L g510 ( .A(n_345), .Y(n_510) );
INVx1_ASAP7_75t_L g846 ( .A(n_346), .Y(n_846) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x6_ASAP7_75t_L g840 ( .A(n_348), .B(n_841), .Y(n_840) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x4_ASAP7_75t_L g833 ( .A(n_349), .B(n_405), .Y(n_833) );
INVx2_ASAP7_75t_L g1160 ( .A(n_350), .Y(n_1160) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_356), .Y(n_350) );
AND2x4_ASAP7_75t_L g375 ( .A(n_351), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g380 ( .A(n_351), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g430 ( .A(n_351), .Y(n_430) );
BUFx2_ASAP7_75t_L g593 ( .A(n_351), .Y(n_593) );
AND2x4_ASAP7_75t_L g649 ( .A(n_351), .B(n_376), .Y(n_649) );
AND2x4_ASAP7_75t_L g651 ( .A(n_351), .B(n_381), .Y(n_651) );
NAND2x1p5_ASAP7_75t_L g810 ( .A(n_351), .B(n_502), .Y(n_810) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_351), .B(n_381), .Y(n_1308) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g405 ( .A(n_354), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g421 ( .A(n_355), .B(n_406), .Y(n_421) );
INVx1_ASAP7_75t_L g1179 ( .A(n_355), .Y(n_1179) );
HB1xp67_ASAP7_75t_L g1184 ( .A(n_355), .Y(n_1184) );
INVx1_ASAP7_75t_L g1188 ( .A(n_355), .Y(n_1188) );
INVx6_ASAP7_75t_L g426 ( .A(n_356), .Y(n_426) );
BUFx2_ASAP7_75t_L g591 ( .A(n_356), .Y(n_591) );
INVx2_ASAP7_75t_L g798 ( .A(n_356), .Y(n_798) );
AND2x4_ASAP7_75t_L g1182 ( .A(n_356), .B(n_1183), .Y(n_1182) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g382 ( .A(n_357), .Y(n_382) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g369 ( .A(n_358), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g412 ( .A(n_358), .B(n_360), .Y(n_412) );
INVx1_ASAP7_75t_L g378 ( .A(n_359), .Y(n_378) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g387 ( .A(n_360), .B(n_388), .Y(n_387) );
AOI31xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_407), .A3(n_431), .B(n_439), .Y(n_362) );
AOI211xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_365), .B(n_373), .C(n_383), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g991 ( .A1(n_365), .A2(n_980), .B(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_367), .Y(n_746) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_367), .A2(n_901), .B1(n_905), .B2(n_908), .C(n_909), .Y(n_900) );
AOI221xp5_ASAP7_75t_L g1054 ( .A1(n_367), .A2(n_1042), .B1(n_1055), .B2(n_1056), .C(n_1058), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1294 ( .A1(n_367), .A2(n_433), .B1(n_1267), .B2(n_1272), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_367), .A2(n_433), .B1(n_1324), .B2(n_1325), .Y(n_1323) );
AOI21xp5_ASAP7_75t_L g1394 ( .A1(n_367), .A2(n_1395), .B(n_1396), .Y(n_1394) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_371), .Y(n_367) );
INVx2_ASAP7_75t_SL g752 ( .A(n_368), .Y(n_752) );
BUFx3_ASAP7_75t_L g906 ( .A(n_368), .Y(n_906) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g389 ( .A(n_369), .Y(n_389) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_369), .Y(n_576) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_369), .Y(n_582) );
INVx2_ASAP7_75t_SL g625 ( .A(n_369), .Y(n_625) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_369), .Y(n_645) );
BUFx3_ASAP7_75t_L g820 ( .A(n_369), .Y(n_820) );
BUFx2_ASAP7_75t_L g995 ( .A(n_369), .Y(n_995) );
AND2x6_ASAP7_75t_L g1206 ( .A(n_369), .B(n_1178), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1290 ( .A(n_369), .Y(n_1290) );
HB1xp67_ASAP7_75t_L g1761 ( .A(n_369), .Y(n_1761) );
INVx1_ASAP7_75t_L g396 ( .A(n_370), .Y(n_396) );
AND2x4_ASAP7_75t_L g410 ( .A(n_371), .B(n_411), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g597 ( .A1(n_371), .A2(n_598), .B(n_602), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g640 ( .A1(n_371), .A2(n_641), .B(n_643), .Y(n_640) );
OAI21xp5_ASAP7_75t_L g1077 ( .A1(n_371), .A2(n_1078), .B(n_1079), .Y(n_1077) );
A2O1A1Ixp33_ASAP7_75t_L g1161 ( .A1(n_371), .A2(n_902), .B(n_1162), .C(n_1163), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_371), .B(n_645), .Y(n_1377) );
AOI221xp5_ASAP7_75t_L g1765 ( .A1(n_371), .A2(n_433), .B1(n_1766), .B2(n_1767), .C(n_1772), .Y(n_1765) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g434 ( .A(n_372), .B(n_394), .Y(n_434) );
OR2x2_ASAP7_75t_L g437 ( .A(n_372), .B(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g789 ( .A(n_372), .B(n_454), .Y(n_789) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_375), .A2(n_380), .B1(n_595), .B2(n_596), .Y(n_594) );
INVx2_ASAP7_75t_SL g748 ( .A(n_375), .Y(n_748) );
INVx2_ASAP7_75t_SL g910 ( .A(n_375), .Y(n_910) );
INVxp67_ASAP7_75t_L g1002 ( .A(n_376), .Y(n_1002) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g808 ( .A(n_377), .Y(n_808) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g1198 ( .A(n_378), .Y(n_1198) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g750 ( .A(n_381), .Y(n_750) );
INVx1_ASAP7_75t_L g1083 ( .A(n_381), .Y(n_1083) );
BUFx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x6_ASAP7_75t_L g1200 ( .A(n_382), .B(n_1179), .Y(n_1200) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g751 ( .A1(n_385), .A2(n_701), .B1(n_752), .B2(n_753), .C(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g1322 ( .A(n_385), .Y(n_1322) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_386), .Y(n_567) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_386), .Y(n_616) );
INVx1_ASAP7_75t_L g772 ( .A(n_386), .Y(n_772) );
INVx1_ASAP7_75t_L g1014 ( .A(n_386), .Y(n_1014) );
AND2x6_ASAP7_75t_L g1186 ( .A(n_386), .B(n_1187), .Y(n_1186) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_387), .Y(n_627) );
INVx1_ASAP7_75t_L g793 ( .A(n_387), .Y(n_793) );
INVx1_ASAP7_75t_L g918 ( .A(n_387), .Y(n_918) );
INVx1_ASAP7_75t_L g395 ( .A(n_388), .Y(n_395) );
OAI21xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_397), .B(n_398), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g1239 ( .A1(n_391), .A2(n_1091), .B1(n_1225), .B2(n_1226), .C(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g599 ( .A(n_393), .Y(n_599) );
INVx2_ASAP7_75t_L g1234 ( .A(n_393), .Y(n_1234) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g587 ( .A(n_394), .Y(n_587) );
OR2x2_ASAP7_75t_L g1701 ( .A(n_394), .B(n_1702), .Y(n_1701) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
AND2x2_ASAP7_75t_L g402 ( .A(n_395), .B(n_396), .Y(n_402) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g573 ( .A(n_402), .Y(n_573) );
BUFx4f_ASAP7_75t_L g585 ( .A(n_402), .Y(n_585) );
INVx2_ASAP7_75t_L g802 ( .A(n_402), .Y(n_802) );
INVx1_ASAP7_75t_L g1769 ( .A(n_402), .Y(n_1769) );
BUFx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_405), .Y(n_588) );
INVx2_ASAP7_75t_SL g632 ( .A(n_405), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_405), .Y(n_904) );
INVx1_ASAP7_75t_L g999 ( .A(n_405), .Y(n_999) );
INVx1_ASAP7_75t_L g1208 ( .A(n_406), .Y(n_1208) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_413), .B1(n_414), .B2(n_422), .C(n_427), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_410), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g911 ( .A1(n_410), .A2(n_428), .B1(n_912), .B2(n_915), .C(n_919), .Y(n_911) );
INVx1_ASAP7_75t_L g1005 ( .A(n_410), .Y(n_1005) );
INVx1_ASAP7_75t_L g1288 ( .A(n_410), .Y(n_1288) );
INVx2_ASAP7_75t_SL g1318 ( .A(n_410), .Y(n_1318) );
BUFx3_ASAP7_75t_L g755 ( .A(n_411), .Y(n_755) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_411), .Y(n_822) );
BUFx4f_ASAP7_75t_L g902 ( .A(n_411), .Y(n_902) );
AND2x4_ASAP7_75t_L g1158 ( .A(n_411), .B(n_593), .Y(n_1158) );
INVx1_ASAP7_75t_L g1279 ( .A(n_411), .Y(n_1279) );
INVx2_ASAP7_75t_SL g1692 ( .A(n_411), .Y(n_1692) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_412), .Y(n_418) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_L g590 ( .A1(n_416), .A2(n_530), .B(n_591), .C(n_592), .Y(n_590) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g428 ( .A(n_417), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g639 ( .A(n_417), .Y(n_639) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g768 ( .A(n_418), .Y(n_768) );
AND2x4_ASAP7_75t_L g1176 ( .A(n_418), .B(n_1177), .Y(n_1176) );
INVx1_ASAP7_75t_L g1408 ( .A(n_418), .Y(n_1408) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g914 ( .A(n_420), .Y(n_914) );
BUFx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_SL g578 ( .A(n_421), .Y(n_578) );
INVx1_ASAP7_75t_L g622 ( .A(n_421), .Y(n_622) );
INVx2_ASAP7_75t_L g817 ( .A(n_421), .Y(n_817) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g757 ( .A(n_425), .Y(n_757) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g570 ( .A(n_426), .Y(n_570) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_426), .Y(n_636) );
INVx1_ASAP7_75t_L g825 ( .A(n_426), .Y(n_825) );
INVx2_ASAP7_75t_SL g1152 ( .A(n_426), .Y(n_1152) );
INVx2_ASAP7_75t_L g1204 ( .A(n_426), .Y(n_1204) );
INVx2_ASAP7_75t_L g1315 ( .A(n_426), .Y(n_1315) );
HB1xp67_ASAP7_75t_L g1764 ( .A(n_426), .Y(n_1764) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g774 ( .A(n_428), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g1003 ( .A1(n_428), .A2(n_985), .B1(n_1004), .B2(n_1006), .C(n_1011), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g1060 ( .A1(n_428), .A2(n_762), .B1(n_1050), .B2(n_1061), .C(n_1062), .Y(n_1060) );
AOI221xp5_ASAP7_75t_L g1286 ( .A1(n_428), .A2(n_1273), .B1(n_1287), .B2(n_1289), .C(n_1291), .Y(n_1286) );
AOI221xp5_ASAP7_75t_L g1316 ( .A1(n_428), .A2(n_1317), .B1(n_1319), .B2(n_1320), .C(n_1321), .Y(n_1316) );
AOI221xp5_ASAP7_75t_L g1378 ( .A1(n_428), .A2(n_1317), .B1(n_1371), .B2(n_1379), .C(n_1380), .Y(n_1378) );
AOI221xp5_ASAP7_75t_L g1401 ( .A1(n_428), .A2(n_762), .B1(n_1402), .B2(n_1403), .C(n_1410), .Y(n_1401) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g749 ( .A(n_430), .B(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_435), .B2(n_436), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_433), .A2(n_436), .B1(n_732), .B2(n_734), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_433), .A2(n_436), .B1(n_921), .B2(n_922), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_433), .A2(n_436), .B1(n_981), .B2(n_983), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_433), .A2(n_436), .B1(n_1045), .B2(n_1047), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g1374 ( .A1(n_433), .A2(n_1367), .B1(n_1370), .B2(n_1375), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1412 ( .A1(n_433), .A2(n_436), .B1(n_1413), .B2(n_1414), .Y(n_1412) );
INVx6_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g1276 ( .A1(n_436), .A2(n_1270), .B1(n_1277), .B2(n_1280), .C(n_1283), .Y(n_1276) );
AOI211xp5_ASAP7_75t_L g1304 ( .A1(n_436), .A2(n_1305), .B(n_1306), .C(n_1309), .Y(n_1304) );
AOI221xp5_ASAP7_75t_L g1381 ( .A1(n_436), .A2(n_1368), .B1(n_1382), .B2(n_1383), .C(n_1384), .Y(n_1381) );
INVx4_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g601 ( .A(n_438), .Y(n_601) );
INVx2_ASAP7_75t_L g997 ( .A(n_438), .Y(n_997) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g1274 ( .A1(n_440), .A2(n_1275), .B1(n_1295), .B2(n_1296), .Y(n_1274) );
INVx5_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI31xp33_ASAP7_75t_L g744 ( .A1(n_441), .A2(n_745), .A3(n_759), .B(n_775), .Y(n_744) );
OAI31xp33_ASAP7_75t_L g848 ( .A1(n_441), .A2(n_849), .A3(n_868), .B(n_889), .Y(n_848) );
AOI31xp33_ASAP7_75t_L g1053 ( .A1(n_441), .A2(n_1054), .A3(n_1060), .B(n_1063), .Y(n_1053) );
AOI221x1_ASAP7_75t_SL g1172 ( .A1(n_441), .A2(n_1173), .B1(n_1207), .B2(n_1209), .C(n_1230), .Y(n_1172) );
BUFx8_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g898 ( .A(n_442), .Y(n_898) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g653 ( .A(n_443), .Y(n_653) );
AND2x4_ASAP7_75t_L g1207 ( .A(n_443), .B(n_1208), .Y(n_1207) );
AND2x4_ASAP7_75t_L g1704 ( .A(n_443), .B(n_1208), .Y(n_1704) );
BUFx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
OR2x6_ASAP7_75t_L g535 ( .A(n_444), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_478), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_448), .A2(n_630), .B(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_448), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_699) );
BUFx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_449), .A2(n_533), .B(n_534), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_449), .A2(n_689), .B1(n_931), .B2(n_932), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_449), .A2(n_529), .B1(n_966), .B2(n_967), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_449), .A2(n_458), .B1(n_1028), .B2(n_1029), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_449), .B(n_1137), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1250 ( .A1(n_449), .A2(n_458), .B1(n_1251), .B2(n_1252), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_449), .A2(n_1342), .B1(n_1343), .B2(n_1344), .Y(n_1341) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_449), .A2(n_1344), .B1(n_1355), .B2(n_1356), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g1420 ( .A1(n_449), .A2(n_689), .B1(n_1421), .B2(n_1422), .Y(n_1420) );
AND2x4_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g487 ( .A(n_451), .Y(n_487) );
INVx2_ASAP7_75t_SL g847 ( .A(n_451), .Y(n_847) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_452), .Y(n_551) );
AND2x2_ASAP7_75t_L g458 ( .A(n_453), .B(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g467 ( .A(n_453), .B(n_468), .Y(n_467) );
AND2x6_ASAP7_75t_L g474 ( .A(n_453), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g529 ( .A(n_453), .B(n_459), .Y(n_529) );
AND2x2_ASAP7_75t_L g689 ( .A(n_453), .B(n_459), .Y(n_689) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_453), .B(n_459), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_453), .B(n_847), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_453), .B(n_1044), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_453), .B(n_859), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_453), .B(n_459), .Y(n_1344) );
AND2x4_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g502 ( .A(n_454), .Y(n_502) );
INVx2_ASAP7_75t_L g853 ( .A(n_455), .Y(n_853) );
AND2x4_ASAP7_75t_L g870 ( .A(n_455), .B(n_551), .Y(n_870) );
AND2x2_ASAP7_75t_L g891 ( .A(n_455), .B(n_460), .Y(n_891) );
INVx1_ASAP7_75t_L g504 ( .A(n_456), .Y(n_504) );
INVx1_ASAP7_75t_L g537 ( .A(n_456), .Y(n_537) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g493 ( .A(n_460), .Y(n_493) );
BUFx6f_ASAP7_75t_L g1108 ( .A(n_460), .Y(n_1108) );
BUFx6f_ASAP7_75t_L g1133 ( .A(n_460), .Y(n_1133) );
AND2x4_ASAP7_75t_L g1719 ( .A(n_460), .B(n_1713), .Y(n_1719) );
BUFx2_ASAP7_75t_L g1730 ( .A(n_460), .Y(n_1730) );
INVx1_ASAP7_75t_L g1788 ( .A(n_460), .Y(n_1788) );
INVx1_ASAP7_75t_L g1795 ( .A(n_460), .Y(n_1795) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g714 ( .A(n_461), .Y(n_714) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_472), .B2(n_473), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g1781 ( .A1(n_466), .A2(n_531), .B1(n_1782), .B2(n_1783), .Y(n_1781) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g525 ( .A(n_467), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_467), .A2(n_474), .B1(n_629), .B2(n_686), .Y(n_685) );
BUFx2_ASAP7_75t_L g703 ( .A(n_467), .Y(n_703) );
BUFx2_ASAP7_75t_L g928 ( .A(n_467), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_467), .A2(n_474), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
BUFx2_ASAP7_75t_L g1248 ( .A(n_467), .Y(n_1248) );
BUFx3_ASAP7_75t_L g952 ( .A(n_468), .Y(n_952) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
INVx3_ASAP7_75t_L g1044 ( .A(n_469), .Y(n_1044) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_470), .Y(n_490) );
INVx1_ASAP7_75t_L g886 ( .A(n_470), .Y(n_886) );
INVx1_ASAP7_75t_L g1723 ( .A(n_470), .Y(n_1723) );
AND2x4_ASAP7_75t_L g476 ( .A(n_471), .B(n_477), .Y(n_476) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_473), .Y(n_698) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_474), .A2(n_524), .B1(n_525), .B2(n_526), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_474), .A2(n_927), .B1(n_928), .B2(n_929), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_474), .A2(n_703), .B1(n_963), .B2(n_964), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_474), .A2(n_1097), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_474), .A2(n_1247), .B1(n_1248), .B2(n_1249), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_474), .A2(n_928), .B1(n_1313), .B2(n_1340), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_474), .A2(n_928), .B1(n_1352), .B2(n_1353), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_474), .A2(n_1248), .B1(n_1398), .B2(n_1419), .Y(n_1418) );
AOI22xp5_ASAP7_75t_L g1778 ( .A1(n_474), .A2(n_1344), .B1(n_1779), .B2(n_1780), .Y(n_1778) );
NAND2x1p5_ASAP7_75t_L g715 ( .A(n_475), .B(n_510), .Y(n_715) );
BUFx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g495 ( .A(n_476), .Y(n_495) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_476), .Y(n_554) );
BUFx3_ASAP7_75t_L g564 ( .A(n_476), .Y(n_564) );
BUFx6f_ASAP7_75t_L g859 ( .A(n_476), .Y(n_859) );
INVx1_ASAP7_75t_L g1129 ( .A(n_476), .Y(n_1129) );
AND2x4_ASAP7_75t_L g1714 ( .A(n_476), .B(n_1715), .Y(n_1714) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_479), .B(n_506), .Y(n_478) );
AOI33xp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_485), .A3(n_491), .B1(n_496), .B2(n_497), .B3(n_498), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
BUFx2_ASAP7_75t_L g606 ( .A(n_483), .Y(n_606) );
OR2x6_ASAP7_75t_L g816 ( .A(n_483), .B(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g842 ( .A(n_483), .Y(n_842) );
AOI31xp33_ASAP7_75t_L g990 ( .A1(n_483), .A2(n_991), .A3(n_1003), .B(n_1015), .Y(n_990) );
AND2x4_ASAP7_75t_L g1111 ( .A(n_483), .B(n_484), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_483), .B(n_862), .Y(n_1135) );
INVx1_ASAP7_75t_L g877 ( .A(n_484), .Y(n_877) );
BUFx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_489), .A2(n_1034), .B1(n_1035), .B2(n_1036), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_489), .A2(n_1263), .B1(n_1363), .B2(n_1364), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_489), .A2(n_1366), .B1(n_1367), .B2(n_1368), .Y(n_1365) );
INVx4_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g560 ( .A(n_490), .Y(n_560) );
INVx2_ASAP7_75t_SL g722 ( .A(n_490), .Y(n_722) );
INVx2_ASAP7_75t_SL g856 ( .A(n_490), .Y(n_856) );
BUFx3_ASAP7_75t_L g1433 ( .A(n_490), .Y(n_1433) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_L g517 ( .A(n_495), .B(n_510), .Y(n_517) );
INVx1_ASAP7_75t_L g738 ( .A(n_498), .Y(n_738) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_499), .A2(n_535), .B1(n_538), .B2(n_555), .Y(n_534) );
OAI33xp33_ASAP7_75t_L g937 ( .A1(n_499), .A2(n_535), .A3(n_938), .B1(n_944), .B2(n_950), .B3(n_953), .Y(n_937) );
OAI33xp33_ASAP7_75t_L g1032 ( .A1(n_499), .A2(n_535), .A3(n_1033), .B1(n_1037), .B2(n_1041), .B3(n_1046), .Y(n_1032) );
OAI33xp33_ASAP7_75t_L g1254 ( .A1(n_499), .A2(n_1255), .A3(n_1256), .B1(n_1261), .B2(n_1266), .B3(n_1271), .Y(n_1254) );
OAI33xp33_ASAP7_75t_L g1358 ( .A1(n_499), .A2(n_1255), .A3(n_1359), .B1(n_1362), .B2(n_1365), .B3(n_1369), .Y(n_1358) );
OAI33xp33_ASAP7_75t_L g1425 ( .A1(n_499), .A2(n_535), .A3(n_1426), .B1(n_1430), .B2(n_1435), .B3(n_1436), .Y(n_1425) );
CKINVDCx8_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
INVx5_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx6_ASAP7_75t_L g683 ( .A(n_501), .Y(n_683) );
OR2x6_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g862 ( .A(n_503), .Y(n_862) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g1716 ( .A(n_504), .Y(n_1716) );
AOI221xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_511), .B1(n_512), .B2(n_516), .C(n_517), .Y(n_506) );
INVx1_ASAP7_75t_L g611 ( .A(n_507), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g1116 ( .A1(n_507), .A2(n_517), .B(n_1117), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_507), .A2(n_512), .B1(n_517), .B2(n_1123), .C(n_1124), .Y(n_1122) );
AOI221xp5_ASAP7_75t_L g1328 ( .A1(n_507), .A2(n_512), .B1(n_517), .B2(n_1329), .C(n_1330), .Y(n_1328) );
AOI221xp5_ASAP7_75t_L g1775 ( .A1(n_507), .A2(n_512), .B1(n_517), .B2(n_1776), .C(n_1777), .Y(n_1775) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
AND2x2_ASAP7_75t_L g865 ( .A(n_508), .B(n_844), .Y(n_865) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g709 ( .A(n_509), .Y(n_709) );
AND2x4_ASAP7_75t_L g512 ( .A(n_510), .B(n_513), .Y(n_512) );
NAND2x1_ASAP7_75t_SL g707 ( .A(n_510), .B(n_708), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g712 ( .A(n_510), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g609 ( .A(n_512), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_512), .A2(n_531), .B1(n_1081), .B2(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g663 ( .A(n_515), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_515), .B(n_664), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_517), .A2(n_595), .B1(n_596), .B2(n_608), .C(n_610), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_517), .A2(n_608), .B1(n_610), .B2(n_650), .C(n_652), .Y(n_690) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
XOR2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_612), .Y(n_519) );
NAND4xp25_ASAP7_75t_L g521 ( .A(n_522), .B(n_532), .C(n_565), .D(n_607), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .Y(n_522) );
OAI221xp5_ASAP7_75t_L g583 ( .A1(n_526), .A2(n_533), .B1(n_584), .B2(n_586), .C(n_588), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_528), .A2(n_529), .B1(n_530), .B2(n_531), .Y(n_527) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_531), .A2(n_637), .B1(n_688), .B2(n_689), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_531), .A2(n_1104), .B1(n_1143), .B2(n_1144), .Y(n_1142) );
OAI33xp33_ASAP7_75t_L g655 ( .A1(n_535), .A2(n_656), .A3(n_665), .B1(n_670), .B2(n_675), .B3(n_682), .Y(n_655) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_535), .Y(n_717) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_535), .Y(n_1255) );
INVx1_ASAP7_75t_L g1713 ( .A(n_537), .Y(n_1713) );
OAI221xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_543), .B1(n_544), .B2(n_547), .C(n_548), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g558 ( .A(n_542), .Y(n_558) );
INVx1_ASAP7_75t_L g668 ( .A(n_542), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g571 ( .A1(n_543), .A2(n_572), .B1(n_574), .B2(n_575), .C(n_577), .Y(n_571) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_546), .A2(n_620), .B1(n_666), .B2(n_669), .Y(n_665) );
INVx3_ASAP7_75t_L g673 ( .A(n_546), .Y(n_673) );
INVx2_ASAP7_75t_L g1131 ( .A(n_546), .Y(n_1131) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_SL g860 ( .A(n_550), .Y(n_860) );
INVx2_ASAP7_75t_L g1127 ( .A(n_550), .Y(n_1127) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx6f_ASAP7_75t_L g1110 ( .A(n_551), .Y(n_1110) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g1333 ( .A(n_553), .Y(n_1333) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
OAI221xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .B1(n_560), .B2(n_561), .C(n_562), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_556), .A2(n_671), .B1(n_672), .B2(n_674), .Y(n_670) );
BUFx2_ASAP7_75t_L g979 ( .A(n_556), .Y(n_979) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g727 ( .A(n_557), .Y(n_727) );
INVx2_ASAP7_75t_L g855 ( .A(n_557), .Y(n_855) );
BUFx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g948 ( .A(n_558), .Y(n_948) );
OAI22xp5_ASAP7_75t_SL g944 ( .A1(n_560), .A2(n_945), .B1(n_946), .B2(n_949), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_560), .A2(n_979), .B1(n_980), .B2(n_981), .Y(n_978) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x4_ASAP7_75t_L g851 ( .A(n_564), .B(n_852), .Y(n_851) );
OAI31xp33_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_579), .A3(n_589), .B(n_605), .Y(n_565) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g1012 ( .A(n_570), .Y(n_1012) );
OAI21xp5_ASAP7_75t_SL g1312 ( .A1(n_572), .A2(n_1313), .B(n_1314), .Y(n_1312) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g618 ( .A(n_573), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_575), .A2(n_618), .B1(n_619), .B2(n_620), .C(n_621), .Y(n_617) );
INVx1_ASAP7_75t_L g1281 ( .A(n_575), .Y(n_1281) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g1409 ( .A(n_577), .Y(n_1409) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g769 ( .A(n_578), .Y(n_769) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g603 ( .A(n_582), .Y(n_603) );
BUFx2_ASAP7_75t_L g764 ( .A(n_582), .Y(n_764) );
BUFx3_ASAP7_75t_L g830 ( .A(n_582), .Y(n_830) );
OAI211xp5_ASAP7_75t_L g1397 ( .A1(n_584), .A2(n_1398), .B(n_1399), .C(n_1400), .Y(n_1397) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_SL g604 ( .A(n_585), .Y(n_604) );
INVx1_ASAP7_75t_L g1150 ( .A(n_585), .Y(n_1150) );
OAI221xp5_ASAP7_75t_L g628 ( .A1(n_586), .A2(n_604), .B1(n_629), .B2(n_630), .C(n_631), .Y(n_628) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_594), .C(n_597), .Y(n_589) );
A2O1A1Ixp33_ASAP7_75t_SL g634 ( .A1(n_592), .A2(n_635), .B(n_637), .C(n_638), .Y(n_634) );
A2O1A1Ixp33_ASAP7_75t_L g1080 ( .A1(n_592), .A2(n_635), .B(n_1081), .C(n_1082), .Y(n_1080) );
BUFx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g1310 ( .A(n_603), .Y(n_1310) );
CKINVDCx8_ASAP7_75t_R g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND4xp25_ASAP7_75t_L g613 ( .A(n_614), .B(n_654), .C(n_684), .D(n_690), .Y(n_613) );
OAI31xp33_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_623), .A3(n_633), .B(n_653), .Y(n_614) );
INVx2_ASAP7_75t_SL g1771 ( .A(n_616), .Y(n_1771) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_619), .A2(n_657), .B1(n_658), .B2(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g787 ( .A(n_625), .Y(n_787) );
BUFx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g642 ( .A(n_627), .Y(n_642) );
INVx1_ASAP7_75t_L g832 ( .A(n_627), .Y(n_832) );
BUFx6f_ASAP7_75t_L g907 ( .A(n_627), .Y(n_907) );
INVx1_ASAP7_75t_L g758 ( .A(n_631), .Y(n_758) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND3xp33_ASAP7_75t_SL g633 ( .A(n_634), .B(n_640), .C(n_646), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g828 ( .A(n_636), .Y(n_828) );
INVx4_ASAP7_75t_L g903 ( .A(n_636), .Y(n_903) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g913 ( .A(n_639), .Y(n_913) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g1405 ( .A(n_645), .Y(n_1405) );
BUFx2_ASAP7_75t_L g1739 ( .A(n_645), .Y(n_1739) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx4_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_649), .A2(n_651), .B1(n_1123), .B2(n_1124), .Y(n_1165) );
INVx2_ASAP7_75t_L g1284 ( .A(n_649), .Y(n_1284) );
INVx1_ASAP7_75t_SL g1773 ( .A(n_649), .Y(n_1773) );
INVx2_ASAP7_75t_SL g1059 ( .A(n_651), .Y(n_1059) );
INVx2_ASAP7_75t_L g1285 ( .A(n_651), .Y(n_1285) );
OAI31xp33_ASAP7_75t_L g1145 ( .A1(n_653), .A2(n_1146), .A3(n_1147), .B(n_1159), .Y(n_1145) );
AOI22xp5_ASAP7_75t_L g1302 ( .A1(n_653), .A2(n_742), .B1(n_1303), .B2(n_1326), .Y(n_1302) );
INVx2_ASAP7_75t_L g1415 ( .A(n_653), .Y(n_1415) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_658), .A2(n_676), .B1(n_677), .B2(n_681), .Y(n_675) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g720 ( .A(n_659), .Y(n_720) );
INVx1_ASAP7_75t_L g1427 ( .A(n_659), .Y(n_1427) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g1215 ( .A(n_661), .Y(n_1215) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g888 ( .A(n_662), .B(n_845), .Y(n_888) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_662), .Y(n_984) );
OR2x6_ASAP7_75t_L g1212 ( .A(n_662), .B(n_845), .Y(n_1212) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g943 ( .A(n_663), .Y(n_943) );
BUFx2_ASAP7_75t_L g955 ( .A(n_663), .Y(n_955) );
INVx3_ASAP7_75t_L g1049 ( .A(n_663), .Y(n_1049) );
BUFx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_668), .Y(n_880) );
INVx2_ASAP7_75t_L g1264 ( .A(n_668), .Y(n_1264) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g729 ( .A(n_678), .Y(n_729) );
INVx1_ASAP7_75t_L g1039 ( .A(n_678), .Y(n_1039) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx3_ASAP7_75t_L g736 ( .A(n_679), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g1789 ( .A1(n_679), .A2(n_1790), .B1(n_1791), .B2(n_1792), .Y(n_1789) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g986 ( .A(n_683), .Y(n_986) );
AOI322xp5_ASAP7_75t_L g1106 ( .A1(n_683), .A2(n_1090), .A3(n_1107), .B1(n_1109), .B2(n_1111), .C1(n_1112), .C2(n_1115), .Y(n_1106) );
AOI33xp33_ASAP7_75t_L g1331 ( .A1(n_683), .A2(n_1111), .A3(n_1332), .B1(n_1334), .B2(n_1335), .B3(n_1338), .Y(n_1331) );
AOI33xp33_ASAP7_75t_L g1725 ( .A1(n_683), .A2(n_1111), .A3(n_1726), .B1(n_1727), .B2(n_1729), .B3(n_1731), .Y(n_1725) );
AOI222xp33_ASAP7_75t_L g1784 ( .A1(n_683), .A2(n_1102), .B1(n_1111), .B2(n_1785), .C1(n_1786), .C2(n_1793), .Y(n_1784) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
XNOR2x1_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_739), .Y(n_695) );
NOR3xp33_ASAP7_75t_SL g696 ( .A(n_697), .B(n_704), .C(n_716), .Y(n_696) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_SL g934 ( .A(n_706), .Y(n_934) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2x1p5_ASAP7_75t_L g1218 ( .A(n_708), .B(n_1219), .Y(n_1218) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx4f_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
BUFx4f_ASAP7_75t_L g935 ( .A(n_712), .Y(n_935) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OR2x6_ASAP7_75t_L g867 ( .A(n_714), .B(n_845), .Y(n_867) );
BUFx3_ASAP7_75t_L g936 ( .A(n_715), .Y(n_936) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_715), .Y(n_1031) );
BUFx2_ASAP7_75t_L g1424 ( .A(n_715), .Y(n_1424) );
OAI33xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .A3(n_723), .B1(n_730), .B2(n_733), .B3(n_738), .Y(n_716) );
OAI33xp33_ASAP7_75t_L g969 ( .A1(n_717), .A2(n_970), .A3(n_973), .B1(n_978), .B2(n_982), .B3(n_986), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g733 ( .A1(n_720), .A2(n_734), .B1(n_735), .B2(n_737), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_722), .A2(n_725), .B1(n_731), .B2(n_732), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g1261 ( .A1(n_722), .A2(n_1262), .B1(n_1263), .B2(n_1265), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_728), .B2(n_729), .Y(n_723) );
OAI22xp33_ASAP7_75t_SL g973 ( .A1(n_725), .A2(n_974), .B1(n_976), .B2(n_977), .Y(n_973) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_727), .A2(n_1267), .B1(n_1268), .B2(n_1270), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g1435 ( .A1(n_727), .A2(n_1268), .B1(n_1395), .B2(n_1414), .Y(n_1435) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_729), .A2(n_856), .B1(n_971), .B2(n_972), .Y(n_970) );
OAI22xp33_ASAP7_75t_L g1369 ( .A1(n_729), .A2(n_1257), .B1(n_1370), .B2(n_1371), .Y(n_1369) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_731), .A2(n_746), .B(n_747), .Y(n_745) );
OAI221xp5_ASAP7_75t_L g871 ( .A1(n_735), .A2(n_872), .B1(n_873), .B2(n_875), .C(n_876), .Y(n_871) );
BUFx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_737), .A2(n_760), .B1(n_763), .B2(n_770), .C(n_773), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_743), .B(n_744), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_742), .A2(n_898), .B1(n_899), .B2(n_923), .Y(n_897) );
AOI21xp33_ASAP7_75t_SL g1051 ( .A1(n_742), .A2(n_1052), .B(n_1053), .Y(n_1051) );
AOI21xp33_ASAP7_75t_SL g1391 ( .A1(n_742), .A2(n_1392), .B(n_1393), .Y(n_1391) );
OR2x6_ASAP7_75t_L g813 ( .A(n_750), .B(n_810), .Y(n_813) );
INVx1_ASAP7_75t_L g1007 ( .A(n_752), .Y(n_1007) );
INVx1_ASAP7_75t_L g1057 ( .A(n_752), .Y(n_1057) );
INVx1_ASAP7_75t_L g1734 ( .A(n_752), .Y(n_1734) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx3_ASAP7_75t_L g1193 ( .A(n_768), .Y(n_1193) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g1066 ( .A(n_777), .Y(n_1066) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_1018), .B2(n_1064), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
XNOR2x1_ASAP7_75t_L g779 ( .A(n_780), .B(n_894), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_838), .C(n_848), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_803), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_794), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_786), .B1(n_790), .B2(n_791), .Y(n_784) );
OAI221xp5_ASAP7_75t_L g854 ( .A1(n_785), .A2(n_790), .B1(n_855), .B2(n_856), .C(n_857), .Y(n_854) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
AND2x2_ASAP7_75t_L g796 ( .A(n_788), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OR2x6_ASAP7_75t_L g792 ( .A(n_789), .B(n_793), .Y(n_792) );
OR2x6_ASAP7_75t_L g801 ( .A(n_789), .B(n_802), .Y(n_801) );
CKINVDCx6p67_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_796), .B1(n_799), .B2(n_800), .Y(n_794) );
INVx2_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g916 ( .A(n_798), .Y(n_916) );
CKINVDCx6p67_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
BUFx3_ASAP7_75t_L g1086 ( .A(n_802), .Y(n_1086) );
INVx1_ASAP7_75t_L g1092 ( .A(n_802), .Y(n_1092) );
NAND3xp33_ASAP7_75t_SL g803 ( .A(n_804), .B(n_814), .C(n_834), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_811), .B2(n_812), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_805), .A2(n_811), .B1(n_864), .B2(n_866), .Y(n_863) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NAND2x1p5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
INVx2_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g837 ( .A(n_810), .Y(n_837) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
AOI33xp33_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_818), .A3(n_823), .B1(n_826), .B2(n_829), .B3(n_833), .Y(n_814) );
AOI33xp33_ASAP7_75t_L g1732 ( .A1(n_815), .A2(n_833), .A3(n_1733), .B1(n_1735), .B2(n_1736), .B3(n_1738), .Y(n_1732) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g1232 ( .A(n_816), .Y(n_1232) );
INVx1_ASAP7_75t_L g1010 ( .A(n_817), .Y(n_1010) );
BUFx3_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_822), .B(n_837), .Y(n_836) );
BUFx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx4_ASAP7_75t_L g1238 ( .A(n_833), .Y(n_1238) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
NOR2xp67_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
AOI211xp5_ASAP7_75t_L g1075 ( .A1(n_842), .A2(n_1076), .B(n_1095), .C(n_1105), .Y(n_1075) );
INVx1_ASAP7_75t_L g1224 ( .A(n_843), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_847), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g1219 ( .A(n_845), .Y(n_1219) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx8_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
AOI222xp33_ASAP7_75t_L g1223 ( .A1(n_851), .A2(n_870), .B1(n_1181), .B2(n_1224), .C1(n_1225), .C2(n_1226), .Y(n_1223) );
AND2x4_ASAP7_75t_L g893 ( .A(n_852), .B(n_885), .Y(n_893) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
BUFx6f_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_SL g861 ( .A(n_862), .Y(n_861) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
CKINVDCx11_ASAP7_75t_R g866 ( .A(n_867), .Y(n_866) );
CKINVDCx6p67_ASAP7_75t_R g869 ( .A(n_870), .Y(n_869) );
OAI22xp33_ASAP7_75t_L g1037 ( .A1(n_873), .A2(n_1038), .B1(n_1039), .B2(n_1040), .Y(n_1037) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_881), .B1(n_882), .B2(n_887), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx3_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_891), .A2(n_893), .B1(n_1228), .B2(n_1229), .Y(n_1227) );
INVx3_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
AO22x2_ASAP7_75t_L g894 ( .A1(n_895), .A2(n_957), .B1(n_1016), .B2(n_1017), .Y(n_894) );
INVx1_ASAP7_75t_L g1017 ( .A(n_895), .Y(n_1017) );
XOR2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_956), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_897), .B(n_924), .Y(n_896) );
NAND3xp33_ASAP7_75t_L g899 ( .A(n_900), .B(n_911), .C(n_920), .Y(n_899) );
BUFx2_ASAP7_75t_L g1008 ( .A(n_902), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g950 ( .A1(n_908), .A2(n_922), .B1(n_946), .B2(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g1282 ( .A(n_918), .Y(n_1282) );
INVx1_ASAP7_75t_L g1311 ( .A(n_918), .Y(n_1311) );
OAI22xp33_ASAP7_75t_L g953 ( .A1(n_919), .A2(n_921), .B1(n_940), .B2(n_954), .Y(n_953) );
NOR3xp33_ASAP7_75t_L g924 ( .A(n_925), .B(n_933), .C(n_937), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_930), .Y(n_925) );
OAI22xp33_ASAP7_75t_L g938 ( .A1(n_939), .A2(n_940), .B1(n_942), .B2(n_943), .Y(n_938) );
BUFx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
OAI22xp33_ASAP7_75t_L g982 ( .A1(n_941), .A2(n_983), .B1(n_984), .B2(n_985), .Y(n_982) );
INVx1_ASAP7_75t_L g1258 ( .A(n_941), .Y(n_1258) );
INVx1_ASAP7_75t_L g1438 ( .A(n_941), .Y(n_1438) );
INVx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx2_ASAP7_75t_L g1035 ( .A(n_947), .Y(n_1035) );
INVx2_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
BUFx2_ASAP7_75t_L g1366 ( .A(n_948), .Y(n_1366) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_952), .Y(n_951) );
OAI22xp33_ASAP7_75t_L g1426 ( .A1(n_954), .A2(n_1427), .B1(n_1428), .B2(n_1429), .Y(n_1426) );
INVx2_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g1016 ( .A(n_957), .Y(n_1016) );
XNOR2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_959), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_960), .B(n_987), .Y(n_959) );
NOR3xp33_ASAP7_75t_SL g960 ( .A(n_961), .B(n_968), .C(n_969), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_962), .B(n_965), .Y(n_961) );
OAI22xp33_ASAP7_75t_L g1046 ( .A1(n_974), .A2(n_1047), .B1(n_1048), .B2(n_1050), .Y(n_1046) );
INVx3_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
AOI21xp5_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_989), .B(n_990), .Y(n_987) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
AOI31xp33_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_998), .A3(n_1000), .B(n_1001), .Y(n_993) );
INVx1_ASAP7_75t_L g1770 ( .A(n_995), .Y(n_1770) );
BUFx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx2_ASAP7_75t_L g1164 ( .A(n_997), .Y(n_1164) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
BUFx2_ASAP7_75t_SL g1019 ( .A(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1020), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1051), .Y(n_1021) );
NOR3xp33_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1030), .C(n_1032), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1027), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_1035), .A2(n_1042), .B1(n_1043), .B2(n_1045), .Y(n_1041) );
INVx2_ASAP7_75t_L g1796 ( .A(n_1043), .Y(n_1796) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1044), .Y(n_1269) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1044), .Y(n_1337) );
OAI22xp33_ASAP7_75t_L g1256 ( .A1(n_1048), .A2(n_1257), .B1(n_1259), .B2(n_1260), .Y(n_1256) );
OAI22xp33_ASAP7_75t_L g1271 ( .A1(n_1048), .A2(n_1257), .B1(n_1272), .B2(n_1273), .Y(n_1271) );
OAI22xp33_ASAP7_75t_L g1359 ( .A1(n_1048), .A2(n_1257), .B1(n_1360), .B2(n_1361), .Y(n_1359) );
OAI22xp33_ASAP7_75t_L g1436 ( .A1(n_1048), .A2(n_1402), .B1(n_1413), .B2(n_1437), .Y(n_1436) );
BUFx2_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1071), .B1(n_1386), .B2(n_1387), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
AOI22xp5_ASAP7_75t_L g1071 ( .A1(n_1072), .A2(n_1073), .B1(n_1167), .B2(n_1168), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
AOI22xp5_ASAP7_75t_L g1073 ( .A1(n_1074), .A2(n_1118), .B1(n_1119), .B2(n_1166), .Y(n_1073) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1074), .Y(n_1166) );
NAND4xp25_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1080), .C(n_1084), .D(n_1089), .Y(n_1076) );
OAI211xp5_ASAP7_75t_L g1084 ( .A1(n_1085), .A2(n_1086), .B(n_1087), .C(n_1088), .Y(n_1084) );
OAI211xp5_ASAP7_75t_L g1154 ( .A1(n_1086), .A2(n_1141), .B(n_1155), .C(n_1156), .Y(n_1154) );
OAI211xp5_ASAP7_75t_L g1089 ( .A1(n_1090), .A2(n_1091), .B(n_1093), .C(n_1094), .Y(n_1089) );
OAI221xp5_ASAP7_75t_L g1233 ( .A1(n_1091), .A2(n_1234), .B1(n_1235), .B2(n_1236), .C(n_1237), .Y(n_1233) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1102), .B1(n_1103), .B2(n_1104), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1116), .Y(n_1105) );
AOI33xp33_ASAP7_75t_L g1125 ( .A1(n_1111), .A2(n_1126), .A3(n_1130), .B1(n_1132), .B2(n_1134), .B3(n_1135), .Y(n_1125) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
NAND3xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1138), .C(n_1145), .Y(n_1120) );
AND3x1_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1125), .C(n_1136), .Y(n_1121) );
INVx2_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1142), .Y(n_1138) );
NAND3xp33_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1154), .C(n_1157), .Y(n_1147) );
OAI211xp5_ASAP7_75t_L g1148 ( .A1(n_1149), .A2(n_1150), .B(n_1151), .C(n_1153), .Y(n_1148) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1152), .Y(n_1293) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1757 ( .A1(n_1158), .A2(n_1758), .B1(n_1759), .B2(n_1760), .C(n_1762), .Y(n_1757) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1164), .Y(n_1241) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
XNOR2xp5_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1298), .Y(n_1168) );
AO22x2_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1171), .B1(n_1242), .B2(n_1297), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
NAND4xp25_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1180), .C(n_1189), .D(n_1201), .Y(n_1173) );
BUFx2_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx5_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
CKINVDCx8_ASAP7_75t_R g1696 ( .A(n_1176), .Y(n_1696) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1178), .Y(n_1702) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_1181), .A2(n_1182), .B1(n_1185), .B2(n_1186), .Y(n_1180) );
INVx4_ASAP7_75t_L g1703 ( .A(n_1182), .Y(n_1703) );
AND2x4_ASAP7_75t_L g1196 ( .A(n_1183), .B(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
INVx4_ASAP7_75t_L g1699 ( .A(n_1186), .Y(n_1699) );
AND2x4_ASAP7_75t_L g1203 ( .A(n_1187), .B(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_SL g1187 ( .A(n_1188), .Y(n_1187) );
AOI222xp33_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1191), .B1(n_1194), .B2(n_1195), .C1(n_1199), .C2(n_1200), .Y(n_1189) );
OAI21xp5_ASAP7_75t_SL g1214 ( .A1(n_1190), .A2(n_1215), .B(n_1216), .Y(n_1214) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
BUFx4f_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1693 ( .A1(n_1196), .A2(n_1200), .B1(n_1694), .B2(n_1695), .Y(n_1693) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_1202), .A2(n_1203), .B1(n_1205), .B2(n_1206), .Y(n_1201) );
CKINVDCx6p67_ASAP7_75t_R g1698 ( .A(n_1206), .Y(n_1698) );
NAND3xp33_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1223), .C(n_1227), .Y(n_1209) );
NOR3xp33_ASAP7_75t_SL g1210 ( .A(n_1211), .B(n_1213), .C(n_1217), .Y(n_1210) );
INVx2_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1222), .Y(n_1220) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_1231), .A2(n_1233), .B1(n_1238), .B2(n_1239), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1242), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1274), .Y(n_1243) );
NOR3xp33_ASAP7_75t_SL g1244 ( .A(n_1245), .B(n_1253), .C(n_1254), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1250), .Y(n_1245) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
BUFx2_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1430 ( .A1(n_1264), .A2(n_1431), .B1(n_1432), .B2(n_1434), .Y(n_1430) );
HB1xp67_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx2_ASAP7_75t_L g1728 ( .A(n_1269), .Y(n_1728) );
NAND3xp33_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1286), .C(n_1294), .Y(n_1275) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
XOR2x2_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1346), .Y(n_1299) );
XNOR2xp5_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1345), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1327), .Y(n_1301) );
NAND3xp33_ASAP7_75t_SL g1303 ( .A(n_1304), .B(n_1316), .C(n_1323), .Y(n_1303) );
INVx2_ASAP7_75t_SL g1307 ( .A(n_1308), .Y(n_1307) );
BUFx3_ASAP7_75t_L g1411 ( .A(n_1315), .Y(n_1411) );
HB1xp67_ASAP7_75t_L g1737 ( .A(n_1315), .Y(n_1737) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
AND4x1_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1331), .C(n_1339), .D(n_1341), .Y(n_1327) );
INVx2_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
XNOR2x1_ASAP7_75t_L g1346 ( .A(n_1347), .B(n_1348), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1349), .B(n_1372), .Y(n_1348) );
NOR3xp33_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1357), .C(n_1358), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1351), .B(n_1354), .Y(n_1350) );
NAND3xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1378), .C(n_1381), .Y(n_1373) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
XNOR2x1_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1439), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1391), .B(n_1416), .Y(n_1390) );
AOI31xp33_ASAP7_75t_L g1393 ( .A1(n_1394), .A2(n_1401), .A3(n_1412), .B(n_1415), .Y(n_1393) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
HB1xp67_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
AOI21xp5_ASAP7_75t_L g1756 ( .A1(n_1415), .A2(n_1757), .B(n_1765), .Y(n_1756) );
NOR3xp33_ASAP7_75t_SL g1416 ( .A(n_1417), .B(n_1423), .C(n_1425), .Y(n_1416) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1420), .Y(n_1417) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
OAI221xp5_ASAP7_75t_L g1441 ( .A1(n_1442), .A2(n_1682), .B1(n_1683), .B2(n_1742), .C(n_1748), .Y(n_1441) );
AOI21xp5_ASAP7_75t_L g1442 ( .A1(n_1443), .A2(n_1587), .B(n_1631), .Y(n_1442) );
NAND5xp2_ASAP7_75t_SL g1443 ( .A(n_1444), .B(n_1526), .C(n_1555), .D(n_1578), .E(n_1582), .Y(n_1443) );
AOI21xp5_ASAP7_75t_L g1444 ( .A1(n_1445), .A2(n_1483), .B(n_1504), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1466), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1446), .B(n_1493), .Y(n_1543) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1446), .B(n_1581), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1605 ( .A(n_1446), .B(n_1515), .Y(n_1605) );
NOR2xp33_ASAP7_75t_L g1616 ( .A(n_1446), .B(n_1493), .Y(n_1616) );
INVx2_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1447), .B(n_1513), .Y(n_1512) );
NAND2xp5_ASAP7_75t_L g1525 ( .A(n_1447), .B(n_1493), .Y(n_1525) );
BUFx2_ASAP7_75t_L g1532 ( .A(n_1447), .Y(n_1532) );
INVx2_ASAP7_75t_L g1539 ( .A(n_1447), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_1447), .B(n_1466), .Y(n_1590) );
OR2x2_ASAP7_75t_L g1614 ( .A(n_1447), .B(n_1523), .Y(n_1614) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1447), .B(n_1515), .Y(n_1647) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1448), .B(n_1460), .Y(n_1447) );
AND2x4_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1455), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
OR2x2_ASAP7_75t_L g1480 ( .A(n_1451), .B(n_1456), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1454), .Y(n_1451) );
HB1xp67_ASAP7_75t_L g1802 ( .A(n_1452), .Y(n_1802) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1454), .Y(n_1463) );
AND2x4_ASAP7_75t_L g1457 ( .A(n_1455), .B(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
OR2x2_ASAP7_75t_L g1482 ( .A(n_1456), .B(n_1459), .Y(n_1482) );
BUFx2_ASAP7_75t_L g1488 ( .A(n_1457), .Y(n_1488) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1461), .Y(n_1502) );
BUFx3_ASAP7_75t_L g1547 ( .A(n_1461), .Y(n_1547) );
AND2x4_ASAP7_75t_L g1461 ( .A(n_1462), .B(n_1464), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1471 ( .A(n_1462), .B(n_1464), .Y(n_1471) );
HB1xp67_ASAP7_75t_L g1803 ( .A(n_1462), .Y(n_1803) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
AND2x4_ASAP7_75t_L g1465 ( .A(n_1463), .B(n_1464), .Y(n_1465) );
INVx2_ASAP7_75t_L g1491 ( .A(n_1465), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1467), .B(n_1472), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1518 ( .A(n_1467), .B(n_1519), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_1467), .B(n_1510), .Y(n_1575) );
A2O1A1Ixp33_ASAP7_75t_L g1648 ( .A1(n_1467), .A2(n_1649), .B(n_1652), .C(n_1653), .Y(n_1648) );
INVxp67_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
BUFx2_ASAP7_75t_L g1513 ( .A(n_1468), .Y(n_1513) );
BUFx3_ASAP7_75t_L g1523 ( .A(n_1468), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1468), .B(n_1510), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1470), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1544 ( .A(n_1472), .B(n_1513), .Y(n_1544) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1472), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1477), .Y(n_1472) );
NAND2xp5_ASAP7_75t_L g1528 ( .A(n_1473), .B(n_1523), .Y(n_1528) );
NOR2xp33_ASAP7_75t_L g1594 ( .A(n_1473), .B(n_1513), .Y(n_1594) );
INVx2_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
OR2x2_ASAP7_75t_L g1511 ( .A(n_1474), .B(n_1477), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_1474), .B(n_1520), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1522 ( .A(n_1474), .B(n_1523), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1474), .B(n_1477), .Y(n_1559) );
NOR2xp33_ASAP7_75t_L g1566 ( .A(n_1474), .B(n_1523), .Y(n_1566) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1475), .B(n_1476), .Y(n_1474) );
INVx2_ASAP7_75t_SL g1520 ( .A(n_1477), .Y(n_1520) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_1477), .B(n_1523), .Y(n_1540) );
OAI22xp5_ASAP7_75t_L g1478 ( .A1(n_1479), .A2(n_1480), .B1(n_1481), .B2(n_1482), .Y(n_1478) );
BUFx6f_ASAP7_75t_L g1496 ( .A(n_1480), .Y(n_1496) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1482), .Y(n_1499) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1483), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1484), .B(n_1492), .Y(n_1483) );
NAND2xp5_ASAP7_75t_L g1553 ( .A(n_1484), .B(n_1554), .Y(n_1553) );
INVx2_ASAP7_75t_L g1570 ( .A(n_1484), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1484), .B(n_1585), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1620 ( .A(n_1484), .B(n_1493), .Y(n_1620) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1485), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1668 ( .A(n_1485), .B(n_1505), .Y(n_1668) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
OR2x2_ASAP7_75t_L g1561 ( .A(n_1486), .B(n_1505), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1486), .B(n_1516), .Y(n_1563) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1486), .Y(n_1643) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1487), .B(n_1489), .Y(n_1486) );
INVx2_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
NAND2xp5_ASAP7_75t_L g1562 ( .A(n_1492), .B(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1492), .Y(n_1630) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1493), .B(n_1505), .Y(n_1533) );
INVx2_ASAP7_75t_SL g1569 ( .A(n_1493), .Y(n_1569) );
AND2x4_ASAP7_75t_L g1585 ( .A(n_1493), .B(n_1516), .Y(n_1585) );
HB1xp67_ASAP7_75t_L g1622 ( .A(n_1493), .Y(n_1622) );
CKINVDCx5p33_ASAP7_75t_R g1493 ( .A(n_1494), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1494), .B(n_1516), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1494), .B(n_1505), .Y(n_1577) );
OR2x2_ASAP7_75t_L g1494 ( .A(n_1495), .B(n_1501), .Y(n_1494) );
OAI22xp5_ASAP7_75t_L g1495 ( .A1(n_1496), .A2(n_1497), .B1(n_1498), .B2(n_1500), .Y(n_1495) );
BUFx3_ASAP7_75t_L g1550 ( .A(n_1496), .Y(n_1550) );
HB1xp67_ASAP7_75t_L g1552 ( .A(n_1498), .Y(n_1552) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
OAI211xp5_ASAP7_75t_SL g1504 ( .A1(n_1505), .A2(n_1508), .B(n_1514), .C(n_1521), .Y(n_1504) );
INVx3_ASAP7_75t_L g1516 ( .A(n_1505), .Y(n_1516) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1505), .Y(n_1607) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1506), .B(n_1507), .Y(n_1505) );
OAI321xp33_ASAP7_75t_L g1613 ( .A1(n_1508), .A2(n_1528), .A3(n_1559), .B1(n_1607), .B2(n_1614), .C(n_1615), .Y(n_1613) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1509), .B(n_1569), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1659 ( .A(n_1509), .B(n_1660), .Y(n_1659) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1512), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1510), .B(n_1539), .Y(n_1624) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
OR2x2_ASAP7_75t_L g1637 ( .A(n_1511), .B(n_1614), .Y(n_1637) );
NAND2xp5_ASAP7_75t_L g1645 ( .A(n_1512), .B(n_1559), .Y(n_1645) );
NOR2x1_ASAP7_75t_L g1612 ( .A(n_1513), .B(n_1520), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1513), .B(n_1559), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g1514 ( .A(n_1515), .B(n_1517), .Y(n_1514) );
AOI221xp5_ASAP7_75t_L g1588 ( .A1(n_1515), .A2(n_1589), .B1(n_1591), .B2(n_1597), .C(n_1598), .Y(n_1588) );
NOR2xp33_ASAP7_75t_L g1524 ( .A(n_1516), .B(n_1525), .Y(n_1524) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1516), .Y(n_1536) );
OR2x2_ASAP7_75t_L g1642 ( .A(n_1516), .B(n_1643), .Y(n_1642) );
AOI221xp5_ASAP7_75t_L g1657 ( .A1(n_1516), .A2(n_1560), .B1(n_1658), .B2(n_1661), .C(n_1664), .Y(n_1657) );
O2A1O1Ixp33_ASAP7_75t_L g1601 ( .A1(n_1517), .A2(n_1584), .B(n_1602), .C(n_1604), .Y(n_1601) );
AOI222xp33_ASAP7_75t_L g1638 ( .A1(n_1517), .A2(n_1563), .B1(n_1639), .B2(n_1641), .C1(n_1644), .C2(n_1646), .Y(n_1638) );
INVx2_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
OR2x2_ASAP7_75t_L g1640 ( .A(n_1518), .B(n_1531), .Y(n_1640) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1519), .B(n_1523), .Y(n_1581) );
NAND2xp5_ASAP7_75t_L g1599 ( .A(n_1519), .B(n_1532), .Y(n_1599) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1519), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1520), .B(n_1523), .Y(n_1663) );
NAND2xp5_ASAP7_75t_L g1521 ( .A(n_1522), .B(n_1524), .Y(n_1521) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1522), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1522), .B(n_1539), .Y(n_1679) );
OR2x2_ASAP7_75t_L g1557 ( .A(n_1523), .B(n_1558), .Y(n_1557) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1523), .B(n_1572), .Y(n_1629) );
AND2x2_ASAP7_75t_L g1652 ( .A(n_1523), .B(n_1624), .Y(n_1652) );
O2A1O1Ixp33_ASAP7_75t_L g1664 ( .A1(n_1525), .A2(n_1665), .B(n_1666), .C(n_1667), .Y(n_1664) );
A2O1A1Ixp33_ASAP7_75t_L g1526 ( .A1(n_1527), .A2(n_1529), .B(n_1534), .C(n_1553), .Y(n_1526) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
NAND2xp5_ASAP7_75t_L g1556 ( .A(n_1528), .B(n_1557), .Y(n_1556) );
O2A1O1Ixp33_ASAP7_75t_L g1598 ( .A1(n_1528), .A2(n_1532), .B(n_1599), .C(n_1600), .Y(n_1598) );
NOR2xp33_ASAP7_75t_L g1604 ( .A(n_1528), .B(n_1605), .Y(n_1604) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1533), .Y(n_1530) );
NAND2xp5_ASAP7_75t_L g1603 ( .A(n_1531), .B(n_1566), .Y(n_1603) );
NAND2xp5_ASAP7_75t_L g1611 ( .A(n_1531), .B(n_1612), .Y(n_1611) );
INVx2_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
AOI321xp33_ASAP7_75t_L g1555 ( .A1(n_1532), .A2(n_1556), .A3(n_1560), .B1(n_1562), .B2(n_1564), .C(n_1573), .Y(n_1555) );
NAND2xp5_ASAP7_75t_L g1576 ( .A(n_1532), .B(n_1577), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1532), .B(n_1594), .Y(n_1593) );
NAND2xp5_ASAP7_75t_SL g1628 ( .A(n_1532), .B(n_1566), .Y(n_1628) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1533), .Y(n_1596) );
OAI211xp5_ASAP7_75t_SL g1534 ( .A1(n_1535), .A2(n_1537), .B(n_1541), .C(n_1545), .Y(n_1534) );
OAI22xp5_ASAP7_75t_L g1591 ( .A1(n_1535), .A2(n_1592), .B1(n_1595), .B2(n_1596), .Y(n_1591) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
A2O1A1Ixp33_ASAP7_75t_L g1626 ( .A1(n_1536), .A2(n_1627), .B(n_1629), .C(n_1630), .Y(n_1626) );
AOI31xp33_ASAP7_75t_L g1677 ( .A1(n_1537), .A2(n_1574), .A3(n_1678), .B(n_1680), .Y(n_1677) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1540), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_1539), .B(n_1559), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1539), .B(n_1569), .Y(n_1674) );
INVxp67_ASAP7_75t_L g1595 ( .A(n_1540), .Y(n_1595) );
INVxp67_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1544), .Y(n_1542) );
INVx2_ASAP7_75t_L g1625 ( .A(n_1545), .Y(n_1625) );
INVx3_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
INVx3_ASAP7_75t_L g1554 ( .A(n_1546), .Y(n_1554) );
CKINVDCx5p33_ASAP7_75t_R g1682 ( .A(n_1547), .Y(n_1682) );
OAI22xp33_ASAP7_75t_L g1548 ( .A1(n_1549), .A2(n_1550), .B1(n_1551), .B2(n_1552), .Y(n_1548) );
AOI21xp5_ASAP7_75t_L g1573 ( .A1(n_1558), .A2(n_1574), .B(n_1576), .Y(n_1573) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1560), .B(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
NOR2xp33_ASAP7_75t_L g1568 ( .A(n_1561), .B(n_1569), .Y(n_1568) );
OAI22xp33_ASAP7_75t_L g1564 ( .A1(n_1565), .A2(n_1567), .B1(n_1570), .B2(n_1571), .Y(n_1564) );
INVxp33_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
NAND2xp5_ASAP7_75t_L g1609 ( .A(n_1569), .B(n_1610), .Y(n_1609) );
NOR2xp33_ASAP7_75t_L g1636 ( .A(n_1569), .B(n_1637), .Y(n_1636) );
INVx2_ASAP7_75t_L g1660 ( .A(n_1569), .Y(n_1660) );
NAND2xp5_ASAP7_75t_L g1662 ( .A(n_1569), .B(n_1663), .Y(n_1662) );
NOR2xp33_ASAP7_75t_L g1681 ( .A(n_1569), .B(n_1642), .Y(n_1681) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1570), .Y(n_1597) );
A2O1A1Ixp33_ASAP7_75t_L g1606 ( .A1(n_1570), .A2(n_1607), .B(n_1608), .C(n_1613), .Y(n_1606) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
NOR2xp33_ASAP7_75t_L g1676 ( .A(n_1575), .B(n_1581), .Y(n_1676) );
AOI221xp5_ASAP7_75t_L g1617 ( .A1(n_1577), .A2(n_1586), .B1(n_1618), .B2(n_1619), .C(n_1621), .Y(n_1617) );
CKINVDCx5p33_ASAP7_75t_R g1656 ( .A(n_1577), .Y(n_1656) );
INVxp67_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVxp67_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1586), .Y(n_1583) );
NAND5xp2_ASAP7_75t_L g1587 ( .A(n_1588), .B(n_1601), .C(n_1606), .D(n_1617), .E(n_1626), .Y(n_1587) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
AOI22xp5_ASAP7_75t_L g1632 ( .A1(n_1597), .A2(n_1633), .B1(n_1635), .B2(n_1636), .Y(n_1632) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1605), .Y(n_1670) );
INVxp67_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1618), .Y(n_1666) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
OAI21xp33_ASAP7_75t_L g1621 ( .A1(n_1622), .A2(n_1623), .B(n_1625), .Y(n_1621) );
NOR2xp33_ASAP7_75t_L g1644 ( .A(n_1622), .B(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1628), .Y(n_1627) );
NAND5xp2_ASAP7_75t_L g1631 ( .A(n_1632), .B(n_1638), .C(n_1648), .D(n_1657), .E(n_1669), .Y(n_1631) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1634), .Y(n_1655) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1634), .Y(n_1673) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
NAND2xp5_ASAP7_75t_L g1649 ( .A(n_1650), .B(n_1651), .Y(n_1649) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
OR2x2_ASAP7_75t_L g1654 ( .A(n_1655), .B(n_1656), .Y(n_1654) );
INVxp67_ASAP7_75t_SL g1658 ( .A(n_1659), .Y(n_1658) );
INVxp67_ASAP7_75t_SL g1661 ( .A(n_1662), .Y(n_1661) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1668), .Y(n_1667) );
O2A1O1Ixp33_ASAP7_75t_L g1669 ( .A1(n_1670), .A2(n_1671), .B(n_1675), .C(n_1677), .Y(n_1669) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_1673), .B(n_1674), .Y(n_1672) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
INVxp67_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
AND4x1_ASAP7_75t_L g1686 ( .A(n_1687), .B(n_1705), .C(n_1725), .D(n_1732), .Y(n_1686) );
NAND4xp25_ASAP7_75t_L g1741 ( .A(n_1687), .B(n_1705), .C(n_1725), .D(n_1732), .Y(n_1741) );
OAI31xp33_ASAP7_75t_L g1687 ( .A1(n_1688), .A2(n_1697), .A3(n_1700), .B(n_1704), .Y(n_1687) );
NAND3xp33_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1693), .C(n_1696), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1689 ( .A(n_1690), .B(n_1691), .Y(n_1689) );
INVx2_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
AO21x1_ASAP7_75t_SL g1705 ( .A1(n_1706), .A2(n_1717), .B(n_1724), .Y(n_1705) );
NOR3xp33_ASAP7_75t_L g1706 ( .A(n_1707), .B(n_1711), .C(n_1714), .Y(n_1706) );
INVx2_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
AND2x4_ASAP7_75t_L g1721 ( .A(n_1713), .B(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
AOI22xp5_ASAP7_75t_L g1717 ( .A1(n_1718), .A2(n_1719), .B1(n_1720), .B2(n_1721), .Y(n_1717) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1723), .Y(n_1722) );
CKINVDCx14_ASAP7_75t_R g1742 ( .A(n_1743), .Y(n_1742) );
INVx4_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
HB1xp67_ASAP7_75t_SL g1749 ( .A(n_1750), .Y(n_1749) );
A2O1A1Ixp33_ASAP7_75t_L g1800 ( .A1(n_1751), .A2(n_1801), .B(n_1803), .C(n_1804), .Y(n_1800) );
INVxp33_ASAP7_75t_SL g1752 ( .A(n_1753), .Y(n_1752) );
HB1xp67_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
NOR2x1_ASAP7_75t_L g1755 ( .A(n_1756), .B(n_1774), .Y(n_1755) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
HB1xp67_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
NAND4xp25_ASAP7_75t_L g1774 ( .A(n_1775), .B(n_1778), .C(n_1781), .D(n_1784), .Y(n_1774) );
INVx2_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
INVx1_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
HB1xp67_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1802), .Y(n_1801) );
endmodule