module fake_ariane_1381_n_909 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_909);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_909;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_670;
wire n_607;
wire n_897;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_761;
wire n_818;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_218;
wire n_839;
wire n_770;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_362;
wire n_260;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_639;
wire n_452;
wire n_217;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_872;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_136),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_24),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_10),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_145),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_132),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_185),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_71),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_98),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_50),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_86),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_26),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_75),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_65),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_22),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_99),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_42),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_102),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_76),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_52),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_16),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_32),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_90),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

BUFx8_ASAP7_75t_SL g223 ( 
.A(n_121),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_150),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_3),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_164),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_36),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_66),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_17),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_162),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_189),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_175),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_56),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_16),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_38),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_100),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_134),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_18),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_126),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_128),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_174),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_2),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_139),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_37),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_0),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_111),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_142),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_165),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_146),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_88),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_79),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_152),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_107),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_122),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_2),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_69),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_91),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_130),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_151),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_96),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_60),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_94),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_54),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_0),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_143),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_51),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_19),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_140),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_192),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_118),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_109),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_39),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_129),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_83),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_125),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_97),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_1),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_195),
.B(n_1),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_3),
.Y(n_282)
);

AND2x6_ASAP7_75t_L g283 ( 
.A(n_212),
.B(n_20),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

AND2x4_ASAP7_75t_L g285 ( 
.A(n_225),
.B(n_4),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_212),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_214),
.A2(n_101),
.B(n_193),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_199),
.Y(n_289)
);

AOI22x1_ASAP7_75t_SL g290 ( 
.A1(n_200),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_219),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_197),
.B(n_21),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_198),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_220),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

OA21x2_ASAP7_75t_L g298 ( 
.A1(n_203),
.A2(n_5),
.B(n_6),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_208),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_196),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_213),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_237),
.B(n_275),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_200),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_234),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_210),
.Y(n_307)
);

BUFx8_ASAP7_75t_SL g308 ( 
.A(n_223),
.Y(n_308)
);

BUFx8_ASAP7_75t_SL g309 ( 
.A(n_223),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_236),
.Y(n_310)
);

BUFx8_ASAP7_75t_L g311 ( 
.A(n_204),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_238),
.Y(n_312)
);

OAI22x1_ASAP7_75t_SL g313 ( 
.A1(n_215),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_201),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_240),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_241),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_242),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_246),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_235),
.Y(n_320)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_243),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_256),
.B(n_10),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_244),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_259),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_264),
.Y(n_329)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_265),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_267),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

BUFx8_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_202),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_205),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_R g338 ( 
.A(n_330),
.B(n_265),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_308),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_308),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_286),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_309),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_309),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_337),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_300),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_300),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_315),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_307),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_315),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_307),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_218),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_291),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_284),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_288),
.Y(n_357)
);

NAND2xp33_ASAP7_75t_SL g358 ( 
.A(n_282),
.B(n_215),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_288),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_326),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_311),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_284),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_307),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_288),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_276),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_311),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_284),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_334),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_334),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_280),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_280),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_327),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_296),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_320),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_316),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_321),
.B(n_207),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_325),
.Y(n_378)
);

AO21x2_ASAP7_75t_L g379 ( 
.A1(n_279),
.A2(n_211),
.B(n_209),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_324),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_296),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_297),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_330),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_295),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_295),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_297),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_297),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_303),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_303),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_317),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_303),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_R g392 ( 
.A(n_330),
.B(n_206),
.Y(n_392)
);

NOR2x1_ASAP7_75t_L g393 ( 
.A(n_317),
.B(n_224),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_313),
.B(n_224),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_306),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_321),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_350),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_341),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_361),
.B(n_321),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_346),
.B(n_321),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_353),
.B(n_325),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_354),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_379),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_340),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_379),
.B(n_302),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_341),
.B(n_302),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_390),
.B(n_279),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_345),
.B(n_285),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_376),
.Y(n_411)
);

NAND3xp33_ASAP7_75t_L g412 ( 
.A(n_366),
.B(n_281),
.C(n_285),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_356),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_348),
.B(n_301),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_357),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_358),
.A2(n_273),
.B1(n_304),
.B2(n_281),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_357),
.B(n_314),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_364),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_380),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_349),
.B(n_318),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_365),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

BUFx6f_ASAP7_75t_SL g426 ( 
.A(n_339),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_351),
.B(n_319),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_387),
.B(n_328),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_333),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_389),
.B(n_306),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_391),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_371),
.B(n_372),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_306),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_384),
.B(n_294),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_362),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

NAND3xp33_ASAP7_75t_L g439 ( 
.A(n_385),
.B(n_375),
.C(n_373),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_360),
.B(n_292),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_395),
.B(n_299),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_378),
.B(n_305),
.Y(n_442)
);

INVxp33_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_396),
.B(n_310),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_386),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_378),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_393),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_338),
.B(n_304),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_338),
.B(n_329),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_392),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_377),
.B(n_331),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_SL g454 ( 
.A(n_342),
.B(n_273),
.C(n_292),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_367),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_369),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_392),
.B(n_312),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_370),
.B(n_312),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_352),
.B(n_312),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_363),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_344),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_354),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_353),
.B(n_322),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_346),
.B(n_322),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_341),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_346),
.B(n_283),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_407),
.Y(n_468)
);

NOR2x1p5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_313),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_397),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_407),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_401),
.A2(n_293),
.B1(n_216),
.B2(n_254),
.Y(n_472)
);

NOR3xp33_ASAP7_75t_SL g473 ( 
.A(n_454),
.B(n_290),
.C(n_221),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_293),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_401),
.A2(n_260),
.B1(n_222),
.B2(n_226),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_428),
.B(n_322),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_440),
.B(n_289),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_323),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_448),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_419),
.Y(n_481)
);

BUFx8_ASAP7_75t_SL g482 ( 
.A(n_426),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_323),
.Y(n_483)
);

NAND2x1p5_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_323),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_419),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_411),
.B(n_332),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_429),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_332),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_436),
.B(n_332),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_403),
.A2(n_252),
.B1(n_227),
.B2(n_228),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_429),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_404),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_421),
.B(n_217),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_461),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_449),
.B(n_409),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_414),
.B(n_289),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_438),
.B(n_298),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_456),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_422),
.B(n_231),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_403),
.A2(n_262),
.B1(n_233),
.B2(n_245),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_442),
.B(n_283),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_434),
.B(n_450),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_426),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_456),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_456),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_412),
.A2(n_268),
.B1(n_248),
.B2(n_249),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_402),
.B(n_463),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_398),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_439),
.B(n_232),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_451),
.B(n_283),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_416),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_458),
.B(n_283),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_457),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_406),
.A2(n_298),
.B1(n_270),
.B2(n_277),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_455),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_430),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_418),
.A2(n_250),
.B1(n_261),
.B2(n_263),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_430),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_458),
.B(n_271),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_405),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_462),
.B(n_11),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_406),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_444),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_405),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_408),
.A2(n_287),
.B1(n_12),
.B2(n_13),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_405),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_417),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_437),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_460),
.B(n_11),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_435),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_445),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_431),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_441),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_453),
.B(n_12),
.Y(n_535)
);

INVx6_ASAP7_75t_L g536 ( 
.A(n_399),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_SL g537 ( 
.A(n_400),
.B(n_13),
.C(n_14),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_413),
.B(n_14),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_435),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_507),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_531),
.Y(n_541)
);

OAI221xp5_ASAP7_75t_L g542 ( 
.A1(n_478),
.A2(n_496),
.B1(n_518),
.B2(n_530),
.C(n_522),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_508),
.Y(n_543)
);

A2O1A1Ixp33_ASAP7_75t_L g544 ( 
.A1(n_468),
.A2(n_467),
.B(n_415),
.C(n_424),
.Y(n_544)
);

OAI21xp33_ASAP7_75t_L g545 ( 
.A1(n_476),
.A2(n_441),
.B(n_423),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_523),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_509),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_474),
.B(n_459),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_471),
.B(n_534),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_502),
.B(n_420),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_539),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_502),
.B(n_427),
.Y(n_552)
);

AOI21x1_ASAP7_75t_L g553 ( 
.A1(n_513),
.A2(n_466),
.B(n_433),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_470),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_512),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_498),
.B(n_431),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_481),
.A2(n_447),
.B1(n_446),
.B2(n_432),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_499),
.A2(n_425),
.B(n_114),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_494),
.Y(n_559)
);

CKINVDCx14_ASAP7_75t_R g560 ( 
.A(n_492),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_528),
.Y(n_561)
);

O2A1O1Ixp5_ASAP7_75t_L g562 ( 
.A1(n_510),
.A2(n_15),
.B(n_17),
.C(n_23),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_482),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g564 ( 
.A(n_503),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_R g565 ( 
.A(n_495),
.B(n_443),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_474),
.B(n_15),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_485),
.B(n_25),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_487),
.A2(n_519),
.B1(n_517),
.B2(n_491),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_495),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_490),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_498),
.B(n_34),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_500),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_472),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_511),
.A2(n_46),
.B(n_47),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_479),
.Y(n_575)
);

A2O1A1Ixp33_ASAP7_75t_SL g576 ( 
.A1(n_538),
.A2(n_194),
.B(n_49),
.C(n_53),
.Y(n_576)
);

OAI221xp5_ASAP7_75t_L g577 ( 
.A1(n_480),
.A2(n_48),
.B1(n_55),
.B2(n_57),
.C(n_58),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_524),
.B(n_59),
.Y(n_578)
);

AOI21x1_ASAP7_75t_L g579 ( 
.A1(n_501),
.A2(n_61),
.B(n_62),
.Y(n_579)
);

A2O1A1Ixp33_ASAP7_75t_L g580 ( 
.A1(n_477),
.A2(n_63),
.B(n_64),
.C(n_67),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_504),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_514),
.B(n_504),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_520),
.A2(n_68),
.B(n_70),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_533),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_483),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_516),
.Y(n_586)
);

AOI21x1_ASAP7_75t_L g587 ( 
.A1(n_488),
.A2(n_72),
.B(n_73),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_505),
.B(n_74),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_505),
.B(n_77),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_529),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_527),
.B(n_78),
.Y(n_591)
);

A2O1A1Ixp33_ASAP7_75t_SL g592 ( 
.A1(n_535),
.A2(n_191),
.B(n_81),
.C(n_82),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_497),
.Y(n_593)
);

NAND2x1p5_ASAP7_75t_L g594 ( 
.A(n_521),
.B(n_80),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_515),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_595)
);

NOR2xp67_ASAP7_75t_L g596 ( 
.A(n_521),
.B(n_89),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_489),
.B(n_92),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_475),
.B(n_93),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_475),
.B(n_95),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_533),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_553),
.A2(n_526),
.B(n_484),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_549),
.A2(n_506),
.B(n_493),
.Y(n_602)
);

NAND2x1p5_ASAP7_75t_L g603 ( 
.A(n_581),
.B(n_532),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_584),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_540),
.B(n_475),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_532),
.Y(n_606)
);

AO21x2_ASAP7_75t_L g607 ( 
.A1(n_544),
.A2(n_486),
.B(n_537),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_554),
.B(n_469),
.Y(n_608)
);

AO21x2_ASAP7_75t_L g609 ( 
.A1(n_567),
.A2(n_475),
.B(n_533),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_568),
.A2(n_525),
.B(n_532),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_582),
.B(n_473),
.Y(n_611)
);

BUFx12f_ASAP7_75t_L g612 ( 
.A(n_563),
.Y(n_612)
);

BUFx8_ASAP7_75t_L g613 ( 
.A(n_564),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_579),
.A2(n_536),
.B(n_105),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_543),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_574),
.A2(n_536),
.B(n_108),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_559),
.B(n_541),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_560),
.Y(n_618)
);

OAI21x1_ASAP7_75t_L g619 ( 
.A1(n_587),
.A2(n_104),
.B(n_110),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_551),
.B(n_112),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_597),
.A2(n_113),
.B(n_115),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_547),
.Y(n_622)
);

AO21x2_ASAP7_75t_L g623 ( 
.A1(n_575),
.A2(n_117),
.B(n_119),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_542),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_581),
.Y(n_625)
);

AOI22x1_ASAP7_75t_L g626 ( 
.A1(n_558),
.A2(n_127),
.B1(n_131),
.B2(n_133),
.Y(n_626)
);

INVx5_ASAP7_75t_L g627 ( 
.A(n_584),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_555),
.Y(n_628)
);

AOI22x1_ASAP7_75t_L g629 ( 
.A1(n_583),
.A2(n_137),
.B1(n_138),
.B2(n_141),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_561),
.Y(n_630)
);

NAND2x1p5_ASAP7_75t_L g631 ( 
.A(n_584),
.B(n_144),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_585),
.A2(n_148),
.B(n_149),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_594),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_590),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_548),
.B(n_153),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_586),
.Y(n_636)
);

INVxp67_ASAP7_75t_SL g637 ( 
.A(n_546),
.Y(n_637)
);

AO21x2_ASAP7_75t_L g638 ( 
.A1(n_593),
.A2(n_154),
.B(n_155),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_600),
.Y(n_639)
);

NAND2x1p5_ASAP7_75t_L g640 ( 
.A(n_588),
.B(n_156),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_548),
.B(n_190),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_545),
.A2(n_157),
.B(n_158),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_591),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_550),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_598),
.A2(n_160),
.B(n_161),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_589),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_599),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_552),
.B(n_163),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_566),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_615),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_622),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_630),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_622),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_624),
.A2(n_648),
.B1(n_642),
.B2(n_602),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_628),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_636),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_628),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_637),
.Y(n_658)
);

NAND2x1p5_ASAP7_75t_L g659 ( 
.A(n_627),
.B(n_596),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_637),
.B(n_545),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_644),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_634),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_646),
.A2(n_578),
.B1(n_569),
.B2(n_595),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_644),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_605),
.B(n_556),
.Y(n_665)
);

AOI21x1_ASAP7_75t_L g666 ( 
.A1(n_601),
.A2(n_596),
.B(n_573),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_635),
.A2(n_571),
.B1(n_570),
.B2(n_572),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_620),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_612),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_617),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_646),
.A2(n_557),
.B1(n_577),
.B2(n_580),
.Y(n_671)
);

AOI21x1_ASAP7_75t_L g672 ( 
.A1(n_601),
.A2(n_576),
.B(n_556),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_636),
.Y(n_673)
);

AOI21x1_ASAP7_75t_L g674 ( 
.A1(n_614),
.A2(n_592),
.B(n_571),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_608),
.B(n_565),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_614),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_618),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_619),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_639),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_619),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_632),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_639),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_612),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_SL g684 ( 
.A1(n_635),
.A2(n_562),
.B1(n_168),
.B2(n_169),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_610),
.B(n_166),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_635),
.B(n_170),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_632),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_608),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_624),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_689)
);

NAND2x1p5_ASAP7_75t_L g690 ( 
.A(n_627),
.B(n_176),
.Y(n_690)
);

CKINVDCx6p67_ASAP7_75t_R g691 ( 
.A(n_618),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_625),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_R g693 ( 
.A(n_669),
.B(n_613),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_683),
.Y(n_694)
);

CKINVDCx16_ASAP7_75t_R g695 ( 
.A(n_673),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_658),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_SL g697 ( 
.A1(n_654),
.A2(n_640),
.B(n_649),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_L g698 ( 
.A(n_654),
.B(n_640),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_650),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_670),
.B(n_611),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_658),
.B(n_608),
.Y(n_701)
);

BUFx12f_ASAP7_75t_L g702 ( 
.A(n_656),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_662),
.B(n_604),
.Y(n_703)
);

CKINVDCx16_ASAP7_75t_R g704 ( 
.A(n_673),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_R g705 ( 
.A(n_691),
.B(n_613),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_688),
.B(n_668),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_660),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_677),
.Y(n_708)
);

OR2x2_ASAP7_75t_SL g709 ( 
.A(n_679),
.B(n_613),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_667),
.A2(n_648),
.B1(n_641),
.B2(n_643),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_682),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_SL g712 ( 
.A(n_689),
.B(n_603),
.C(n_631),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_661),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_675),
.B(n_604),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_652),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_R g716 ( 
.A(n_692),
.B(n_643),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_661),
.B(n_604),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_692),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_686),
.Y(n_719)
);

CKINVDCx9p33_ASAP7_75t_R g720 ( 
.A(n_665),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_686),
.B(n_648),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_657),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_686),
.B(n_606),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_692),
.Y(n_724)
);

XNOR2xp5_ASAP7_75t_L g725 ( 
.A(n_664),
.B(n_606),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_692),
.Y(n_726)
);

OAI21x1_ASAP7_75t_SL g727 ( 
.A1(n_689),
.A2(n_674),
.B(n_663),
.Y(n_727)
);

CKINVDCx16_ASAP7_75t_R g728 ( 
.A(n_665),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_651),
.B(n_609),
.Y(n_729)
);

AO31x2_ASAP7_75t_L g730 ( 
.A1(n_676),
.A2(n_609),
.A3(n_638),
.B(n_623),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_651),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_SL g732 ( 
.A(n_684),
.B(n_603),
.C(n_631),
.Y(n_732)
);

AO32x1_ASAP7_75t_L g733 ( 
.A1(n_681),
.A2(n_625),
.A3(n_638),
.B1(n_623),
.B2(n_607),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_653),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_653),
.A2(n_647),
.B1(n_607),
.B2(n_633),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_655),
.Y(n_736)
);

CKINVDCx9p33_ASAP7_75t_R g737 ( 
.A(n_655),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_676),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_671),
.Y(n_739)
);

AND2x2_ASAP7_75t_SL g740 ( 
.A(n_685),
.B(n_625),
.Y(n_740)
);

AO31x2_ASAP7_75t_L g741 ( 
.A1(n_681),
.A2(n_647),
.A3(n_616),
.B(n_621),
.Y(n_741)
);

INVx5_ASAP7_75t_L g742 ( 
.A(n_687),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_685),
.B(n_633),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_699),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_728),
.B(n_687),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_707),
.B(n_627),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_701),
.B(n_680),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_715),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_707),
.B(n_680),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_706),
.B(n_739),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_713),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_722),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_696),
.B(n_678),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_696),
.B(n_678),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_711),
.B(n_690),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_703),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_700),
.B(n_690),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_702),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_713),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_SL g760 ( 
.A(n_716),
.B(n_633),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_734),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_714),
.B(n_627),
.Y(n_762)
);

OAI21x1_ASAP7_75t_L g763 ( 
.A1(n_727),
.A2(n_672),
.B(n_666),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_742),
.B(n_721),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_742),
.B(n_645),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_742),
.B(n_645),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_695),
.B(n_606),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_734),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_741),
.Y(n_769)
);

AO31x2_ASAP7_75t_L g770 ( 
.A1(n_738),
.A2(n_616),
.A3(n_621),
.B(n_629),
.Y(n_770)
);

INVx3_ASAP7_75t_SL g771 ( 
.A(n_694),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_693),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_704),
.B(n_659),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_719),
.B(n_659),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_717),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_731),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_743),
.Y(n_777)
);

NOR2xp67_ASAP7_75t_SL g778 ( 
.A(n_697),
.B(n_626),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_718),
.B(n_177),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_709),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_725),
.B(n_178),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_724),
.Y(n_782)
);

INVxp67_ASAP7_75t_SL g783 ( 
.A(n_729),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_723),
.B(n_179),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_710),
.B(n_180),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_752),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_751),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_751),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_756),
.B(n_708),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_760),
.B(n_740),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_768),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_744),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_760),
.B(n_726),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_775),
.B(n_698),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_753),
.B(n_741),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_753),
.B(n_741),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_754),
.B(n_735),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_777),
.B(n_736),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_765),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_782),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_754),
.B(n_730),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_745),
.B(n_712),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_764),
.B(n_750),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_764),
.B(n_730),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_748),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_755),
.B(n_732),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_768),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_759),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_749),
.B(n_747),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_755),
.B(n_705),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_761),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_749),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_787),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_787),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_799),
.B(n_780),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_800),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_808),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_788),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_809),
.B(n_783),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_786),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_792),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_803),
.B(n_758),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_812),
.B(n_765),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_809),
.B(n_773),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_788),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_799),
.B(n_795),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_789),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_795),
.Y(n_828)
);

OAI22xp33_ASAP7_75t_SL g829 ( 
.A1(n_806),
.A2(n_781),
.B1(n_785),
.B2(n_767),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_815),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_815),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_813),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_819),
.B(n_798),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_816),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_817),
.B(n_811),
.Y(n_835)
);

OA222x2_ASAP7_75t_L g836 ( 
.A1(n_828),
.A2(n_794),
.B1(n_802),
.B2(n_799),
.C1(n_790),
.C2(n_793),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_829),
.B(n_790),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_813),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_827),
.B(n_771),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_827),
.B(n_773),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_832),
.Y(n_841)
);

XOR2xp5_ASAP7_75t_L g842 ( 
.A(n_837),
.B(n_772),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_840),
.A2(n_828),
.B1(n_757),
.B2(n_797),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_840),
.A2(n_836),
.B1(n_834),
.B2(n_839),
.Y(n_844)
);

AOI21xp33_ASAP7_75t_SL g845 ( 
.A1(n_830),
.A2(n_771),
.B(n_772),
.Y(n_845)
);

AOI21xp33_ASAP7_75t_L g846 ( 
.A1(n_835),
.A2(n_821),
.B(n_820),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_846),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_841),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_842),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_843),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_844),
.B(n_810),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_845),
.A2(n_793),
.B(n_817),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_847),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_848),
.Y(n_854)
);

NAND3xp33_ASAP7_75t_SL g855 ( 
.A(n_849),
.B(n_852),
.C(n_850),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_L g856 ( 
.A(n_851),
.B(n_784),
.C(n_823),
.Y(n_856)
);

NOR2x1_ASAP7_75t_L g857 ( 
.A(n_855),
.B(n_831),
.Y(n_857)
);

NOR3xp33_ASAP7_75t_L g858 ( 
.A(n_853),
.B(n_784),
.C(n_779),
.Y(n_858)
);

AOI221xp5_ASAP7_75t_L g859 ( 
.A1(n_858),
.A2(n_854),
.B1(n_856),
.B2(n_857),
.C(n_778),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_858),
.B(n_822),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_857),
.B(n_831),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_860),
.B(n_830),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_861),
.Y(n_863)
);

INVxp33_ASAP7_75t_SL g864 ( 
.A(n_859),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_861),
.Y(n_865)
);

INVxp33_ASAP7_75t_SL g866 ( 
.A(n_861),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_859),
.B(n_826),
.Y(n_867)
);

NOR3xp33_ASAP7_75t_L g868 ( 
.A(n_865),
.B(n_779),
.C(n_757),
.Y(n_868)
);

NOR2x1_ASAP7_75t_L g869 ( 
.A(n_863),
.B(n_779),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_864),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_862),
.Y(n_871)
);

OAI221xp5_ASAP7_75t_L g872 ( 
.A1(n_867),
.A2(n_833),
.B1(n_823),
.B2(n_805),
.C(n_746),
.Y(n_872)
);

NOR2xp67_ASAP7_75t_L g873 ( 
.A(n_866),
.B(n_824),
.Y(n_873)
);

NAND4xp75_ASAP7_75t_L g874 ( 
.A(n_863),
.B(n_762),
.C(n_720),
.D(n_766),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_873),
.Y(n_875)
);

NAND2xp33_ASAP7_75t_L g876 ( 
.A(n_871),
.B(n_838),
.Y(n_876)
);

NOR2xp67_ASAP7_75t_L g877 ( 
.A(n_870),
.B(n_826),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_869),
.B(n_796),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_874),
.Y(n_879)
);

NAND4xp25_ASAP7_75t_L g880 ( 
.A(n_872),
.B(n_766),
.C(n_797),
.D(n_774),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_868),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_875),
.Y(n_882)
);

OA22x2_ASAP7_75t_L g883 ( 
.A1(n_881),
.A2(n_763),
.B1(n_818),
.B2(n_814),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_879),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_876),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_877),
.A2(n_769),
.B1(n_818),
.B2(n_825),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_878),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_880),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_875),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_875),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_887),
.A2(n_796),
.B1(n_804),
.B2(n_801),
.Y(n_891)
);

BUFx4f_ASAP7_75t_SL g892 ( 
.A(n_882),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_889),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_890),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_888),
.A2(n_804),
.B1(n_801),
.B2(n_774),
.Y(n_895)
);

AOI31xp33_ASAP7_75t_L g896 ( 
.A1(n_884),
.A2(n_737),
.A3(n_807),
.B(n_791),
.Y(n_896)
);

AOI31xp33_ASAP7_75t_L g897 ( 
.A1(n_885),
.A2(n_791),
.A3(n_807),
.B(n_184),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_883),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_886),
.B(n_181),
.Y(n_899)
);

OAI22x1_ASAP7_75t_SL g900 ( 
.A1(n_893),
.A2(n_182),
.B1(n_186),
.B2(n_187),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_892),
.B(n_769),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_894),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_898),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_903),
.A2(n_899),
.B1(n_895),
.B2(n_891),
.Y(n_904)
);

XNOR2x1_ASAP7_75t_L g905 ( 
.A(n_901),
.B(n_897),
.Y(n_905)
);

NOR2xp67_ASAP7_75t_SL g906 ( 
.A(n_905),
.B(n_902),
.Y(n_906)
);

AOI222xp33_ASAP7_75t_L g907 ( 
.A1(n_906),
.A2(n_900),
.B1(n_904),
.B2(n_896),
.C1(n_769),
.C2(n_776),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_907),
.B(n_188),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_908),
.A2(n_763),
.B1(n_733),
.B2(n_770),
.Y(n_909)
);


endmodule