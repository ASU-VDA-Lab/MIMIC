module fake_jpeg_20001_n_292 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_265;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_8),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_29),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_37),
.Y(n_94)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_25),
.B1(n_19),
.B2(n_26),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_61),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_25),
.B1(n_19),
.B2(n_26),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_25),
.B1(n_19),
.B2(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_32),
.B1(n_25),
.B2(n_33),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_17),
.B1(n_21),
.B2(n_20),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_31),
.B1(n_22),
.B2(n_23),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_39),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_31),
.B1(n_23),
.B2(n_33),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_68),
.A2(n_51),
.B1(n_49),
.B2(n_47),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_40),
.B1(n_38),
.B2(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_39),
.B(n_40),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_94),
.B(n_21),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_34),
.B1(n_20),
.B2(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_20),
.B1(n_34),
.B2(n_21),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_46),
.B1(n_61),
.B2(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_41),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_33),
.B(n_32),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_95),
.B(n_50),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_34),
.B1(n_20),
.B2(n_21),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_49),
.B1(n_58),
.B2(n_60),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_42),
.B1(n_37),
.B2(n_17),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_47),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_84),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_17),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_91),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_60),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_90),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_114),
.B1(n_95),
.B2(n_94),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_48),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_115),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_51),
.B1(n_49),
.B2(n_52),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_89),
.B1(n_81),
.B2(n_93),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_17),
.A3(n_28),
.B1(n_34),
.B2(n_27),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_116),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_123),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_124),
.B1(n_74),
.B2(n_80),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_27),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_27),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_28),
.B(n_1),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_81),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_28),
.B1(n_1),
.B2(n_2),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_127),
.B1(n_145),
.B2(n_114),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_126),
.A2(n_135),
.B1(n_146),
.B2(n_149),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_113),
.A2(n_66),
.B1(n_73),
.B2(n_69),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_82),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_129),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_94),
.B1(n_66),
.B2(n_83),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_98),
.B(n_78),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_137),
.B(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_142),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_98),
.B(n_76),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_86),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_96),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_147),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_82),
.B1(n_91),
.B2(n_92),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_65),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_77),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_154),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_65),
.B1(n_77),
.B2(n_67),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_67),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_112),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_9),
.C(n_15),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_14),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_77),
.A3(n_72),
.B1(n_14),
.B2(n_13),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_9),
.Y(n_179)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_14),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_107),
.B(n_117),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_175),
.B(n_184),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_156),
.A2(n_170),
.B1(n_179),
.B2(n_11),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_157),
.B(n_154),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_115),
.C(n_108),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_162),
.C(n_180),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_115),
.C(n_108),
.Y(n_162)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_141),
.B(n_106),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_169),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_102),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_108),
.B1(n_115),
.B2(n_110),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_121),
.B(n_99),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_177),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_102),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_101),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_181),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_101),
.C(n_111),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_119),
.B1(n_99),
.B2(n_111),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_128),
.B1(n_148),
.B2(n_134),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_127),
.B(n_13),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_152),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_72),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_137),
.B(n_140),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_170),
.B1(n_164),
.B2(n_168),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_144),
.B(n_134),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_192),
.B(n_201),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_130),
.C(n_132),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_200),
.C(n_202),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_126),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_199),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_128),
.C(n_146),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_129),
.C(n_147),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_206),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_149),
.C(n_145),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_205),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_153),
.C(n_11),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_163),
.B(n_11),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_155),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_191),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_183),
.B1(n_167),
.B2(n_159),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_197),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_211),
.B(n_224),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_191),
.A2(n_165),
.B1(n_171),
.B2(n_182),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_214),
.B1(n_219),
.B2(n_220),
.Y(n_236)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_215),
.A2(n_229),
.B1(n_176),
.B2(n_181),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_167),
.B1(n_158),
.B2(n_156),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_158),
.B1(n_164),
.B2(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_159),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_169),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_230),
.C(n_226),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_237),
.C(n_238),
.Y(n_252)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_199),
.B(n_194),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_223),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_233),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_193),
.C(n_204),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_202),
.C(n_200),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_207),
.C(n_190),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_240),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_209),
.C(n_186),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_209),
.C(n_205),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_0),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_219),
.A2(n_179),
.B1(n_209),
.B2(n_172),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_236),
.B1(n_217),
.B2(n_239),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_178),
.B(n_177),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_212),
.B(n_227),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_245),
.B(n_3),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_220),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_172),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_214),
.B(n_225),
.C(n_215),
.Y(n_250)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_250),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_257),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_255),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_210),
.B1(n_213),
.B2(n_10),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_238),
.CI(n_236),
.CON(n_256),
.SN(n_256)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_258),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_10),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_3),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_231),
.C(n_245),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_261),
.Y(n_272)
);

AOI31xp67_ASAP7_75t_SL g261 ( 
.A1(n_255),
.A2(n_243),
.A3(n_241),
.B(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_258),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_2),
.C(n_3),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_266),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_4),
.B(n_5),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_4),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_248),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_273),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_256),
.C(n_253),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_276),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_270),
.Y(n_276)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_249),
.B(n_264),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_256),
.C(n_254),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_265),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_247),
.CI(n_264),
.CON(n_279),
.SN(n_279)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_283),
.C(n_250),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_250),
.B(n_5),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_284),
.A2(n_4),
.B(n_6),
.Y(n_288)
);

OAI321xp33_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_287),
.A3(n_288),
.B1(n_279),
.B2(n_282),
.C(n_281),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_274),
.C(n_250),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_6),
.C(n_7),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_290),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_7),
.Y(n_292)
);


endmodule