module fake_jpeg_18655_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_37),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_15),
.B(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_43),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_32),
.B1(n_21),
.B2(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_45),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_51),
.B1(n_58),
.B2(n_16),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_33),
.B1(n_24),
.B2(n_20),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_55),
.B1(n_56),
.B2(n_61),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_33),
.B1(n_24),
.B2(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_57),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_33),
.B1(n_24),
.B2(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_24),
.B1(n_20),
.B2(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_29),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_32),
.B1(n_21),
.B2(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_61),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_62),
.B(n_63),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_61),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_74),
.Y(n_109)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_23),
.B1(n_15),
.B2(n_43),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_77),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_82),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_45),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_46),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_44),
.B1(n_36),
.B2(n_21),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_90),
.B1(n_59),
.B2(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_23),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_83),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_23),
.B1(n_44),
.B2(n_36),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_87),
.B1(n_89),
.B2(n_93),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_56),
.A2(n_36),
.B1(n_44),
.B2(n_16),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_32),
.B1(n_16),
.B2(n_22),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_45),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_92),
.CI(n_45),
.CON(n_98),
.SN(n_98)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_45),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_22),
.B1(n_30),
.B2(n_58),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_30),
.Y(n_94)
);

AND2x4_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_35),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_98),
.B(n_102),
.Y(n_143)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_122),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_108),
.B1(n_96),
.B2(n_94),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_35),
.Y(n_102)
);

OAI21x1_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_91),
.B(n_74),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_59),
.B1(n_39),
.B2(n_18),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_62),
.A2(n_18),
.B1(n_31),
.B2(n_19),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_124),
.B1(n_126),
.B2(n_95),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_65),
.A2(n_39),
.B1(n_18),
.B2(n_47),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_65),
.A2(n_39),
.B1(n_18),
.B2(n_47),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_79),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_151),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_141),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_106),
.B1(n_103),
.B2(n_124),
.Y(n_154)
);

XNOR2x1_ASAP7_75t_SL g171 ( 
.A(n_135),
.B(n_98),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_63),
.B(n_91),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_144),
.B(n_106),
.Y(n_160)
);

AOI21x1_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_75),
.B(n_66),
.Y(n_137)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_64),
.B1(n_80),
.B2(n_67),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_72),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_86),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_153),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_116),
.B(n_102),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_94),
.B1(n_87),
.B2(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_82),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_73),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_92),
.C(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_154),
.B(n_168),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_108),
.B1(n_118),
.B2(n_101),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_173),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_163),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_160),
.A2(n_145),
.B(n_133),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_111),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_167),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_78),
.C(n_70),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_149),
.Y(n_168)
);

OAI21x1_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_155),
.B(n_162),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_114),
.B1(n_126),
.B2(n_90),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_129),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_179),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_114),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_80),
.B1(n_64),
.B2(n_71),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_176),
.A2(n_138),
.B1(n_130),
.B2(n_142),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_129),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_184),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_18),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_182),
.C(n_133),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_18),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_115),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_143),
.B(n_144),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_187),
.B(n_189),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_143),
.B(n_137),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_137),
.B(n_139),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_201),
.B(n_203),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_200),
.B1(n_210),
.B2(n_125),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_85),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_148),
.C(n_145),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_198),
.C(n_182),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_145),
.C(n_135),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_145),
.B1(n_134),
.B2(n_141),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_178),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_104),
.B(n_100),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_169),
.B(n_150),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_177),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

FAx1_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_85),
.CI(n_88),
.CON(n_207),
.SN(n_207)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_170),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_132),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_166),
.A2(n_152),
.B1(n_125),
.B2(n_99),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_215),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_154),
.B1(n_184),
.B2(n_156),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_231),
.B1(n_186),
.B2(n_189),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_181),
.C(n_173),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_220),
.C(n_222),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_170),
.C(n_159),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_183),
.C(n_178),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_201),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_225),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_176),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_183),
.C(n_161),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_228),
.C(n_230),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_107),
.C(n_67),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_229),
.A2(n_226),
.B1(n_208),
.B2(n_211),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_200),
.B(n_31),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_191),
.A2(n_11),
.B1(n_12),
.B2(n_10),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_232),
.B(n_185),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_207),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_248),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_190),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_191),
.B1(n_195),
.B2(n_199),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_240),
.B1(n_219),
.B2(n_207),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_199),
.B1(n_210),
.B2(n_205),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_216),
.B(n_194),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_244),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_204),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_246),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_188),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_251),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_224),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_220),
.C(n_222),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_258),
.C(n_259),
.Y(n_270)
);

NAND4xp25_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_192),
.C(n_207),
.D(n_227),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_256),
.A2(n_19),
.B(n_17),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_257),
.B(n_29),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_212),
.C(n_232),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_250),
.C(n_248),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_215),
.C(n_227),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_263),
.C(n_266),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_213),
.C(n_107),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_17),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_100),
.C(n_127),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_12),
.B(n_11),
.C(n_3),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_267),
.A2(n_246),
.B(n_235),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_0),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_238),
.B1(n_243),
.B2(n_236),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_271),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_243),
.B1(n_239),
.B2(n_4),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_100),
.B(n_11),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_274),
.B(n_277),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_17),
.C(n_29),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_260),
.C(n_258),
.Y(n_280)
);

NAND4xp25_ASAP7_75t_SL g276 ( 
.A(n_267),
.B(n_31),
.C(n_19),
.D(n_29),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_278),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_261),
.B1(n_263),
.B2(n_259),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_273),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_282),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_262),
.C(n_266),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_0),
.B(n_2),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_276),
.B(n_5),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_269),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_0),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_288),
.B(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_278),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_291),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_293),
.B1(n_296),
.B2(n_7),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_270),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_295),
.A3(n_273),
.B1(n_275),
.B2(n_17),
.C1(n_7),
.C2(n_4),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_9),
.B(n_6),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_297),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_17),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_300),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_301),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_299),
.C(n_6),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_305),
.A2(n_306),
.B(n_303),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_302),
.A2(n_4),
.B(n_8),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_304),
.C(n_9),
.Y(n_308)
);


endmodule