module fake_jpeg_13283_n_299 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_1),
.Y(n_68)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_21),
.Y(n_71)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_19),
.B1(n_29),
.B2(n_20),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_33),
.B1(n_22),
.B2(n_19),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_46),
.A2(n_57),
.B1(n_58),
.B2(n_65),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_47),
.B(n_53),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_29),
.B(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_68),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_66),
.B1(n_43),
.B2(n_37),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_28),
.B1(n_26),
.B2(n_30),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_31),
.B1(n_26),
.B2(n_28),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_28),
.B1(n_26),
.B2(n_30),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_59),
.A2(n_61),
.B1(n_32),
.B2(n_7),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_18),
.B1(n_30),
.B2(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_3),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_18),
.B1(n_23),
.B2(n_17),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_18),
.B1(n_20),
.B2(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_40),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_27),
.B(n_21),
.C(n_32),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_32),
.B(n_7),
.C(n_8),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_78),
.B1(n_58),
.B2(n_46),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_75),
.B(n_82),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_40),
.B1(n_27),
.B2(n_21),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_95),
.Y(n_119)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_40),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_87),
.B(n_99),
.Y(n_131)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_90),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_62),
.B(n_5),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_105),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_5),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_98),
.Y(n_128)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_27),
.B1(n_32),
.B2(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_5),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_53),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_112),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_73),
.B1(n_71),
.B2(n_100),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_121),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_106),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_55),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_132),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g129 ( 
.A1(n_84),
.A2(n_72),
.A3(n_60),
.B1(n_49),
.B2(n_68),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_71),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_135),
.B(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_137),
.B(n_139),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_87),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_84),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_140),
.B(n_145),
.Y(n_195)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_152),
.Y(n_189)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_98),
.B(n_105),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_103),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_103),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_157),
.C(n_114),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_89),
.B1(n_105),
.B2(n_98),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_148),
.A2(n_156),
.B1(n_166),
.B2(n_6),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_89),
.B(n_95),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_160),
.B(n_133),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_91),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_91),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_120),
.B1(n_117),
.B2(n_126),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_85),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_163),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_109),
.A2(n_57),
.B1(n_65),
.B2(n_92),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_93),
.C(n_85),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_108),
.B(n_71),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_102),
.B(n_79),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_165),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_81),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_110),
.A2(n_77),
.B1(n_67),
.B2(n_83),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_164),
.A2(n_120),
.B1(n_117),
.B2(n_134),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_97),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_113),
.A2(n_76),
.B1(n_94),
.B2(n_83),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_137),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_180),
.C(n_159),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_151),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_148),
.A2(n_118),
.B1(n_134),
.B2(n_130),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_176),
.B(n_179),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_167),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_192),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_127),
.B(n_123),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_130),
.B(n_118),
.C(n_127),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_161),
.B(n_147),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_118),
.C(n_133),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_183),
.B1(n_188),
.B2(n_166),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_194),
.B1(n_165),
.B2(n_141),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_131),
.B1(n_117),
.B2(n_126),
.Y(n_183)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_107),
.B(n_9),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_149),
.B(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_155),
.A2(n_32),
.B1(n_9),
.B2(n_11),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_193),
.A2(n_144),
.B(n_142),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_6),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_197),
.A2(n_219),
.B(n_190),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_218),
.B(n_179),
.Y(n_224)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_202),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_209),
.C(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_206),
.Y(n_221)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_183),
.B1(n_178),
.B2(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_216),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_172),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_220),
.B1(n_194),
.B2(n_186),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_153),
.C(n_156),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_214),
.C(n_215),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_152),
.C(n_143),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_144),
.C(n_162),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_175),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_144),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_176),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_231),
.B1(n_233),
.B2(n_12),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_203),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_170),
.B(n_174),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_228),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_220),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_199),
.Y(n_230)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_170),
.B1(n_192),
.B2(n_171),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_188),
.B1(n_208),
.B2(n_13),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_171),
.B1(n_181),
.B2(n_191),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_191),
.C(n_169),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_204),
.C(n_197),
.Y(n_247)
);

AO21x1_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_184),
.B(n_173),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_236),
.A2(n_237),
.B(n_212),
.Y(n_248)
);

NOR4xp25_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_195),
.C(n_184),
.D(n_190),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_208),
.B(n_218),
.C(n_199),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_211),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_255),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_249),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_198),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_223),
.C(n_226),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_11),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_233),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_16),
.C(n_13),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_236),
.C(n_221),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_267),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_240),
.C(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_263),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_231),
.C(n_224),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_237),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_251),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_228),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_269),
.B(n_261),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_245),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_271),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_243),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_256),
.A2(n_243),
.B1(n_232),
.B2(n_229),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_256),
.Y(n_281)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_254),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_274),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_278),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_280),
.B(n_276),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_260),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_246),
.B1(n_260),
.B2(n_252),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_249),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_287),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_248),
.B1(n_272),
.B2(n_225),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_288),
.B(n_289),
.Y(n_293)
);

NOR3xp33_ASAP7_75t_SL g292 ( 
.A(n_290),
.B(n_281),
.C(n_235),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_288),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_295),
.B(n_284),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_291),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_293),
.A3(n_239),
.B1(n_242),
.B2(n_235),
.C1(n_15),
.C2(n_16),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_239),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_14),
.Y(n_299)
);


endmodule