module real_jpeg_9566_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_213;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_1),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_1),
.A2(n_52),
.B(n_66),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_1),
.A2(n_64),
.B1(n_70),
.B2(n_139),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_1),
.B(n_73),
.Y(n_188)
);

A2O1A1O1Ixp25_ASAP7_75t_L g200 ( 
.A1(n_1),
.A2(n_36),
.B(n_40),
.C(n_201),
.D(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_1),
.B(n_36),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_1),
.B(n_59),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_1),
.A2(n_25),
.B(n_216),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g247 ( 
.A1(n_1),
.A2(n_54),
.B(n_55),
.C(n_149),
.D(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_1),
.B(n_54),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_2),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_4),
.A2(n_64),
.B1(n_70),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_4),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_4),
.A2(n_52),
.B1(n_54),
.B2(n_75),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_75),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_75),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_5),
.A2(n_143),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_5),
.B(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_5),
.A2(n_190),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_5),
.A2(n_191),
.B(n_232),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_10),
.A2(n_64),
.B1(n_70),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_10),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_10),
.A2(n_52),
.B1(n_54),
.B2(n_91),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_91),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_91),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_11),
.A2(n_38),
.B1(n_52),
.B2(n_54),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_38),
.Y(n_143)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_13),
.A2(n_27),
.B1(n_30),
.B2(n_46),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_13),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_14),
.A2(n_64),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_14),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_14),
.A2(n_52),
.B1(n_54),
.B2(n_71),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_71),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_71),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_15),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_15),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_16),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_16),
.A2(n_53),
.B1(n_64),
.B2(n_70),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_16),
.A2(n_27),
.B1(n_30),
.B2(n_53),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_99),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_20),
.B(n_99),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.C(n_82),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_21),
.A2(n_22),
.B1(n_76),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_23),
.B(n_50),
.C(n_61),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_24),
.B(n_34),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_25),
.A2(n_26),
.B(n_32),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_25),
.A2(n_26),
.B1(n_85),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_25),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_25),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_25),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_26),
.A2(n_223),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_26),
.B(n_139),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_27),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_27),
.A2(n_43),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_30),
.B(n_41),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_30),
.B(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_35),
.A2(n_39),
.B1(n_47),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_37),
.B1(n_56),
.B2(n_57),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_36),
.A2(n_248),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_37),
.B(n_57),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_39),
.A2(n_45),
.B1(n_47),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_39),
.A2(n_47),
.B1(n_213),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_39),
.A2(n_246),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_40),
.A2(n_44),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_40),
.B(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_47),
.A2(n_87),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_47),
.B(n_166),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_47),
.A2(n_164),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_47),
.B(n_139),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_61),
.B2(n_62),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_56),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_55),
.A2(n_59),
.B1(n_60),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_55),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_58),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_59),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_69),
.B(n_72),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_68),
.B1(n_69),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_67),
.C(n_68),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_64),
.A2(n_65),
.B(n_139),
.C(n_140),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_68),
.A2(n_90),
.B(n_119),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_72),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_76),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_78),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_79),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_80),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_82),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.C(n_92),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_84),
.B(n_86),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B(n_96),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_98),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_95),
.A2(n_146),
.B1(n_147),
.B2(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_95),
.A2(n_96),
.B(n_172),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_122),
.B2(n_123),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_111),
.B2(n_112),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_108),
.B(n_110),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_108),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_121),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_122),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_153),
.B(n_277),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_150),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_128),
.B(n_150),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.C(n_132),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_131),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_133),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_144),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_135),
.B1(n_144),
.B2(n_145),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_137),
.A2(n_138),
.B1(n_141),
.B2(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_141),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B(n_148),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_193),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_176),
.B(n_192),
.Y(n_155)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_156),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_173),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_173),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_161),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_161),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.C(n_170),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_163),
.B1(n_170),
.B2(n_171),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_177),
.B(n_179),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_184),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_180),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_182),
.A2(n_184),
.B1(n_185),
.B2(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_182),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_189),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_186),
.A2(n_187),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_188),
.B(n_189),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_275),
.C(n_276),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_269),
.B(n_274),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_258),
.B(n_268),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_240),
.B(n_257),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_219),
.B(n_239),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_199),
.B(n_207),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_200),
.A2(n_203),
.B1(n_204),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_214),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_212),
.C(n_214),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_215),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_227),
.B(n_238),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_225),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_233),
.B(n_237),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_241),
.B(n_242),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_251),
.B2(n_256),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_250),
.C(n_256),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_255),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_259),
.B(n_260),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_265),
.C(n_266),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_262),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);


endmodule