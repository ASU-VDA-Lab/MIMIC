module fake_ariane_1595_n_1646 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1646);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1646;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_143;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_144;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_145;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_142;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_141;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_133),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_3),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_62),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_51),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_52),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_37),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_60),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_125),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_42),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_32),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_46),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_24),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_138),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_103),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_91),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_66),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_37),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_26),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_32),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_3),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_6),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_65),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_9),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_49),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_5),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_0),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_105),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_132),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_12),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_131),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_92),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_40),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_53),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_95),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_13),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_7),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_28),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_124),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_70),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_48),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_8),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_34),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_122),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_86),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_63),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_10),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_42),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_104),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_109),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_58),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_6),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_10),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_59),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_45),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_29),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_83),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_117),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_33),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_99),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_67),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_38),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_80),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_7),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_85),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_57),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_134),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_8),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_11),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_50),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_39),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_38),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_23),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_19),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_118),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_26),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_44),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_123),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_89),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_23),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_14),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_9),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_77),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_54),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_61),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_126),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_101),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_98),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_16),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_40),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_112),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_22),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_19),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_97),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_29),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_13),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_31),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_68),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_31),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_18),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_120),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_41),
.Y(n_257)
);

BUFx8_ASAP7_75t_SL g258 ( 
.A(n_79),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_39),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_28),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_4),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_55),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_81),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_69),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_72),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_128),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_18),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_47),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_74),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_64),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_1),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_114),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_33),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_4),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_14),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_0),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_30),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_15),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_191),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_251),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_258),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_195),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_251),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_236),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_261),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_177),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_261),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_142),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_142),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_216),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_216),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_152),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_177),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_163),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_145),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_145),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_182),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_164),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_165),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_200),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_182),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_237),
.Y(n_311)
);

INVx4_ASAP7_75t_R g312 ( 
.A(n_224),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_200),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_147),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_154),
.Y(n_315)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_161),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_167),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_160),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_207),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_197),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_213),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_218),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_170),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_222),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_151),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_237),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_242),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_242),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_225),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_227),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_172),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_235),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_247),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_207),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_175),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_183),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_161),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_201),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_184),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_253),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_190),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_257),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_260),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_276),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_158),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_168),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_171),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_179),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_180),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_196),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_203),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_206),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_284),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_256),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_282),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_282),
.Y(n_358)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_350),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_287),
.A2(n_151),
.B1(n_178),
.B2(n_185),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_283),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_284),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_208),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_283),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_281),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_292),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_280),
.B(n_211),
.Y(n_367)
);

NOR2x1_ASAP7_75t_L g368 ( 
.A(n_304),
.B(n_155),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_292),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_290),
.Y(n_370)
);

OR2x6_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_224),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

AND2x2_ASAP7_75t_SL g373 ( 
.A(n_279),
.B(n_212),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_293),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_294),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_215),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_316),
.B(n_264),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_294),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_304),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_325),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_348),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_288),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_306),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_347),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_286),
.B(n_232),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_306),
.Y(n_389)
);

BUFx10_ASAP7_75t_L g390 ( 
.A(n_300),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_310),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_310),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_301),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_309),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_348),
.B(n_239),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_321),
.B(n_349),
.Y(n_398)
);

AND3x2_ASAP7_75t_L g399 ( 
.A(n_287),
.B(n_248),
.C(n_241),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_313),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_319),
.A2(n_185),
.B1(n_255),
.B2(n_244),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_334),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_289),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_351),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_291),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_295),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_295),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_338),
.A2(n_178),
.B1(n_210),
.B2(n_244),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_296),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_296),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_297),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_303),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_297),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_352),
.B(n_271),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_361),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_361),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_373),
.B(n_307),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_366),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_373),
.B(n_308),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_373),
.B(n_363),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_363),
.B(n_317),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_420),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_382),
.B(n_352),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_354),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_353),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_374),
.Y(n_436)
);

AND3x2_ASAP7_75t_L g437 ( 
.A(n_377),
.B(n_330),
.C(n_329),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_366),
.Y(n_438)
);

CKINVDCx6p67_ASAP7_75t_R g439 ( 
.A(n_390),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_411),
.B(n_353),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_370),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_382),
.B(n_330),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_364),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_R g445 ( 
.A(n_365),
.B(n_323),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_364),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_369),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_374),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_386),
.Y(n_449)
);

AOI21x1_ASAP7_75t_L g450 ( 
.A1(n_369),
.A2(n_265),
.B(n_252),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_374),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

OAI22xp33_ASAP7_75t_L g453 ( 
.A1(n_377),
.A2(n_210),
.B1(n_255),
.B2(n_339),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_413),
.B(n_398),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_398),
.B(n_285),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_360),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_407),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_378),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_354),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_378),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_382),
.B(n_339),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_382),
.B(n_331),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_356),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_363),
.B(n_336),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_423),
.B(n_332),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_357),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_423),
.B(n_337),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_371),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_357),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_356),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_356),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_387),
.B(n_340),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_374),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_375),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_407),
.B(n_332),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_355),
.B(n_333),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_358),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_363),
.B(n_342),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_371),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_358),
.Y(n_485)
);

OAI22xp33_ASAP7_75t_L g486 ( 
.A1(n_416),
.A2(n_264),
.B1(n_162),
.B2(n_275),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_386),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_375),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_375),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_375),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_375),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_355),
.A2(n_318),
.B1(n_315),
.B2(n_320),
.Y(n_493)
);

AOI21x1_ASAP7_75t_L g494 ( 
.A1(n_367),
.A2(n_388),
.B(n_385),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_375),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_416),
.B(n_162),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_356),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_386),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_386),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_386),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_404),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_404),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_404),
.Y(n_504)
);

BUFx8_ASAP7_75t_SL g505 ( 
.A(n_401),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_422),
.B(n_156),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_404),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_387),
.B(n_333),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_404),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_408),
.Y(n_510)
);

AND2x6_ASAP7_75t_L g511 ( 
.A(n_368),
.B(n_376),
.Y(n_511)
);

BUFx6f_ASAP7_75t_SL g512 ( 
.A(n_390),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_371),
.B(n_335),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_387),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_422),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_380),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_376),
.B(n_397),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_408),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_408),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_379),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_L g524 ( 
.A(n_384),
.B(n_156),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_379),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_371),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_SL g528 ( 
.A1(n_371),
.A2(n_360),
.B1(n_385),
.B2(n_400),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_415),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_415),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_376),
.B(n_335),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_412),
.B(n_322),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_379),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_412),
.B(n_341),
.Y(n_534)
);

BUFx6f_ASAP7_75t_SL g535 ( 
.A(n_390),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_383),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_383),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_412),
.B(n_341),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_383),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_415),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_380),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_395),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_394),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_394),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_405),
.B(n_324),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g547 ( 
.A(n_359),
.B(n_278),
.C(n_275),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_368),
.B(n_343),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_362),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_394),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_362),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_409),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_409),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_409),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_393),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_393),
.Y(n_556)
);

NOR2x1p5_ASAP7_75t_L g557 ( 
.A(n_390),
.B(n_278),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_376),
.A2(n_271),
.B1(n_233),
.B2(n_272),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_393),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_396),
.Y(n_560)
);

NAND2x1_ASAP7_75t_L g561 ( 
.A(n_397),
.B(n_312),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_393),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_406),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_397),
.B(n_157),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_406),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_406),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_362),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_362),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_406),
.Y(n_569)
);

AND3x1_ASAP7_75t_L g570 ( 
.A(n_410),
.B(n_345),
.C(n_344),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_415),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_516),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_472),
.B(n_430),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_513),
.B(n_397),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_513),
.B(n_359),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_516),
.Y(n_576)
);

BUFx6f_ASAP7_75t_SL g577 ( 
.A(n_505),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_427),
.B(n_367),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_516),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_429),
.B(n_388),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_517),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_471),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_541),
.B(n_403),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_467),
.B(n_359),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_473),
.B(n_359),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_432),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_471),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_513),
.B(n_157),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_513),
.B(n_381),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_477),
.B(n_410),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_518),
.B(n_381),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_481),
.B(n_381),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_518),
.B(n_381),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_546),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_560),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_445),
.Y(n_596)
);

INVx8_ASAP7_75t_L g597 ( 
.A(n_512),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_434),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_458),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_434),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_532),
.B(n_410),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_433),
.B(n_410),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_474),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_474),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_441),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_434),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_463),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_465),
.B(n_389),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_473),
.B(n_159),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_484),
.B(n_159),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_482),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_482),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_433),
.B(n_389),
.Y(n_613)
);

O2A1O1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_508),
.A2(n_538),
.B(n_534),
.C(n_454),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_484),
.B(n_198),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_497),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_497),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_547),
.B(n_391),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_497),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_527),
.B(n_415),
.Y(n_620)
);

AND2x6_ASAP7_75t_SL g621 ( 
.A(n_543),
.B(n_343),
.Y(n_621)
);

AOI22x1_ASAP7_75t_L g622 ( 
.A1(n_555),
.A2(n_391),
.B1(n_392),
.B2(n_400),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_549),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_485),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_481),
.B(n_344),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_511),
.B(n_392),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_511),
.B(n_417),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_449),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_511),
.B(n_417),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_437),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_527),
.A2(n_249),
.B1(n_205),
.B2(n_209),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_549),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_470),
.B(n_345),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_560),
.B(n_402),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_485),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_453),
.B(n_402),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_465),
.B(n_417),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_470),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_465),
.B(n_417),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_L g640 ( 
.A(n_557),
.B(n_204),
.Y(n_640)
);

INVxp33_ASAP7_75t_L g641 ( 
.A(n_496),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_511),
.B(n_480),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_425),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_511),
.B(n_417),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_456),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_511),
.B(n_418),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_465),
.B(n_418),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_515),
.B(n_418),
.Y(n_648)
);

O2A1O1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_442),
.A2(n_414),
.B(n_419),
.C(n_298),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_549),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_511),
.B(n_480),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_570),
.B(n_418),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_449),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_531),
.B(n_418),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_551),
.Y(n_655)
);

INVx8_ASAP7_75t_L g656 ( 
.A(n_512),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_442),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_548),
.B(n_421),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_562),
.B(n_421),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_515),
.B(n_421),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_466),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_431),
.B(n_228),
.C(n_259),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_426),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_562),
.B(n_421),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_562),
.B(n_421),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_506),
.A2(n_269),
.B1(n_214),
.B2(n_270),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_426),
.Y(n_667)
);

BUFx8_ASAP7_75t_L g668 ( 
.A(n_512),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_428),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_563),
.B(n_421),
.Y(n_670)
);

BUFx8_ASAP7_75t_L g671 ( 
.A(n_512),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_555),
.A2(n_419),
.B(n_414),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_515),
.B(n_399),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_428),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_438),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_561),
.Y(n_676)
);

NOR2xp67_ASAP7_75t_L g677 ( 
.A(n_469),
.B(n_419),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_493),
.B(n_439),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_458),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_535),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_483),
.B(n_223),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_563),
.B(n_226),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_569),
.B(n_230),
.Y(n_683)
);

OR2x6_ASAP7_75t_L g684 ( 
.A(n_561),
.B(n_298),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_515),
.B(n_231),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_569),
.B(n_243),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_449),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_556),
.A2(n_169),
.B(n_268),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_557),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_569),
.B(n_246),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_556),
.B(n_559),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_565),
.B(n_254),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_458),
.B(n_267),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_565),
.B(n_566),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_524),
.A2(n_150),
.B1(n_149),
.B2(n_148),
.Y(n_695)
);

INVxp67_ASAP7_75t_SL g696 ( 
.A(n_461),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_447),
.Y(n_697)
);

AOI21x1_ASAP7_75t_L g698 ( 
.A1(n_450),
.A2(n_302),
.B(n_299),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_528),
.A2(n_233),
.B1(n_272),
.B2(n_271),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_462),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_461),
.B(n_273),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_542),
.B(n_202),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_462),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_464),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_461),
.B(n_274),
.Y(n_705)
);

O2A1O1Ixp5_ASAP7_75t_L g706 ( 
.A1(n_450),
.A2(n_302),
.B(n_299),
.C(n_202),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_464),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_564),
.B(n_1),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_435),
.B(n_141),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_440),
.B(n_143),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_542),
.B(n_233),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_496),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_542),
.B(n_144),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_542),
.B(n_202),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_533),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_468),
.B(n_475),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_535),
.A2(n_146),
.B1(n_266),
.B2(n_263),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_494),
.B(n_272),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_551),
.Y(n_719)
);

NAND2x1p5_ASAP7_75t_L g720 ( 
.A(n_498),
.B(n_212),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_551),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_449),
.B(n_202),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_468),
.B(n_153),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_494),
.B(n_2),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_535),
.B(n_5),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_533),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_449),
.B(n_202),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_567),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_475),
.B(n_166),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_539),
.Y(n_730)
);

AND2x6_ASAP7_75t_L g731 ( 
.A(n_539),
.B(n_212),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_581),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_583),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_643),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_594),
.B(n_457),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_599),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_702),
.A2(n_476),
.B(n_498),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_597),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_663),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_573),
.B(n_545),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_586),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_605),
.B(n_486),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_594),
.B(n_528),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_636),
.A2(n_558),
.B1(n_523),
.B2(n_526),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_597),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_SL g746 ( 
.A(n_596),
.B(n_174),
.C(n_173),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_599),
.Y(n_747)
);

NAND2x1p5_ASAP7_75t_L g748 ( 
.A(n_575),
.B(n_498),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_628),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_634),
.B(n_597),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_598),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_667),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_628),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_625),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_600),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_633),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_696),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_573),
.B(n_449),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_577),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_606),
.Y(n_760)
);

NOR2x2_ASAP7_75t_L g761 ( 
.A(n_634),
.B(n_535),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_657),
.B(n_476),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_669),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_628),
.Y(n_764)
);

AND2x4_ASAP7_75t_SL g765 ( 
.A(n_634),
.B(n_498),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_592),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_628),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_595),
.B(n_545),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_638),
.B(n_500),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_674),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_675),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_578),
.B(n_550),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_578),
.B(n_550),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_616),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_617),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_L g776 ( 
.A(n_653),
.B(n_540),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_699),
.A2(n_536),
.B1(n_523),
.B2(n_526),
.Y(n_777)
);

AND3x1_ASAP7_75t_L g778 ( 
.A(n_662),
.B(n_500),
.C(n_525),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_678),
.B(n_500),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_580),
.B(n_552),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_697),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_653),
.Y(n_782)
);

INVx5_ASAP7_75t_L g783 ( 
.A(n_656),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_580),
.B(n_552),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_653),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_700),
.A2(n_553),
.B1(n_554),
.B2(n_529),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_621),
.Y(n_787)
);

NOR2x1p5_ASAP7_75t_L g788 ( 
.A(n_680),
.B(n_708),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_685),
.A2(n_708),
.B1(n_651),
.B2(n_642),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_630),
.B(n_689),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_673),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_619),
.Y(n_792)
);

BUFx10_ASAP7_75t_L g793 ( 
.A(n_577),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_703),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_613),
.A2(n_554),
.B(n_553),
.C(n_544),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_704),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_645),
.B(n_500),
.Y(n_797)
);

AND2x6_ASAP7_75t_SL g798 ( 
.A(n_725),
.B(n_487),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_707),
.B(n_536),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_645),
.B(n_537),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_582),
.B(n_587),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_574),
.B(n_540),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_656),
.B(n_537),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_661),
.B(n_540),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_589),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_603),
.B(n_544),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_604),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_656),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_611),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_612),
.B(n_444),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_687),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_685),
.A2(n_525),
.B1(n_529),
.B2(n_530),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_624),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_666),
.B(n_540),
.Y(n_814)
);

AND3x1_ASAP7_75t_L g815 ( 
.A(n_662),
.B(n_529),
.C(n_530),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_635),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_588),
.B(n_529),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_602),
.B(n_444),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_668),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_687),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_SL g821 ( 
.A1(n_641),
.A2(n_217),
.B1(n_176),
.B2(n_181),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_584),
.A2(n_615),
.B1(n_673),
.B2(n_696),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_715),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_726),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_681),
.B(n_530),
.Y(n_825)
);

NOR2xp67_ASAP7_75t_L g826 ( 
.A(n_717),
.B(n_530),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_631),
.B(n_609),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_730),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_671),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_725),
.B(n_540),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_687),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_590),
.B(n_446),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_687),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_607),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_584),
.B(n_540),
.Y(n_835)
);

AND2x6_ASAP7_75t_L g836 ( 
.A(n_724),
.B(n_499),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_684),
.B(n_499),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_679),
.B(n_424),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_591),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_572),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_593),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_671),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_SL g843 ( 
.A1(n_608),
.A2(n_519),
.B(n_487),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_679),
.B(n_424),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_654),
.Y(n_845)
);

AND2x6_ASAP7_75t_L g846 ( 
.A(n_724),
.B(n_499),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_626),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_590),
.B(n_446),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_614),
.B(n_452),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_608),
.B(n_452),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_716),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_601),
.B(n_455),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_712),
.B(n_455),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_709),
.B(n_424),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_682),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_623),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_632),
.Y(n_857)
);

INVx5_ASAP7_75t_L g858 ( 
.A(n_684),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_610),
.B(n_424),
.Y(n_859)
);

NOR2x1p5_ASAP7_75t_L g860 ( 
.A(n_683),
.B(n_436),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_686),
.B(n_436),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_684),
.B(n_501),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_690),
.B(n_711),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_712),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_650),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_699),
.B(n_459),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_655),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_693),
.B(n_436),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_647),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_719),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_676),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_710),
.B(n_436),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_691),
.B(n_459),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_627),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_576),
.B(n_443),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_579),
.B(n_443),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_728),
.Y(n_877)
);

BUFx6f_ASAP7_75t_SL g878 ( 
.A(n_731),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_695),
.B(n_443),
.Y(n_879)
);

AND2x6_ASAP7_75t_L g880 ( 
.A(n_629),
.B(n_501),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_677),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_701),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_694),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_658),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_718),
.B(n_460),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_647),
.B(n_501),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_640),
.B(n_567),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_SL g888 ( 
.A(n_649),
.B(n_713),
.C(n_692),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_644),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_721),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_659),
.Y(n_891)
);

CKINVDCx16_ASAP7_75t_R g892 ( 
.A(n_731),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_622),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_664),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_648),
.B(n_522),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_705),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_585),
.B(n_443),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_585),
.B(n_448),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_648),
.B(n_522),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_672),
.B(n_618),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_620),
.A2(n_519),
.B1(n_488),
.B2(n_509),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_646),
.B(n_448),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_665),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_652),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_670),
.B(n_522),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_723),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_750),
.B(n_637),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_735),
.B(n_637),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_754),
.B(n_639),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_850),
.A2(n_714),
.B(n_702),
.Y(n_910)
);

NOR2xp67_ASAP7_75t_SL g911 ( 
.A(n_741),
.B(n_639),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_801),
.A2(n_660),
.B1(n_729),
.B2(n_714),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_756),
.B(n_660),
.Y(n_913)
);

OAI22x1_ASAP7_75t_L g914 ( 
.A1(n_788),
.A2(n_727),
.B1(n_722),
.B2(n_698),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_783),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_883),
.B(n_488),
.Y(n_916)
);

BUFx12f_ASAP7_75t_L g917 ( 
.A(n_793),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_819),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_734),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_801),
.A2(n_509),
.B1(n_504),
.B2(n_507),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_733),
.B(n_568),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_822),
.B(n_789),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_843),
.A2(n_706),
.B(n_740),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_791),
.B(n_688),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_850),
.A2(n_727),
.B(n_722),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_783),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_751),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_783),
.Y(n_928)
);

AND2x6_ASAP7_75t_L g929 ( 
.A(n_837),
.B(n_571),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_863),
.A2(n_507),
.B(n_510),
.C(n_521),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_772),
.A2(n_510),
.B1(n_514),
.B2(n_521),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_772),
.A2(n_720),
.B1(n_448),
.B2(n_451),
.Y(n_932)
);

O2A1O1Ixp5_ASAP7_75t_L g933 ( 
.A1(n_835),
.A2(n_571),
.B(n_502),
.C(n_520),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_733),
.B(n_451),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_739),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_752),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_763),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_770),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_855),
.B(n_451),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_864),
.B(n_742),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_853),
.B(n_768),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_783),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_759),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_750),
.B(n_502),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_906),
.A2(n_503),
.B(n_479),
.C(n_478),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_832),
.A2(n_503),
.B(n_492),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_SL g947 ( 
.A1(n_882),
.A2(n_821),
.B1(n_787),
.B2(n_750),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_755),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_779),
.B(n_478),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_779),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_858),
.B(n_490),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_858),
.B(n_490),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_839),
.B(n_479),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_766),
.B(n_489),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_760),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_773),
.B(n_491),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_841),
.B(n_491),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_774),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_732),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_832),
.A2(n_495),
.B(n_492),
.Y(n_960)
);

BUFx2_ASAP7_75t_SL g961 ( 
.A(n_793),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_805),
.B(n_491),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_764),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_771),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_845),
.B(n_495),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_888),
.A2(n_495),
.B(n_720),
.C(n_16),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_848),
.A2(n_490),
.B(n_221),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_738),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_858),
.B(n_490),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_829),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_848),
.A2(n_869),
.B(n_780),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_790),
.B(n_12),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_773),
.A2(n_490),
.B1(n_188),
.B2(n_187),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_780),
.B(n_490),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_890),
.B(n_186),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_790),
.B(n_15),
.Y(n_976)
);

O2A1O1Ixp5_ASAP7_75t_L g977 ( 
.A1(n_879),
.A2(n_731),
.B(n_20),
.C(n_21),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_764),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_784),
.A2(n_740),
.B1(n_796),
.B2(n_781),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_R g980 ( 
.A(n_842),
.B(n_731),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_837),
.Y(n_981)
);

AOI21x1_ASAP7_75t_L g982 ( 
.A1(n_885),
.A2(n_849),
.B(n_893),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_784),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_888),
.A2(n_17),
.B(n_20),
.C(n_21),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_852),
.A2(n_229),
.B(n_262),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_904),
.B(n_194),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_778),
.B(n_220),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_797),
.A2(n_219),
.B(n_245),
.C(n_199),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_794),
.B(n_731),
.Y(n_989)
);

OA22x2_ASAP7_75t_L g990 ( 
.A1(n_765),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_849),
.A2(n_240),
.B(n_238),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_823),
.A2(n_27),
.B(n_30),
.C(n_34),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_795),
.A2(n_240),
.B(n_238),
.C(n_212),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_775),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_792),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_745),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_762),
.B(n_36),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_745),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_886),
.A2(n_899),
.B(n_895),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_896),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_851),
.B(n_884),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_815),
.B(n_202),
.Y(n_1002)
);

AOI21x1_ASAP7_75t_L g1003 ( 
.A1(n_885),
.A2(n_240),
.B(n_238),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_769),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_807),
.B(n_36),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_862),
.B(n_800),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_SL g1007 ( 
.A(n_746),
.B(n_41),
.C(n_43),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_809),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_813),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_862),
.B(n_240),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_764),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_SL g1012 ( 
.A1(n_861),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_870),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_762),
.Y(n_1014)
);

AOI33xp33_ASAP7_75t_L g1015 ( 
.A1(n_816),
.A2(n_238),
.A3(n_212),
.B1(n_56),
.B2(n_71),
.B3(n_75),
.Y(n_1015)
);

AOI21x1_ASAP7_75t_L g1016 ( 
.A1(n_758),
.A2(n_76),
.B(n_78),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_834),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_798),
.B(n_82),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_824),
.A2(n_87),
.B(n_88),
.C(n_90),
.Y(n_1019)
);

BUFx2_ASAP7_75t_SL g1020 ( 
.A(n_808),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_776),
.A2(n_93),
.B(n_94),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_757),
.A2(n_96),
.B(n_102),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_803),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_795),
.A2(n_110),
.B(n_115),
.C(n_116),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_782),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_SL g1026 ( 
.A1(n_744),
.A2(n_121),
.B1(n_135),
.B2(n_136),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_828),
.Y(n_1027)
);

INVx6_ASAP7_75t_L g1028 ( 
.A(n_803),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_769),
.B(n_140),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_786),
.A2(n_872),
.B(n_854),
.C(n_844),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_873),
.A2(n_899),
.B(n_895),
.Y(n_1031)
);

INVx3_ASAP7_75t_SL g1032 ( 
.A(n_761),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_803),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_873),
.A2(n_886),
.B(n_818),
.Y(n_1034)
);

NOR4xp25_ASAP7_75t_L g1035 ( 
.A(n_984),
.B(n_830),
.C(n_866),
.D(n_786),
.Y(n_1035)
);

AOI221x1_ASAP7_75t_L g1036 ( 
.A1(n_1026),
.A2(n_900),
.B1(n_737),
.B2(n_817),
.C(n_859),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_979),
.B(n_820),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_1031),
.A2(n_818),
.B(n_905),
.Y(n_1038)
);

AO31x2_ASAP7_75t_L g1039 ( 
.A1(n_1034),
.A2(n_903),
.A3(n_891),
.B(n_894),
.Y(n_1039)
);

AO21x1_ASAP7_75t_L g1040 ( 
.A1(n_922),
.A2(n_814),
.B(n_804),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_971),
.A2(n_810),
.B(n_806),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_1003),
.A2(n_799),
.B(n_810),
.Y(n_1042)
);

OA21x2_ASAP7_75t_L g1043 ( 
.A1(n_923),
.A2(n_806),
.B(n_799),
.Y(n_1043)
);

INVx3_ASAP7_75t_SL g1044 ( 
.A(n_943),
.Y(n_1044)
);

AO31x2_ASAP7_75t_L g1045 ( 
.A1(n_979),
.A2(n_902),
.A3(n_898),
.B(n_897),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_982),
.A2(n_802),
.B(n_875),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_918),
.Y(n_1047)
);

INVxp67_ASAP7_75t_SL g1048 ( 
.A(n_1006),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_919),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_941),
.B(n_847),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_999),
.A2(n_836),
.B(n_846),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_L g1052 ( 
.A(n_908),
.B(n_782),
.Y(n_1052)
);

NAND3xp33_ASAP7_75t_L g1053 ( 
.A(n_983),
.B(n_825),
.C(n_868),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_960),
.A2(n_875),
.B(n_831),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_917),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1017),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_966),
.A2(n_826),
.B(n_887),
.C(n_860),
.Y(n_1057)
);

AOI221xp5_ASAP7_75t_SL g1058 ( 
.A1(n_992),
.A2(n_838),
.B1(n_876),
.B2(n_777),
.C(n_840),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_999),
.A2(n_923),
.B(n_912),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_940),
.B(n_871),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_SL g1061 ( 
.A(n_1018),
.B(n_881),
.C(n_748),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_970),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_983),
.A2(n_840),
.B1(n_748),
.B2(n_812),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_921),
.B(n_877),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_946),
.A2(n_925),
.B(n_933),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_L g1066 ( 
.A(n_1001),
.B(n_749),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_1015),
.A2(n_901),
.B(n_874),
.C(n_736),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_981),
.B(n_871),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_910),
.A2(n_836),
.B(n_846),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_959),
.Y(n_1070)
);

AOI221xp5_ASAP7_75t_SL g1071 ( 
.A1(n_912),
.A2(n_736),
.B1(n_747),
.B2(n_867),
.C(n_865),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_1032),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1001),
.B(n_874),
.Y(n_1073)
);

AOI221x1_ASAP7_75t_L g1074 ( 
.A1(n_1024),
.A2(n_856),
.B1(n_857),
.B2(n_889),
.C(n_767),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_956),
.A2(n_820),
.B(n_785),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1016),
.A2(n_833),
.B(n_749),
.Y(n_1076)
);

AO32x2_ASAP7_75t_L g1077 ( 
.A1(n_931),
.A2(n_846),
.A3(n_836),
.B1(n_880),
.B2(n_889),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_SL g1078 ( 
.A(n_929),
.B(n_892),
.Y(n_1078)
);

NAND3x1_ASAP7_75t_L g1079 ( 
.A(n_972),
.B(n_747),
.C(n_753),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_950),
.B(n_782),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_907),
.Y(n_1081)
);

AO22x2_ASAP7_75t_L g1082 ( 
.A1(n_950),
.A2(n_846),
.B1(n_836),
.B2(n_811),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_915),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1014),
.B(n_889),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_986),
.A2(n_811),
.B(n_785),
.C(n_880),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_935),
.B(n_880),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_915),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_932),
.A2(n_880),
.B(n_878),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_936),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_932),
.A2(n_878),
.B(n_974),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_937),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_938),
.B(n_964),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_993),
.A2(n_920),
.B(n_945),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_907),
.B(n_944),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_L g1095 ( 
.A(n_915),
.B(n_926),
.Y(n_1095)
);

INVx3_ASAP7_75t_SL g1096 ( 
.A(n_976),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_1000),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1012),
.A2(n_924),
.B(n_1007),
.C(n_930),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1002),
.A2(n_1021),
.B(n_967),
.Y(n_1099)
);

AOI21x1_ASAP7_75t_SL g1100 ( 
.A1(n_1005),
.A2(n_909),
.B(n_913),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_920),
.A2(n_977),
.B(n_953),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1027),
.B(n_1004),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_926),
.B(n_928),
.Y(n_1104)
);

AO32x2_ASAP7_75t_L g1105 ( 
.A1(n_973),
.A2(n_947),
.A3(n_990),
.B1(n_996),
.B2(n_914),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1022),
.A2(n_953),
.B(n_965),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_997),
.B(n_939),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1029),
.A2(n_916),
.B(n_1019),
.Y(n_1108)
);

BUFx4f_ASAP7_75t_L g1109 ( 
.A(n_926),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_957),
.B(n_911),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1023),
.A2(n_1033),
.B(n_989),
.Y(n_1111)
);

CKINVDCx11_ASAP7_75t_R g1112 ( 
.A(n_963),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_985),
.A2(n_987),
.B(n_1010),
.Y(n_1113)
);

AOI21xp33_ASAP7_75t_L g1114 ( 
.A1(n_962),
.A2(n_954),
.B(n_988),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_928),
.B(n_942),
.Y(n_1115)
);

INVxp67_ASAP7_75t_SL g1116 ( 
.A(n_949),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_927),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_990),
.A2(n_996),
.B1(n_1020),
.B2(n_968),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_951),
.A2(n_952),
.B(n_969),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_975),
.B(n_934),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_929),
.A2(n_1028),
.B1(n_1033),
.B2(n_961),
.Y(n_1121)
);

AOI221x1_ASAP7_75t_L g1122 ( 
.A1(n_948),
.A2(n_1013),
.B1(n_995),
.B2(n_994),
.C(n_955),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1028),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_958),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_968),
.A2(n_998),
.B(n_929),
.Y(n_1125)
);

AO32x2_ASAP7_75t_L g1126 ( 
.A1(n_929),
.A2(n_1025),
.A3(n_963),
.B1(n_978),
.B2(n_1011),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_963),
.B(n_978),
.Y(n_1127)
);

BUFx4_ASAP7_75t_SL g1128 ( 
.A(n_980),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_1025),
.A2(n_991),
.B(n_923),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_942),
.A2(n_991),
.B(n_1003),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_942),
.A2(n_724),
.B(n_971),
.Y(n_1131)
);

OAI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_979),
.A2(n_377),
.B(n_594),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_941),
.B(n_735),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_941),
.B(n_735),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_SL g1135 ( 
.A1(n_979),
.A2(n_1030),
.B(n_999),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_941),
.B(n_735),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_991),
.A2(n_1003),
.B(n_982),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_1031),
.A2(n_1034),
.A3(n_991),
.B(n_979),
.Y(n_1138)
);

NAND2x1_ASAP7_75t_L g1139 ( 
.A(n_963),
.B(n_749),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_922),
.A2(n_827),
.B(n_573),
.C(n_735),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_940),
.B(n_432),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_940),
.B(n_432),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_940),
.B(n_432),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_979),
.B(n_822),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_941),
.B(n_735),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_950),
.B(n_738),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_991),
.A2(n_1003),
.B(n_982),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_915),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_919),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1031),
.A2(n_971),
.B(n_1034),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_991),
.A2(n_1003),
.B(n_982),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_991),
.A2(n_1003),
.B(n_982),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1031),
.A2(n_1034),
.A3(n_991),
.B(n_979),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_991),
.A2(n_1003),
.B(n_982),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_979),
.A2(n_594),
.B(n_735),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_979),
.A2(n_594),
.B1(n_735),
.B2(n_595),
.Y(n_1156)
);

NOR2xp67_ASAP7_75t_L g1157 ( 
.A(n_979),
.B(n_783),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_922),
.A2(n_827),
.B(n_573),
.C(n_735),
.Y(n_1158)
);

OA21x2_ASAP7_75t_L g1159 ( 
.A1(n_991),
.A2(n_923),
.B(n_982),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1003),
.A2(n_982),
.B(n_991),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_941),
.B(n_733),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_941),
.B(n_733),
.Y(n_1162)
);

AOI211x1_ASAP7_75t_L g1163 ( 
.A1(n_908),
.A2(n_979),
.B(n_743),
.C(n_1005),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1031),
.A2(n_971),
.B(n_1034),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_941),
.B(n_735),
.Y(n_1165)
);

NAND2xp33_ASAP7_75t_L g1166 ( 
.A(n_979),
.B(n_432),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_941),
.B(n_735),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1073),
.B(n_1155),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1132),
.A2(n_1144),
.B1(n_1166),
.B2(n_1133),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1160),
.A2(n_1147),
.B(n_1137),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1132),
.B(n_1140),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1151),
.A2(n_1154),
.B(n_1152),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1130),
.A2(n_1065),
.B(n_1042),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1045),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1150),
.A2(n_1164),
.B(n_1099),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1055),
.Y(n_1176)
);

CKINVDCx6p67_ASAP7_75t_R g1177 ( 
.A(n_1044),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1158),
.A2(n_1059),
.B(n_1053),
.Y(n_1178)
);

BUFx12f_ASAP7_75t_L g1179 ( 
.A(n_1112),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1163),
.B(n_1135),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1163),
.B(n_1045),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1156),
.B(n_1141),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1094),
.B(n_1081),
.Y(n_1183)
);

NOR3xp33_ASAP7_75t_SL g1184 ( 
.A(n_1142),
.B(n_1143),
.C(n_1098),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1102),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1126),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1128),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1134),
.A2(n_1136),
.B(n_1165),
.C(n_1145),
.Y(n_1188)
);

BUFx2_ASAP7_75t_R g1189 ( 
.A(n_1062),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1053),
.A2(n_1101),
.B(n_1093),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1040),
.A2(n_1038),
.A3(n_1036),
.B(n_1041),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1049),
.Y(n_1192)
);

OAI222xp33_ASAP7_75t_L g1193 ( 
.A1(n_1161),
.A2(n_1162),
.B1(n_1050),
.B2(n_1116),
.C1(n_1121),
.C2(n_1167),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1045),
.B(n_1064),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1101),
.A2(n_1093),
.B(n_1131),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1054),
.A2(n_1106),
.B(n_1046),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_SL g1197 ( 
.A1(n_1110),
.A2(n_1125),
.B(n_1051),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1107),
.A2(n_1067),
.B(n_1037),
.C(n_1114),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1071),
.A2(n_1131),
.B(n_1069),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1069),
.A2(n_1111),
.B(n_1076),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1072),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_1082),
.B(n_1125),
.Y(n_1202)
);

NOR2x1_ASAP7_75t_R g1203 ( 
.A(n_1070),
.B(n_1047),
.Y(n_1203)
);

NAND2x1p5_ASAP7_75t_L g1204 ( 
.A(n_1109),
.B(n_1121),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_1097),
.Y(n_1205)
);

AOI222xp33_ASAP7_75t_SL g1206 ( 
.A1(n_1089),
.A2(n_1091),
.B1(n_1149),
.B2(n_1118),
.C1(n_1063),
.C2(n_1105),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1123),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1061),
.A2(n_1096),
.B1(n_1117),
.B2(n_1124),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1090),
.A2(n_1088),
.B(n_1100),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1103),
.B(n_1060),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1157),
.A2(n_1108),
.B1(n_1120),
.B2(n_1043),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_SL g1212 ( 
.A1(n_1119),
.A2(n_1075),
.B(n_1113),
.Y(n_1212)
);

OR2x6_ASAP7_75t_L g1213 ( 
.A(n_1079),
.B(n_1066),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1048),
.B(n_1084),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1086),
.B(n_1146),
.Y(n_1215)
);

AO21x1_ASAP7_75t_L g1216 ( 
.A1(n_1052),
.A2(n_1080),
.B(n_1068),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1058),
.A2(n_1057),
.B(n_1122),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_1109),
.B(n_1148),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1085),
.A2(n_1035),
.B1(n_1159),
.B2(n_1105),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1129),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1039),
.Y(n_1221)
);

AO21x2_ASAP7_75t_L g1222 ( 
.A1(n_1035),
.A2(n_1115),
.B(n_1104),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1078),
.A2(n_1105),
.B1(n_1058),
.B2(n_1087),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1083),
.A2(n_1127),
.B1(n_1139),
.B2(n_1077),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1039),
.Y(n_1225)
);

BUFx12f_ASAP7_75t_L g1226 ( 
.A(n_1083),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1138),
.A2(n_1153),
.B(n_1077),
.Y(n_1227)
);

AOI222xp33_ASAP7_75t_L g1228 ( 
.A1(n_1078),
.A2(n_1095),
.B1(n_1077),
.B2(n_1126),
.C1(n_1138),
.C2(n_1153),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1126),
.A2(n_1071),
.B(n_1137),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1132),
.A2(n_1158),
.B(n_1140),
.C(n_827),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1073),
.B(n_1155),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1074),
.A2(n_1040),
.A3(n_1164),
.B(n_1150),
.Y(n_1232)
);

NAND2x1p5_ASAP7_75t_L g1233 ( 
.A(n_1109),
.B(n_858),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1133),
.B(n_1167),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1160),
.A2(n_1147),
.B(n_1137),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1133),
.B(n_1167),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1092),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1132),
.A2(n_402),
.B1(n_636),
.B2(n_453),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1166),
.A2(n_377),
.B1(n_735),
.B2(n_636),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_SL g1240 ( 
.A1(n_1155),
.A2(n_1135),
.B(n_1059),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1160),
.A2(n_1147),
.B(n_1137),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1133),
.B(n_1167),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1132),
.B(n_377),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_1112),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1092),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1086),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1071),
.A2(n_1147),
.B(n_1137),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1056),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1092),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1064),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1166),
.A2(n_377),
.B1(n_735),
.B2(n_636),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1073),
.B(n_1155),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1160),
.A2(n_1147),
.B(n_1137),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1070),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1160),
.A2(n_1147),
.B(n_1137),
.Y(n_1255)
);

AO22x2_ASAP7_75t_L g1256 ( 
.A1(n_1163),
.A2(n_1144),
.B1(n_1135),
.B2(n_1059),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1140),
.A2(n_1158),
.B(n_1132),
.Y(n_1257)
);

CKINVDCx6p67_ASAP7_75t_R g1258 ( 
.A(n_1044),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1128),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1073),
.B(n_1155),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_SL g1261 ( 
.A1(n_1155),
.A2(n_1135),
.B(n_1059),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1140),
.A2(n_1158),
.B(n_1132),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1160),
.A2(n_1147),
.B(n_1137),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1166),
.A2(n_377),
.B1(n_735),
.B2(n_636),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1045),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1092),
.Y(n_1266)
);

OAI22x1_ASAP7_75t_L g1267 ( 
.A1(n_1121),
.A2(n_416),
.B1(n_360),
.B2(n_496),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1064),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1092),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1112),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1140),
.A2(n_1158),
.B(n_1132),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1112),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1112),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1070),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_SL g1275 ( 
.A1(n_1140),
.A2(n_1158),
.B(n_1144),
.C(n_1155),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1132),
.A2(n_402),
.B1(n_636),
.B2(n_453),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1160),
.A2(n_1147),
.B(n_1137),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1140),
.A2(n_1158),
.B(n_1132),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1132),
.B(n_377),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1160),
.A2(n_1147),
.B(n_1137),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1192),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1239),
.A2(n_1264),
.B1(n_1251),
.B2(n_1169),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1170),
.A2(n_1241),
.B(n_1235),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1169),
.A2(n_1182),
.B1(n_1230),
.B2(n_1238),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1184),
.B(n_1168),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1238),
.A2(n_1276),
.B1(n_1184),
.B2(n_1190),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1243),
.A2(n_1279),
.B(n_1198),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1276),
.A2(n_1190),
.B1(n_1243),
.B2(n_1279),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_SL g1289 ( 
.A1(n_1198),
.A2(n_1188),
.B(n_1257),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1275),
.A2(n_1178),
.B(n_1195),
.Y(n_1290)
);

BUFx12f_ASAP7_75t_L g1291 ( 
.A(n_1270),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1178),
.A2(n_1271),
.B1(n_1278),
.B2(n_1257),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1168),
.B(n_1231),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1262),
.A2(n_1271),
.B1(n_1278),
.B2(n_1231),
.Y(n_1294)
);

O2A1O1Ixp5_ASAP7_75t_L g1295 ( 
.A1(n_1262),
.A2(n_1171),
.B(n_1195),
.C(n_1219),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1226),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1252),
.A2(n_1260),
.B1(n_1256),
.B2(n_1171),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1240),
.A2(n_1261),
.B(n_1188),
.C(n_1180),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1268),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1253),
.A2(n_1255),
.B(n_1277),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1176),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1194),
.B(n_1234),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1206),
.A2(n_1267),
.B1(n_1208),
.B2(n_1215),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1236),
.B(n_1242),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1254),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1183),
.B(n_1274),
.Y(n_1306)
);

O2A1O1Ixp5_ASAP7_75t_L g1307 ( 
.A1(n_1219),
.A2(n_1211),
.B(n_1181),
.C(n_1224),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1260),
.B(n_1256),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1256),
.A2(n_1223),
.B1(n_1208),
.B2(n_1237),
.Y(n_1309)
);

AND2x4_ASAP7_75t_SL g1310 ( 
.A(n_1177),
.B(n_1258),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1223),
.A2(n_1245),
.B1(n_1185),
.B2(n_1249),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1173),
.A2(n_1172),
.B(n_1175),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1270),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1197),
.A2(n_1212),
.B(n_1246),
.C(n_1193),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1266),
.B(n_1269),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1246),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1189),
.A2(n_1244),
.B1(n_1202),
.B2(n_1199),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1207),
.Y(n_1318)
);

AOI221xp5_ASAP7_75t_L g1319 ( 
.A1(n_1174),
.A2(n_1265),
.B1(n_1193),
.B2(n_1206),
.C(n_1214),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1205),
.Y(n_1320)
);

CKINVDCx6p67_ASAP7_75t_R g1321 ( 
.A(n_1179),
.Y(n_1321)
);

AOI221xp5_ASAP7_75t_L g1322 ( 
.A1(n_1224),
.A2(n_1186),
.B1(n_1220),
.B2(n_1221),
.C(n_1225),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1272),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1209),
.A2(n_1196),
.B(n_1200),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1189),
.A2(n_1244),
.B1(n_1199),
.B2(n_1273),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1201),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1272),
.A2(n_1273),
.B1(n_1204),
.B2(n_1217),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1187),
.A2(n_1259),
.B(n_1222),
.C(n_1204),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1228),
.B(n_1227),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1203),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1217),
.A2(n_1213),
.B1(n_1227),
.B2(n_1233),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1233),
.A2(n_1218),
.B(n_1229),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1218),
.A2(n_1248),
.B1(n_1247),
.B2(n_1228),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1247),
.A2(n_1191),
.B1(n_1232),
.B2(n_1216),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1232),
.B(n_1191),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1191),
.B(n_1232),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1263),
.B(n_1280),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1239),
.A2(n_1264),
.B1(n_1251),
.B2(n_1158),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1230),
.A2(n_1132),
.B(n_1140),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1230),
.A2(n_1132),
.B(n_1140),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1234),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1210),
.B(n_1250),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1210),
.B(n_1250),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1250),
.B(n_1268),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1239),
.A2(n_1264),
.B1(n_1251),
.B2(n_1158),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1210),
.B(n_1250),
.Y(n_1346)
);

BUFx4_ASAP7_75t_R g1347 ( 
.A(n_1189),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1239),
.A2(n_1264),
.B1(n_1251),
.B2(n_1158),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1250),
.B(n_1268),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1192),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1230),
.A2(n_1132),
.B(n_1140),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1210),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1210),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1210),
.B(n_1250),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1230),
.A2(n_1132),
.B(n_1140),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1170),
.A2(n_1241),
.B(n_1235),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1170),
.A2(n_1241),
.B(n_1235),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1210),
.B(n_1250),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1281),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1335),
.B(n_1308),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1286),
.A2(n_1339),
.B(n_1355),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1307),
.A2(n_1295),
.B(n_1329),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1337),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1305),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1297),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1334),
.A2(n_1329),
.B(n_1297),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1293),
.B(n_1294),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1336),
.B(n_1302),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1333),
.A2(n_1288),
.B(n_1309),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1290),
.A2(n_1322),
.B(n_1333),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1350),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1352),
.B(n_1353),
.Y(n_1372)
);

AO21x2_ASAP7_75t_L g1373 ( 
.A1(n_1288),
.A2(n_1309),
.B(n_1287),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1316),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1293),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1324),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1292),
.A2(n_1311),
.B(n_1331),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1292),
.B(n_1324),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1294),
.B(n_1285),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1315),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1319),
.A2(n_1331),
.B(n_1311),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1283),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1312),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1283),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1286),
.A2(n_1284),
.B1(n_1282),
.B2(n_1348),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1342),
.B(n_1343),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1327),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1327),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1299),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1346),
.B(n_1358),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1317),
.A2(n_1340),
.B(n_1351),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1289),
.A2(n_1282),
.B(n_1303),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1300),
.B(n_1357),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1332),
.B(n_1328),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1357),
.B(n_1356),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1356),
.Y(n_1396)
);

NAND3xp33_ASAP7_75t_L g1397 ( 
.A(n_1284),
.B(n_1338),
.C(n_1348),
.Y(n_1397)
);

OR2x6_ASAP7_75t_L g1398 ( 
.A(n_1314),
.B(n_1345),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1326),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1338),
.A2(n_1345),
.B(n_1298),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1379),
.B(n_1397),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1359),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1378),
.B(n_1306),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1378),
.B(n_1304),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1378),
.B(n_1341),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1396),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1385),
.A2(n_1397),
.B1(n_1400),
.B2(n_1379),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1383),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1359),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1367),
.B(n_1375),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1391),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1372),
.B(n_1365),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1372),
.B(n_1344),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1382),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1384),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1363),
.B(n_1325),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1363),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1363),
.B(n_1325),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1364),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1367),
.B(n_1354),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1372),
.B(n_1349),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1382),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1375),
.B(n_1365),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1362),
.B(n_1366),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1366),
.B(n_1368),
.Y(n_1425)
);

OR2x6_ASAP7_75t_L g1426 ( 
.A(n_1411),
.B(n_1394),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1402),
.Y(n_1427)
);

NAND3xp33_ASAP7_75t_L g1428 ( 
.A(n_1401),
.B(n_1361),
.C(n_1385),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1401),
.A2(n_1392),
.B1(n_1361),
.B2(n_1373),
.Y(n_1429)
);

AOI21xp33_ASAP7_75t_L g1430 ( 
.A1(n_1424),
.A2(n_1366),
.B(n_1373),
.Y(n_1430)
);

NOR2xp67_ASAP7_75t_L g1431 ( 
.A(n_1417),
.B(n_1387),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1407),
.A2(n_1392),
.B1(n_1373),
.B2(n_1369),
.Y(n_1432)
);

AOI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1407),
.A2(n_1366),
.B1(n_1392),
.B2(n_1373),
.C(n_1377),
.Y(n_1433)
);

AOI221xp5_ASAP7_75t_L g1434 ( 
.A1(n_1425),
.A2(n_1392),
.B1(n_1373),
.B2(n_1377),
.C(n_1369),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1420),
.A2(n_1400),
.B1(n_1398),
.B2(n_1388),
.Y(n_1435)
);

AOI211x1_ASAP7_75t_L g1436 ( 
.A1(n_1420),
.A2(n_1390),
.B(n_1386),
.C(n_1374),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1404),
.B(n_1364),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1404),
.B(n_1386),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1411),
.A2(n_1398),
.B1(n_1388),
.B2(n_1381),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1412),
.B(n_1413),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1409),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1408),
.Y(n_1442)
);

AOI221xp5_ASAP7_75t_L g1443 ( 
.A1(n_1425),
.A2(n_1392),
.B1(n_1377),
.B2(n_1369),
.C(n_1360),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1419),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1415),
.A2(n_1395),
.B(n_1393),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1411),
.A2(n_1369),
.B1(n_1391),
.B2(n_1377),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1410),
.B(n_1362),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1411),
.A2(n_1398),
.B1(n_1388),
.B2(n_1381),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1409),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1423),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1423),
.B(n_1362),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1412),
.B(n_1374),
.Y(n_1452)
);

OAI221xp5_ASAP7_75t_L g1453 ( 
.A1(n_1425),
.A2(n_1381),
.B1(n_1370),
.B2(n_1362),
.C(n_1387),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_L g1454 ( 
.A(n_1414),
.B(n_1362),
.C(n_1370),
.Y(n_1454)
);

OAI221xp5_ASAP7_75t_L g1455 ( 
.A1(n_1416),
.A2(n_1381),
.B1(n_1370),
.B2(n_1387),
.C(n_1394),
.Y(n_1455)
);

AO21x1_ASAP7_75t_SL g1456 ( 
.A1(n_1412),
.A2(n_1376),
.B(n_1371),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1403),
.B(n_1360),
.Y(n_1457)
);

AOI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1416),
.A2(n_1360),
.B1(n_1391),
.B2(n_1380),
.C(n_1389),
.Y(n_1458)
);

OAI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1416),
.A2(n_1381),
.B1(n_1370),
.B2(n_1394),
.C(n_1398),
.Y(n_1459)
);

OA21x2_ASAP7_75t_L g1460 ( 
.A1(n_1434),
.A2(n_1393),
.B(n_1395),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1457),
.B(n_1404),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1427),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1441),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1445),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1449),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1440),
.Y(n_1466)
);

NAND3xp33_ASAP7_75t_SL g1467 ( 
.A(n_1433),
.B(n_1418),
.C(n_1399),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1457),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1431),
.B(n_1403),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1450),
.B(n_1405),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1452),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1452),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1447),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1436),
.B(n_1405),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1438),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1451),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1454),
.B(n_1413),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1442),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1428),
.B(n_1321),
.Y(n_1479)
);

NOR2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1444),
.B(n_1291),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1456),
.B(n_1437),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_L g1482 ( 
.A(n_1443),
.B(n_1398),
.C(n_1370),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1435),
.B(n_1413),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1430),
.A2(n_1393),
.B(n_1395),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1444),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1481),
.B(n_1437),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1466),
.B(n_1421),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1472),
.B(n_1432),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1460),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1481),
.B(n_1403),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1462),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1462),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1482),
.A2(n_1459),
.B1(n_1448),
.B2(n_1439),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1479),
.B(n_1399),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1480),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1471),
.B(n_1432),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1461),
.B(n_1403),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1471),
.B(n_1429),
.Y(n_1498)
);

CKINVDCx16_ASAP7_75t_R g1499 ( 
.A(n_1467),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1473),
.B(n_1429),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1469),
.B(n_1426),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1485),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1461),
.B(n_1403),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1483),
.B(n_1318),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1473),
.B(n_1458),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1460),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1460),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1460),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1463),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1463),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1466),
.B(n_1421),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1476),
.B(n_1465),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1474),
.B(n_1421),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1464),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1483),
.B(n_1310),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1486),
.B(n_1468),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1486),
.B(n_1474),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1497),
.B(n_1480),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1504),
.B(n_1330),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1502),
.B(n_1498),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1506),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1502),
.B(n_1477),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1498),
.B(n_1475),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1513),
.B(n_1470),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1494),
.B(n_1499),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1492),
.Y(n_1526)
);

NOR2xp67_ASAP7_75t_SL g1527 ( 
.A(n_1499),
.B(n_1296),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1506),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1513),
.B(n_1470),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1503),
.B(n_1478),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1496),
.B(n_1482),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1496),
.B(n_1467),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1487),
.B(n_1484),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1488),
.B(n_1422),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1492),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1488),
.B(n_1464),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1509),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1509),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1487),
.B(n_1484),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1493),
.A2(n_1453),
.B(n_1446),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1510),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1506),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1510),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1507),
.Y(n_1544)
);

NOR2xp67_ASAP7_75t_L g1545 ( 
.A(n_1495),
.B(n_1490),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1511),
.B(n_1484),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1491),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1491),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1500),
.B(n_1406),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1531),
.B(n_1507),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1520),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1533),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1524),
.B(n_1512),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1547),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1548),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1525),
.B(n_1515),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1533),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1525),
.B(n_1507),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1521),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1526),
.B(n_1505),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1521),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1528),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1524),
.B(n_1512),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1516),
.B(n_1495),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1540),
.A2(n_1493),
.B1(n_1508),
.B2(n_1489),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1528),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1516),
.B(n_1490),
.Y(n_1567)
);

AND2x6_ASAP7_75t_L g1568 ( 
.A(n_1518),
.B(n_1501),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1536),
.A2(n_1508),
.B(n_1489),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1535),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1537),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1518),
.B(n_1503),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1539),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1517),
.B(n_1495),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1551),
.B(n_1538),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1562),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_SL g1577 ( 
.A1(n_1551),
.A2(n_1560),
.B(n_1550),
.C(n_1522),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1567),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1565),
.A2(n_1532),
.B(n_1500),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1574),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1558),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1550),
.A2(n_1508),
.B1(n_1489),
.B2(n_1542),
.Y(n_1582)
);

A2O1A1Ixp33_ASAP7_75t_SL g1583 ( 
.A1(n_1558),
.A2(n_1544),
.B(n_1542),
.C(n_1527),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1562),
.Y(n_1584)
);

AOI221xp5_ASAP7_75t_L g1585 ( 
.A1(n_1558),
.A2(n_1544),
.B1(n_1505),
.B2(n_1523),
.C(n_1534),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1560),
.A2(n_1545),
.B(n_1519),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1554),
.Y(n_1587)
);

AOI211xp5_ASAP7_75t_L g1588 ( 
.A1(n_1556),
.A2(n_1546),
.B(n_1539),
.C(n_1549),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1553),
.B(n_1529),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1554),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1572),
.B(n_1517),
.Y(n_1591)
);

NAND2x1p5_ASAP7_75t_L g1592 ( 
.A(n_1561),
.B(n_1296),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1555),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1591),
.B(n_1564),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1581),
.B(n_1580),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1578),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1589),
.B(n_1561),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1585),
.B(n_1561),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1586),
.B(n_1564),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1577),
.B(n_1566),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1576),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1584),
.B(n_1566),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1575),
.B(n_1553),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1579),
.B(n_1559),
.Y(n_1604)
);

INVxp67_ASAP7_75t_SL g1605 ( 
.A(n_1604),
.Y(n_1605)
);

AOI221xp5_ASAP7_75t_L g1606 ( 
.A1(n_1604),
.A2(n_1582),
.B1(n_1583),
.B2(n_1588),
.C(n_1575),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1600),
.A2(n_1582),
.B(n_1559),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1598),
.A2(n_1529),
.B1(n_1572),
.B2(n_1567),
.Y(n_1608)
);

OAI211xp5_ASAP7_75t_L g1609 ( 
.A1(n_1597),
.A2(n_1595),
.B(n_1602),
.C(n_1599),
.Y(n_1609)
);

AOI211xp5_ASAP7_75t_L g1610 ( 
.A1(n_1603),
.A2(n_1559),
.B(n_1574),
.C(n_1552),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1594),
.A2(n_1569),
.B(n_1557),
.Y(n_1611)
);

AOI221x1_ASAP7_75t_L g1612 ( 
.A1(n_1601),
.A2(n_1571),
.B1(n_1570),
.B2(n_1590),
.C(n_1587),
.Y(n_1612)
);

NOR3xp33_ASAP7_75t_L g1613 ( 
.A(n_1596),
.B(n_1593),
.C(n_1571),
.Y(n_1613)
);

AOI31xp33_ASAP7_75t_L g1614 ( 
.A1(n_1605),
.A2(n_1592),
.A3(n_1570),
.B(n_1519),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1611),
.A2(n_1606),
.B(n_1607),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1610),
.A2(n_1592),
.B(n_1569),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1608),
.Y(n_1617)
);

NOR2x1_ASAP7_75t_L g1618 ( 
.A(n_1609),
.B(n_1555),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1618),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1617),
.B(n_1572),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1614),
.B(n_1563),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1615),
.B(n_1612),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1616),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1618),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1619),
.B(n_1613),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1620),
.B(n_1567),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1624),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1621),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_SL g1629 ( 
.A1(n_1622),
.A2(n_1541),
.B(n_1543),
.Y(n_1629)
);

OAI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1627),
.A2(n_1622),
.B1(n_1623),
.B2(n_1629),
.Y(n_1630)
);

NAND5xp2_ASAP7_75t_L g1631 ( 
.A(n_1628),
.B(n_1568),
.C(n_1347),
.D(n_1530),
.E(n_1455),
.Y(n_1631)
);

NOR3xp33_ASAP7_75t_L g1632 ( 
.A(n_1625),
.B(n_1573),
.C(n_1557),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1632),
.Y(n_1633)
);

AOI322xp5_ASAP7_75t_L g1634 ( 
.A1(n_1633),
.A2(n_1630),
.A3(n_1626),
.B1(n_1573),
.B2(n_1557),
.C1(n_1552),
.C2(n_1514),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1634),
.Y(n_1635)
);

NOR2xp67_ASAP7_75t_L g1636 ( 
.A(n_1634),
.B(n_1631),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1635),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1636),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1637),
.B(n_1552),
.Y(n_1639)
);

CKINVDCx20_ASAP7_75t_R g1640 ( 
.A(n_1638),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1639),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1641),
.Y(n_1642)
);

OAI211xp5_ASAP7_75t_L g1643 ( 
.A1(n_1642),
.A2(n_1640),
.B(n_1573),
.C(n_1301),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1643),
.A2(n_1569),
.B1(n_1568),
.B2(n_1563),
.Y(n_1644)
);

AOI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1644),
.A2(n_1320),
.B1(n_1514),
.B2(n_1313),
.C(n_1323),
.Y(n_1645)
);

AOI211xp5_ASAP7_75t_L g1646 ( 
.A1(n_1645),
.A2(n_1296),
.B(n_1546),
.C(n_1514),
.Y(n_1646)
);


endmodule