module fake_jpeg_24230_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_18),
.B1(n_31),
.B2(n_24),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_54),
.B1(n_16),
.B2(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_51),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_50),
.B1(n_57),
.B2(n_20),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_18),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_39),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_24),
.B1(n_31),
.B2(n_19),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_24),
.B1(n_31),
.B2(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_35),
.B1(n_41),
.B2(n_20),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_21),
.B(n_23),
.C(n_56),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_43),
.B1(n_34),
.B2(n_19),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_36),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_70),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_33),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_39),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_79),
.B(n_80),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_34),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_39),
.B(n_36),
.C(n_35),
.Y(n_80)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_44),
.B(n_39),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_85),
.B(n_48),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_84),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_55),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_87),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_95),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_92),
.B1(n_102),
.B2(n_84),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_93),
.B(n_99),
.Y(n_133)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_59),
.B1(n_36),
.B2(n_62),
.Y(n_92)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_36),
.B(n_35),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_56),
.B1(n_59),
.B2(n_58),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_106),
.B1(n_80),
.B2(n_64),
.Y(n_113)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_100),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_59),
.B1(n_16),
.B2(n_32),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_104),
.A2(n_110),
.B(n_28),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_61),
.B1(n_34),
.B2(n_30),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_66),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_112),
.B(n_29),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_102),
.B1(n_93),
.B2(n_106),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_114),
.A2(n_123),
.B1(n_124),
.B2(n_23),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_85),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_116),
.B(n_119),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_85),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_129),
.Y(n_160)
);

NAND2x1_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_36),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_78),
.B(n_82),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_125),
.B(n_130),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_89),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_65),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_77),
.B1(n_75),
.B2(n_83),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_107),
.B1(n_99),
.B2(n_93),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_81),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_75),
.C(n_77),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_65),
.C(n_70),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_81),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_100),
.B(n_87),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_22),
.B(n_109),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_137),
.B(n_27),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_86),
.B1(n_67),
.B2(n_111),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_163),
.B1(n_118),
.B2(n_113),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_140),
.B1(n_114),
.B2(n_123),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_93),
.B1(n_98),
.B2(n_103),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_98),
.B(n_72),
.C(n_101),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_143),
.B(n_147),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_101),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_155),
.C(n_157),
.Y(n_187)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_149),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_148),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_67),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_150),
.A2(n_158),
.B(n_162),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_67),
.Y(n_152)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_156),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_70),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_161),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_65),
.C(n_86),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_124),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_23),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_21),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_130),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_119),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_142),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_119),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_179),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_181),
.B1(n_157),
.B2(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_170),
.B(n_172),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_133),
.B1(n_130),
.B2(n_121),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_182),
.B1(n_184),
.B2(n_188),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_186),
.B1(n_139),
.B2(n_148),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_163),
.C(n_145),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_134),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_179),
.B(n_169),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_141),
.A2(n_133),
.B(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_127),
.B1(n_117),
.B2(n_28),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_180),
.C(n_181),
.Y(n_222)
);

OAI22x1_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_162),
.B1(n_147),
.B2(n_145),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_194),
.A2(n_205),
.B(n_206),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_164),
.B1(n_161),
.B2(n_150),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_165),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_208),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_178),
.Y(n_205)
);

XOR2x2_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_151),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_183),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_187),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_146),
.C(n_22),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_173),
.C(n_186),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_146),
.B1(n_0),
.B2(n_2),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_173),
.Y(n_225)
);

OAI21x1_ASAP7_75t_SL g211 ( 
.A1(n_166),
.A2(n_7),
.B(n_1),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_8),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_185),
.C(n_183),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_199),
.C(n_192),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_226),
.C(n_8),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_177),
.C(n_180),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_15),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_212),
.B1(n_194),
.B2(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_220),
.A2(n_193),
.B1(n_197),
.B2(n_209),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_234),
.B1(n_239),
.B2(n_213),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_241),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_168),
.B1(n_198),
.B2(n_203),
.Y(n_234)
);

BUFx12f_ASAP7_75t_SL g235 ( 
.A(n_221),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_218),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_240),
.C(n_10),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_9),
.C(n_3),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_226),
.C(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_244),
.B(n_246),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_216),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_0),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_223),
.C(n_224),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_250),
.C(n_11),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_228),
.C(n_0),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_9),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_252),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_235),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_253),
.A2(n_241),
.B1(n_238),
.B2(n_232),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_231),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_255),
.C(n_258),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_247),
.A2(n_240),
.B(n_236),
.C(n_6),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_257),
.B(n_260),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_261),
.B(n_11),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_263),
.B(n_261),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_245),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_266),
.B(n_267),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_243),
.Y(n_266)
);

NOR2x1_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_249),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_270),
.B(n_271),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_268),
.A2(n_257),
.B(n_254),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_268),
.Y(n_274)
);

OAI31xp33_ASAP7_75t_SL g275 ( 
.A1(n_274),
.A2(n_269),
.A3(n_258),
.B(n_15),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_273),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_12),
.B(n_14),
.Y(n_277)
);

OAI31xp33_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_12),
.A3(n_14),
.B(n_15),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_12),
.Y(n_279)
);


endmodule