module fake_jpeg_23254_n_348 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_46),
.Y(n_53)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx9p33_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_43),
.B(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_50),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_24),
.B1(n_31),
.B2(n_20),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_52),
.A2(n_64),
.B1(n_41),
.B2(n_39),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_24),
.B1(n_31),
.B2(n_36),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_41),
.B1(n_46),
.B2(n_39),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_24),
.B1(n_19),
.B2(n_21),
.Y(n_61)
);

OAI22x1_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_20),
.B1(n_18),
.B2(n_28),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_24),
.B1(n_41),
.B2(n_46),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_19),
.B(n_21),
.C(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_68),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_19),
.Y(n_67)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_26),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_73),
.A2(n_98),
.B(n_101),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_74),
.A2(n_84),
.B1(n_102),
.B2(n_62),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_75),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_83),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_36),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_81),
.A2(n_97),
.B1(n_32),
.B2(n_30),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_17),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_67),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_0),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_25),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_112)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_48),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_32),
.C(n_44),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_32),
.B1(n_29),
.B2(n_25),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_18),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_70),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_42),
.B1(n_48),
.B2(n_45),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_36),
.B1(n_25),
.B2(n_29),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_68),
.B1(n_57),
.B2(n_66),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_110),
.B1(n_131),
.B2(n_119),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_57),
.B1(n_70),
.B2(n_55),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_130),
.B(n_85),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_117),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_60),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_121),
.B(n_17),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_55),
.B1(n_60),
.B2(n_48),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_104),
.B1(n_100),
.B2(n_84),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_130),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_80),
.C(n_105),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_0),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_78),
.A2(n_30),
.B1(n_22),
.B2(n_23),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_135),
.B1(n_84),
.B2(n_102),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_74),
.A2(n_22),
.B1(n_34),
.B2(n_33),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_85),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_138),
.C(n_145),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_94),
.C(n_73),
.Y(n_138)
);

XOR2x2_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_165),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_116),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_140),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_79),
.B1(n_86),
.B2(n_92),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_153),
.B1(n_124),
.B2(n_125),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_94),
.A3(n_101),
.B1(n_87),
.B2(n_90),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_17),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_76),
.B(n_75),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_128),
.B(n_114),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_129),
.B1(n_133),
.B2(n_120),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_166),
.B(n_119),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_109),
.A2(n_104),
.B1(n_106),
.B2(n_81),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_88),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_44),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_44),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_160),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_37),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_37),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_110),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_96),
.B1(n_28),
.B2(n_11),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_118),
.B(n_23),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_182),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_187),
.B(n_200),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_193),
.B1(n_196),
.B2(n_201),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_112),
.A3(n_129),
.B1(n_120),
.B2(n_115),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_115),
.C(n_124),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_170),
.C(n_188),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_169),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_199),
.B1(n_164),
.B2(n_157),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_34),
.B(n_33),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_152),
.B(n_166),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_140),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_191),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_144),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_195),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_133),
.B1(n_125),
.B2(n_95),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_28),
.B1(n_5),
.B2(n_11),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_159),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_1),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_142),
.A2(n_95),
.B1(n_96),
.B2(n_28),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_138),
.A2(n_0),
.B(n_1),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_153),
.B(n_165),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_204),
.A2(n_187),
.B(n_196),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_205),
.A2(n_212),
.B1(n_220),
.B2(n_228),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_207),
.B(n_221),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_168),
.B(n_170),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_226),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_210),
.A2(n_190),
.B(n_168),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_141),
.B1(n_150),
.B2(n_156),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_139),
.Y(n_214)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_160),
.B(n_2),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_187),
.B(n_175),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_177),
.A2(n_1),
.B(n_2),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_218),
.A2(n_174),
.B(n_172),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_173),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_222),
.B(n_223),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_227),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_16),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_183),
.C(n_172),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_229)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_240),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_249),
.C(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_241),
.Y(n_262)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_202),
.A2(n_186),
.B(n_174),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_213),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_182),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_247),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_256),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_230),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_202),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_176),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_187),
.B(n_6),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_266),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_228),
.Y(n_261)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_231),
.C(n_214),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_268),
.C(n_263),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_205),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_208),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_212),
.C(n_210),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_215),
.Y(n_269)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_220),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_218),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_275),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_204),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_276),
.B(n_250),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_239),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_240),
.B(n_238),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_289),
.C(n_290),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_221),
.B(n_258),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_286),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_246),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_287),
.B(n_297),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_236),
.C(n_234),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_254),
.C(n_243),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_247),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_292),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_266),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

BUFx12_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_270),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_254),
.C(n_248),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_277),
.C(n_278),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_259),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_296),
.A2(n_260),
.B1(n_262),
.B2(n_223),
.Y(n_299)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_307),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_281),
.A2(n_251),
.B(n_256),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_305),
.C(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_310),
.Y(n_314)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_3),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_278),
.C(n_274),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_255),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_289),
.A2(n_203),
.B1(n_204),
.B2(n_241),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_290),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_313),
.B(n_321),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_280),
.Y(n_315)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_304),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_318),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_293),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_288),
.C(n_283),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_322),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_211),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_320),
.B(n_299),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_325),
.B(n_331),
.C(n_332),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_324),
.A2(n_306),
.B1(n_298),
.B2(n_302),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_326),
.B(n_327),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_316),
.Y(n_330)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_330),
.A2(n_9),
.B(n_12),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_314),
.A2(n_302),
.B(n_305),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_308),
.C(n_307),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_322),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_334),
.B(n_335),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_323),
.B(n_300),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_333),
.B(n_312),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_339),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_12),
.Y(n_340)
);

AOI21x1_ASAP7_75t_L g342 ( 
.A1(n_340),
.A2(n_330),
.B(n_14),
.Y(n_342)
);

AOI31xp33_ASAP7_75t_L g344 ( 
.A1(n_342),
.A2(n_339),
.A3(n_16),
.B(n_13),
.Y(n_344)
);

NOR2x1_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_341),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_337),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_346),
.A2(n_343),
.B(n_336),
.Y(n_347)
);

FAx1_ASAP7_75t_SL g348 ( 
.A(n_347),
.B(n_16),
.CI(n_337),
.CON(n_348),
.SN(n_348)
);


endmodule