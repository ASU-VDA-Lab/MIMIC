module real_aes_15332_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_911, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_911;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_0), .Y(n_533) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_1), .A2(n_53), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g237 ( .A(n_1), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_2), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g196 ( .A(n_3), .B(n_186), .Y(n_196) );
BUFx6f_ASAP7_75t_SL g525 ( .A(n_4), .Y(n_525) );
NAND2xp33_ASAP7_75t_L g657 ( .A(n_5), .B(n_184), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g229 ( .A1(n_6), .A2(n_101), .B1(n_217), .B2(n_230), .C(n_231), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_7), .A2(n_105), .B1(n_900), .B2(n_908), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_8), .B(n_171), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_9), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_10), .B(n_140), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_11), .B(n_175), .Y(n_174) );
AOI21xp33_ASAP7_75t_L g537 ( .A1(n_12), .A2(n_532), .B(n_538), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_13), .Y(n_672) );
BUFx3_ASAP7_75t_L g142 ( .A(n_14), .Y(n_142) );
INVx1_ASAP7_75t_L g153 ( .A(n_14), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_15), .B(n_155), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_16), .A2(n_187), .B(n_579), .C(n_633), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_17), .Y(n_279) );
BUFx10_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_19), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_20), .B(n_262), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_21), .A2(n_524), .B1(n_525), .B2(n_526), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_21), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_22), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_23), .B(n_163), .Y(n_276) );
OAI21xp33_ASAP7_75t_L g320 ( .A1(n_23), .A2(n_70), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_24), .B(n_260), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_25), .A2(n_548), .B1(n_551), .B2(n_552), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_25), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_26), .B(n_600), .Y(n_599) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_27), .A2(n_624), .B(n_625), .C(n_627), .Y(n_623) );
O2A1O1Ixp5_ASAP7_75t_L g232 ( .A1(n_28), .A2(n_188), .B(n_222), .C(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g610 ( .A(n_29), .B(n_171), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_30), .B(n_163), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_31), .A2(n_80), .B1(n_140), .B2(n_144), .Y(n_680) );
INVx1_ASAP7_75t_L g161 ( .A(n_32), .Y(n_161) );
INVx1_ASAP7_75t_L g646 ( .A(n_33), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_34), .B(n_145), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_35), .B(n_144), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_36), .B(n_163), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_37), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g121 ( .A(n_38), .Y(n_121) );
AND3x2_ASAP7_75t_L g542 ( .A(n_38), .B(n_543), .C(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_39), .B(n_217), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_40), .B(n_163), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_41), .B(n_222), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_42), .B(n_155), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_43), .Y(n_634) );
AND2x4_ASAP7_75t_L g160 ( .A(n_44), .B(n_161), .Y(n_160) );
NAND2x1_ASAP7_75t_L g185 ( .A(n_45), .B(n_186), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_46), .Y(n_285) );
INVx1_ASAP7_75t_L g180 ( .A(n_47), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_48), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_49), .A2(n_59), .B1(n_549), .B2(n_550), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_49), .Y(n_549) );
AND2x2_ASAP7_75t_L g195 ( .A(n_50), .B(n_151), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_51), .B(n_144), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_52), .A2(n_95), .B1(n_144), .B2(n_587), .Y(n_678) );
INVx1_ASAP7_75t_L g236 ( .A(n_53), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_54), .B(n_171), .Y(n_266) );
INVx1_ASAP7_75t_L g136 ( .A(n_55), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_56), .B(n_151), .Y(n_202) );
AND2x4_ASAP7_75t_L g906 ( .A(n_57), .B(n_907), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_58), .B(n_163), .Y(n_310) );
INVx1_ASAP7_75t_L g550 ( .A(n_59), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_60), .B(n_184), .Y(n_183) );
NOR2xp67_ASAP7_75t_L g122 ( .A(n_61), .B(n_83), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_62), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g605 ( .A(n_63), .B(n_164), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_64), .B(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_65), .B(n_600), .Y(n_617) );
INVx1_ASAP7_75t_L g907 ( .A(n_66), .Y(n_907) );
NAND2x1_ASAP7_75t_L g578 ( .A(n_67), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g200 ( .A(n_68), .B(n_171), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_69), .B(n_155), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_70), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_71), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_72), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_73), .B(n_144), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_74), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_75), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_76), .B(n_251), .Y(n_639) );
INVx2_ASAP7_75t_L g119 ( .A(n_77), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_78), .B(n_214), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_79), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_81), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_82), .B(n_217), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_84), .B(n_163), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_85), .A2(n_522), .B1(n_523), .B2(n_527), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_85), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_86), .B(n_164), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_87), .B(n_151), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_88), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_89), .B(n_262), .Y(n_575) );
NAND2xp33_ASAP7_75t_SL g641 ( .A(n_90), .B(n_263), .Y(n_641) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_91), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_92), .B(n_151), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_93), .B(n_216), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_94), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g148 ( .A(n_96), .Y(n_148) );
BUFx3_ASAP7_75t_L g158 ( .A(n_96), .Y(n_158) );
INVx1_ASAP7_75t_L g189 ( .A(n_96), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_97), .B(n_286), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_98), .Y(n_626) );
INVx1_ASAP7_75t_L g113 ( .A(n_99), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_99), .B(n_530), .Y(n_529) );
NAND2xp33_ASAP7_75t_L g654 ( .A(n_100), .B(n_181), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_102), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_103), .B(n_151), .Y(n_614) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_545), .Y(n_105) );
OAI21xp33_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_112), .B(n_537), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
CKINVDCx11_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_111), .B(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g899 ( .A(n_111), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_114), .B(n_528), .Y(n_112) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_123), .Y(n_114) );
BUFx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx12f_ASAP7_75t_L g530 ( .A(n_116), .Y(n_530) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g536 ( .A(n_117), .Y(n_536) );
NOR2x1p5_ASAP7_75t_L g117 ( .A(n_118), .B(n_120), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g543 ( .A(n_119), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
BUFx2_ASAP7_75t_L g558 ( .A(n_121), .Y(n_558) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_122), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_123), .A2(n_529), .B(n_531), .Y(n_528) );
XOR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_521), .Y(n_123) );
XNOR2xp5_ASAP7_75t_L g559 ( .A(n_124), .B(n_526), .Y(n_559) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_450), .Y(n_124) );
NOR3xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_397), .C(n_427), .Y(n_125) );
NAND4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_325), .C(n_364), .D(n_377), .Y(n_126) );
AOI332xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_225), .A3(n_242), .B1(n_267), .B2(n_272), .B3(n_293), .C1(n_311), .C2(n_315), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_191), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_166), .Y(n_129) );
INVx2_ASAP7_75t_L g268 ( .A(n_130), .Y(n_268) );
AND2x2_ASAP7_75t_L g382 ( .A(n_130), .B(n_167), .Y(n_382) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx3_ASAP7_75t_L g337 ( .A(n_131), .Y(n_337) );
OAI21x1_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_137), .B(n_162), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_133), .A2(n_159), .B(n_645), .Y(n_648) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx3_ASAP7_75t_L g321 ( .A(n_134), .Y(n_321) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_135), .Y(n_171) );
INVxp33_ASAP7_75t_L g647 ( .A(n_135), .Y(n_647) );
INVx1_ASAP7_75t_L g238 ( .A(n_136), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_149), .B(n_159), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B(n_146), .Y(n_138) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_141), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g251 ( .A(n_141), .Y(n_251) );
INVx2_ASAP7_75t_L g260 ( .A(n_141), .Y(n_260) );
INVx2_ASAP7_75t_L g286 ( .A(n_141), .Y(n_286) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g145 ( .A(n_142), .Y(n_145) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_142), .Y(n_156) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
INVx1_ASAP7_75t_L g214 ( .A(n_145), .Y(n_214) );
INVx2_ASAP7_75t_L g281 ( .A(n_145), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_146), .A2(n_213), .B(n_215), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_146), .A2(n_258), .B(n_261), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_146), .A2(n_306), .B(n_308), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_146), .A2(n_574), .B(n_575), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_146), .A2(n_589), .B(n_591), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_146), .A2(n_616), .B(n_617), .Y(n_615) );
AO21x1_ASAP7_75t_L g637 ( .A1(n_146), .A2(n_638), .B(n_639), .Y(n_637) );
BUFx10_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx3_ASAP7_75t_L g231 ( .A(n_148), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_154), .B(n_157), .Y(n_149) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx2_ASAP7_75t_L g222 ( .A(n_152), .Y(n_222) );
INVx2_ASAP7_75t_L g263 ( .A(n_152), .Y(n_263) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
INVx3_ASAP7_75t_L g186 ( .A(n_156), .Y(n_186) );
INVx2_ASAP7_75t_L g587 ( .A(n_156), .Y(n_587) );
INVx2_ASAP7_75t_L g600 ( .A(n_156), .Y(n_600) );
INVx2_ASAP7_75t_L g643 ( .A(n_156), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_157), .A2(n_585), .B(n_586), .Y(n_584) );
AO21x1_ASAP7_75t_L g640 ( .A1(n_157), .A2(n_641), .B(n_642), .Y(n_640) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g175 ( .A(n_158), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_158), .B(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g283 ( .A(n_158), .Y(n_283) );
AOI211x1_ASAP7_75t_L g611 ( .A1(n_158), .A2(n_610), .B(n_612), .C(n_615), .Y(n_611) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_159), .A2(n_173), .B(n_182), .Y(n_172) );
INVx1_ASAP7_75t_L g224 ( .A(n_159), .Y(n_224) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_159), .A2(n_584), .B(n_588), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_159), .A2(n_609), .B(n_610), .Y(n_608) );
OAI21x1_ASAP7_75t_L g651 ( .A1(n_159), .A2(n_652), .B(n_655), .Y(n_651) );
BUFx6f_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g208 ( .A(n_160), .Y(n_208) );
INVx2_ASAP7_75t_L g265 ( .A(n_160), .Y(n_265) );
INVx1_ASAP7_75t_L g290 ( .A(n_160), .Y(n_290) );
INVx1_ASAP7_75t_L g676 ( .A(n_160), .Y(n_676) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_164), .B(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g388 ( .A(n_166), .B(n_337), .Y(n_388) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g271 ( .A(n_167), .Y(n_271) );
AND2x4_ASAP7_75t_SL g312 ( .A(n_167), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_167), .B(n_193), .Y(n_340) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_167), .Y(n_358) );
AND2x2_ASAP7_75t_L g384 ( .A(n_167), .B(n_337), .Y(n_384) );
INVx1_ASAP7_75t_L g431 ( .A(n_167), .Y(n_431) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_190), .Y(n_168) );
INVx1_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVxp33_ASAP7_75t_L g206 ( .A(n_171), .Y(n_206) );
INVx1_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_171), .Y(n_247) );
NOR2xp67_ASAP7_75t_SL g596 ( .A(n_171), .B(n_290), .Y(n_596) );
INVxp67_ASAP7_75t_SL g609 ( .A(n_171), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_176), .B(n_178), .Y(n_173) );
INVx1_ASAP7_75t_L g627 ( .A(n_175), .Y(n_627) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_181), .Y(n_178) );
AOI21x1_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_185), .B(n_187), .Y(n_182) );
INVx1_ASAP7_75t_L g303 ( .A(n_184), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_187), .A2(n_220), .B(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g304 ( .A(n_188), .Y(n_304) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx3_ASAP7_75t_L g198 ( .A(n_189), .Y(n_198) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g354 ( .A(n_192), .Y(n_354) );
INVx1_ASAP7_75t_L g485 ( .A(n_192), .Y(n_485) );
OR2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_209), .Y(n_192) );
INVx2_ASAP7_75t_L g313 ( .A(n_193), .Y(n_313) );
AND2x2_ASAP7_75t_L g359 ( .A(n_193), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g414 ( .A(n_193), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_193), .B(n_431), .Y(n_462) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_199), .B(n_205), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .Y(n_194) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g204 ( .A(n_198), .Y(n_204) );
O2A1O1Ixp5_ASAP7_75t_L g576 ( .A1(n_198), .A2(n_250), .B(n_577), .C(n_578), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_198), .B(n_324), .C(n_675), .Y(n_679) );
NOR2xp67_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
AOI21xp33_ASAP7_75t_L g205 ( .A1(n_200), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_204), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_204), .A2(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR3xp33_ASAP7_75t_L g228 ( .A(n_208), .B(n_229), .C(n_232), .Y(n_228) );
INVx1_ASAP7_75t_L g270 ( .A(n_209), .Y(n_270) );
AND2x2_ASAP7_75t_L g335 ( .A(n_209), .B(n_336), .Y(n_335) );
INVx3_ASAP7_75t_L g360 ( .A(n_209), .Y(n_360) );
INVx1_ASAP7_75t_L g381 ( .A(n_209), .Y(n_381) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_209), .Y(n_385) );
AND2x2_ASAP7_75t_L g395 ( .A(n_209), .B(n_313), .Y(n_395) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_219), .B(n_223), .Y(n_211) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g624 ( .A(n_217), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_217), .B(n_634), .Y(n_633) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx3_ASAP7_75t_L g230 ( .A(n_218), .Y(n_230) );
INVx1_ASAP7_75t_L g437 ( .A(n_225), .Y(n_437) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g295 ( .A(n_226), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g446 ( .A(n_226), .B(n_420), .Y(n_446) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g331 ( .A(n_227), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g370 ( .A(n_227), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g403 ( .A(n_227), .B(n_297), .Y(n_403) );
INVx1_ASAP7_75t_L g493 ( .A(n_227), .Y(n_493) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_235), .B(n_239), .Y(n_227) );
NAND2xp33_ASAP7_75t_L g322 ( .A(n_228), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g307 ( .A(n_230), .Y(n_307) );
INVx2_ASAP7_75t_L g579 ( .A(n_230), .Y(n_579) );
INVx2_ASAP7_75t_L g590 ( .A(n_230), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_230), .B(n_626), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_231), .A2(n_250), .B1(n_252), .B2(n_256), .Y(n_249) );
INVx2_ASAP7_75t_SL g255 ( .A(n_231), .Y(n_255) );
INVx1_ASAP7_75t_L g288 ( .A(n_231), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_235), .B(n_264), .Y(n_628) );
INVx2_ASAP7_75t_L g630 ( .A(n_235), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_235), .B(n_672), .Y(n_671) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_238), .Y(n_235) );
AOI21x1_ASAP7_75t_L g291 ( .A1(n_236), .A2(n_237), .B(n_238), .Y(n_291) );
NOR2xp33_ASAP7_75t_R g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_244), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g369 ( .A(n_244), .Y(n_369) );
INVx2_ASAP7_75t_L g391 ( .A(n_244), .Y(n_391) );
OR2x2_ASAP7_75t_L g465 ( .A(n_244), .B(n_319), .Y(n_465) );
AND2x2_ASAP7_75t_L g504 ( .A(n_244), .B(n_295), .Y(n_504) );
BUFx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g344 ( .A(n_245), .Y(n_344) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_248), .B(n_266), .Y(n_245) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_246), .A2(n_248), .B(n_266), .Y(n_292) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_246), .A2(n_299), .B(n_310), .Y(n_298) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_246), .A2(n_299), .B(n_310), .Y(n_332) );
OAI21x1_ASAP7_75t_L g571 ( .A1(n_246), .A2(n_572), .B(n_580), .Y(n_571) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_246), .A2(n_583), .B(n_592), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_246), .A2(n_583), .B(n_592), .Y(n_719) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_257), .B(n_264), .Y(n_248) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OAI221xp5_ASAP7_75t_L g284 ( .A1(n_263), .A2(n_285), .B1(n_286), .B2(n_287), .C(n_288), .Y(n_284) );
INVx2_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g309 ( .A(n_265), .Y(n_309) );
NOR2x1_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g314 ( .A(n_268), .Y(n_314) );
AND2x2_ASAP7_75t_L g436 ( .A(n_268), .B(n_421), .Y(n_436) );
AND2x2_ASAP7_75t_L g441 ( .A(n_268), .B(n_312), .Y(n_441) );
AND2x2_ASAP7_75t_L g516 ( .A(n_268), .B(n_359), .Y(n_516) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g408 ( .A(n_270), .Y(n_408) );
INVx1_ASAP7_75t_L g467 ( .A(n_271), .Y(n_467) );
AND2x2_ASAP7_75t_L g482 ( .A(n_271), .B(n_483), .Y(n_482) );
OAI211xp5_ASAP7_75t_SL g500 ( .A1(n_272), .A2(n_501), .B(n_503), .C(n_505), .Y(n_500) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_SL g386 ( .A(n_273), .B(n_295), .Y(n_386) );
AND2x2_ASAP7_75t_L g426 ( .A(n_273), .B(n_331), .Y(n_426) );
AND2x2_ASAP7_75t_L g438 ( .A(n_273), .B(n_403), .Y(n_438) );
AND2x2_ASAP7_75t_L g445 ( .A(n_273), .B(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_292), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g330 ( .A(n_275), .Y(n_330) );
AND2x2_ASAP7_75t_L g343 ( .A(n_275), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g372 ( .A(n_275), .Y(n_372) );
AND2x2_ASAP7_75t_L g475 ( .A(n_275), .B(n_292), .Y(n_475) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NAND3xp33_ASAP7_75t_L g319 ( .A(n_277), .B(n_320), .C(n_322), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_284), .C(n_289), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B(n_282), .C(n_283), .Y(n_278) );
INVx2_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_283), .A2(n_603), .B(n_604), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_283), .A2(n_653), .B(n_654), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx2_ASAP7_75t_L g324 ( .A(n_291), .Y(n_324) );
INVx1_ASAP7_75t_L g422 ( .A(n_292), .Y(n_422) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_293), .A2(n_421), .B(n_441), .C(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g345 ( .A(n_296), .Y(n_345) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVxp67_ASAP7_75t_L g317 ( .A(n_298), .Y(n_317) );
OAI21x1_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_305), .B(n_309), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B(n_304), .Y(n_300) );
INVx1_ASAP7_75t_L g677 ( .A(n_304), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_307), .A2(n_613), .B(n_614), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g572 ( .A1(n_309), .A2(n_573), .B(n_576), .Y(n_572) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx2_ASAP7_75t_L g479 ( .A(n_312), .Y(n_479) );
AND2x2_ASAP7_75t_L g499 ( .A(n_312), .B(n_385), .Y(n_499) );
BUFx2_ASAP7_75t_L g448 ( .A(n_313), .Y(n_448) );
OR2x2_ASAP7_75t_L g461 ( .A(n_314), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g509 ( .A(n_315), .Y(n_509) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g367 ( .A(n_316), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_316), .B(n_368), .Y(n_396) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g362 ( .A(n_317), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g363 ( .A(n_319), .Y(n_363) );
OR2x2_ASAP7_75t_L g390 ( .A(n_319), .B(n_391), .Y(n_390) );
OAI21x1_ASAP7_75t_L g650 ( .A1(n_321), .A2(n_651), .B(n_658), .Y(n_650) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_324), .B(n_675), .C(n_677), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_333), .B1(n_341), .B2(n_346), .C(n_348), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g421 ( .A(n_330), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g432 ( .A(n_331), .B(n_369), .Y(n_432) );
AND2x2_ASAP7_75t_L g468 ( .A(n_331), .B(n_421), .Y(n_468) );
AND2x2_ASAP7_75t_L g515 ( .A(n_331), .B(n_475), .Y(n_515) );
INVx1_ASAP7_75t_L g420 ( .A(n_332), .Y(n_420) );
NOR2xp67_ASAP7_75t_SL g333 ( .A(n_334), .B(n_338), .Y(n_333) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_334), .B(n_413), .C(n_460), .D(n_461), .Y(n_459) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g346 ( .A(n_335), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_335), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g352 ( .A(n_336), .Y(n_352) );
INVx1_ASAP7_75t_L g394 ( .A(n_336), .Y(n_394) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_336), .Y(n_449) );
AND2x2_ASAP7_75t_L g458 ( .A(n_336), .B(n_347), .Y(n_458) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g483 ( .A(n_337), .B(n_414), .Y(n_483) );
INVx1_ASAP7_75t_L g406 ( .A(n_338), .Y(n_406) );
BUFx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g424 ( .A(n_339), .B(n_381), .Y(n_424) );
AND2x4_ASAP7_75t_L g439 ( .A(n_339), .B(n_408), .Y(n_439) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g347 ( .A(n_340), .Y(n_347) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_343), .B(n_403), .Y(n_410) );
INVx1_ASAP7_75t_L g507 ( .A(n_343), .Y(n_507) );
BUFx3_ASAP7_75t_L g401 ( .A(n_344), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_345), .B(n_436), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_353), .B(n_355), .C(n_361), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI21xp33_ASAP7_75t_L g508 ( .A1(n_351), .A2(n_509), .B(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g376 ( .A(n_352), .Y(n_376) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g387 ( .A(n_354), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g429 ( .A(n_354), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g433 ( .A(n_354), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2x1_ASAP7_75t_L g374 ( .A(n_356), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_358), .Y(n_416) );
INVx1_ASAP7_75t_L g398 ( .A(n_359), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_359), .B(n_376), .Y(n_473) );
OR2x2_ASAP7_75t_L g413 ( .A(n_360), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g488 ( .A(n_360), .Y(n_488) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_370), .B(n_373), .Y(n_364) );
INVxp33_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_370), .A2(n_429), .B1(n_432), .B2(n_433), .Y(n_428) );
AND2x2_ASAP7_75t_L g402 ( .A(n_371), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g456 ( .A(n_371), .Y(n_456) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI222xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_386), .B1(n_387), .B2(n_389), .C1(n_392), .C2(n_396), .Y(n_377) );
NAND2xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_383), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
AND2x2_ASAP7_75t_L g425 ( .A(n_381), .B(n_384), .Y(n_425) );
AND2x2_ASAP7_75t_L g496 ( .A(n_381), .B(n_467), .Y(n_496) );
INVx1_ASAP7_75t_L g460 ( .A(n_382), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_384), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_388), .B(n_412), .Y(n_443) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_392), .A2(n_426), .B1(n_515), .B2(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
OAI211xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B(n_404), .C(n_423), .Y(n_397) );
NAND2x1p5_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_402), .A2(n_441), .B1(n_445), .B2(n_447), .Y(n_444) );
INVx1_ASAP7_75t_L g502 ( .A(n_403), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_409), .B1(n_411), .B2(n_417), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
AND2x2_ASAP7_75t_L g457 ( .A(n_407), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g520 ( .A(n_408), .B(n_479), .Y(n_520) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .Y(n_411) );
AOI32xp33_ASAP7_75t_L g435 ( .A1(n_412), .A2(n_436), .A3(n_437), .B1(n_438), .B2(n_439), .Y(n_435) );
INVx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx2_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_421), .B(n_437), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_421), .B(n_455), .Y(n_510) );
OAI21xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B(n_426), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_424), .A2(n_499), .B1(n_500), .B2(n_508), .Y(n_498) );
NAND4xp25_ASAP7_75t_SL g427 ( .A(n_428), .B(n_435), .C(n_440), .D(n_444), .Y(n_427) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_437), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_SL g486 ( .A(n_438), .Y(n_486) );
OAI21xp5_ASAP7_75t_SL g487 ( .A1(n_438), .A2(n_488), .B(n_489), .Y(n_487) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_497), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_469), .C(n_487), .Y(n_451) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_457), .B1(n_459), .B2(n_463), .C1(n_466), .C2(n_468), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
OR2x2_ASAP7_75t_L g464 ( .A(n_455), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g474 ( .A(n_455), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g518 ( .A(n_465), .Y(n_518) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_472), .B1(n_474), .B2(n_476), .C(n_480), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g491 ( .A(n_475), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_484), .B(n_486), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_488), .A2(n_490), .B(n_494), .C(n_496), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_488), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND4xp25_ASAP7_75t_L g497 ( .A(n_498), .B(n_511), .C(n_514), .D(n_517), .Y(n_497) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVxp67_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
OAI21xp33_ASAP7_75t_SL g517 ( .A1(n_515), .A2(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g527 ( .A(n_523), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_525), .Y(n_526) );
INVxp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
BUFx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g901 ( .A(n_542), .B(n_902), .Y(n_901) );
AND2x2_ASAP7_75t_L g898 ( .A(n_543), .B(n_544), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_896), .Y(n_545) );
XNOR2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_553), .Y(n_546) );
INVx1_ASAP7_75t_L g552 ( .A(n_548), .Y(n_552) );
OAI21x1_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_559), .B(n_560), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_555), .Y(n_561) );
CKINVDCx10_ASAP7_75t_R g555 ( .A(n_556), .Y(n_555) );
BUFx6f_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_835), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_779), .Y(n_564) );
NAND4xp25_ASAP7_75t_L g565 ( .A(n_566), .B(n_695), .C(n_722), .D(n_747), .Y(n_565) );
AOI221x1_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_618), .B1(n_659), .B2(n_666), .C(n_683), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_593), .Y(n_567) );
INVx1_ASAP7_75t_L g790 ( .A(n_568), .Y(n_790) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g688 ( .A(n_569), .Y(n_688) );
OR2x2_ASAP7_75t_L g869 ( .A(n_569), .B(n_870), .Y(n_869) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_581), .Y(n_569) );
BUFx2_ASAP7_75t_L g704 ( .A(n_570), .Y(n_704) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g663 ( .A(n_571), .Y(n_663) );
INVx1_ASAP7_75t_L g745 ( .A(n_571), .Y(n_745) );
AND2x2_ASAP7_75t_L g665 ( .A(n_581), .B(n_594), .Y(n_665) );
INVx1_ASAP7_75t_L g778 ( .A(n_581), .Y(n_778) );
AND2x2_ASAP7_75t_L g809 ( .A(n_581), .B(n_745), .Y(n_809) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g711 ( .A(n_582), .B(n_594), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_593), .B(n_826), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_593), .B(n_809), .Y(n_834) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_606), .Y(n_593) );
INVx2_ASAP7_75t_L g718 ( .A(n_594), .Y(n_718) );
INVx1_ASAP7_75t_L g762 ( .A(n_594), .Y(n_762) );
AND2x4_ASAP7_75t_L g594 ( .A(n_595), .B(n_601), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_596), .A2(n_602), .B(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g687 ( .A(n_607), .Y(n_687) );
INVx1_ASAP7_75t_L g692 ( .A(n_607), .Y(n_692) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_607), .Y(n_703) );
BUFx2_ASAP7_75t_L g715 ( .A(n_607), .Y(n_715) );
AND2x2_ASAP7_75t_L g746 ( .A(n_607), .B(n_718), .Y(n_746) );
INVx2_ASAP7_75t_L g840 ( .A(n_607), .Y(n_840) );
AND2x2_ASAP7_75t_L g856 ( .A(n_607), .B(n_719), .Y(n_856) );
OR2x6_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_635), .Y(n_618) );
OR2x2_ASAP7_75t_L g758 ( .A(n_619), .B(n_721), .Y(n_758) );
NAND2x1p5_ASAP7_75t_L g819 ( .A(n_619), .B(n_820), .Y(n_819) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g708 ( .A(n_621), .Y(n_708) );
AND2x2_ASAP7_75t_L g739 ( .A(n_621), .B(n_740), .Y(n_739) );
BUFx2_ASAP7_75t_L g766 ( .A(n_621), .Y(n_766) );
AND2x2_ASAP7_75t_L g814 ( .A(n_621), .B(n_687), .Y(n_814) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_621), .Y(n_850) );
NAND2x1p5_ASAP7_75t_L g621 ( .A(n_622), .B(n_631), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g682 ( .A(n_622), .B(n_631), .Y(n_682) );
OA21x2_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_628), .B(n_629), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_627), .A2(n_656), .B(n_657), .Y(n_655) );
OR2x2_ASAP7_75t_L g631 ( .A(n_628), .B(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g721 ( .A(n_635), .Y(n_721) );
AND2x2_ASAP7_75t_L g801 ( .A(n_635), .B(n_753), .Y(n_801) );
AND2x2_ASAP7_75t_L g891 ( .A(n_635), .B(n_765), .Y(n_891) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_649), .Y(n_635) );
OR2x2_ASAP7_75t_L g681 ( .A(n_636), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g694 ( .A(n_636), .B(n_650), .Y(n_694) );
AND2x2_ASAP7_75t_L g707 ( .A(n_636), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g730 ( .A(n_636), .B(n_682), .Y(n_730) );
INVx2_ASAP7_75t_L g740 ( .A(n_636), .Y(n_740) );
INVx1_ASAP7_75t_L g787 ( .A(n_636), .Y(n_787) );
AO31x2_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_640), .A3(n_644), .B(n_648), .Y(n_636) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g742 ( .A(n_650), .Y(n_742) );
AND2x2_ASAP7_75t_L g767 ( .A(n_650), .B(n_670), .Y(n_767) );
INVx1_ASAP7_75t_L g794 ( .A(n_650), .Y(n_794) );
AND2x2_ASAP7_75t_L g847 ( .A(n_650), .B(n_822), .Y(n_847) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_664), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g691 ( .A(n_662), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g712 ( .A(n_662), .B(n_692), .Y(n_712) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g735 ( .A(n_663), .Y(n_735) );
OR2x2_ASAP7_75t_L g803 ( .A(n_664), .B(n_751), .Y(n_803) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g690 ( .A(n_665), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g886 ( .A(n_665), .B(n_686), .Y(n_886) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_681), .Y(n_667) );
OR2x2_ASAP7_75t_L g720 ( .A(n_668), .B(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g879 ( .A(n_668), .B(n_721), .Y(n_879) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g698 ( .A(n_670), .Y(n_698) );
INVxp67_ASAP7_75t_L g729 ( .A(n_670), .Y(n_729) );
AND2x2_ASAP7_75t_L g741 ( .A(n_670), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g753 ( .A(n_670), .Y(n_753) );
AND2x2_ASAP7_75t_L g775 ( .A(n_670), .B(n_682), .Y(n_775) );
INVx1_ASAP7_75t_L g822 ( .A(n_670), .Y(n_822) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_678), .B1(n_679), .B2(n_680), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g702 ( .A(n_681), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g754 ( .A(n_681), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_681), .B(n_800), .Y(n_799) );
OR2x2_ASAP7_75t_L g872 ( .A(n_681), .B(n_873), .Y(n_872) );
AND2x2_ASAP7_75t_L g737 ( .A(n_682), .B(n_698), .Y(n_737) );
INVx2_ASAP7_75t_L g868 ( .A(n_682), .Y(n_868) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_689), .B(n_693), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g875 ( .A(n_685), .B(n_749), .C(n_750), .Y(n_875) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_686), .B(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_686), .B(n_733), .Y(n_842) );
BUFx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g870 ( .A(n_687), .B(n_718), .Y(n_870) );
AND2x4_ASAP7_75t_SL g760 ( .A(n_688), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g812 ( .A(n_688), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_689), .A2(n_790), .B1(n_791), .B2(n_795), .Y(n_789) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g736 ( .A(n_694), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g774 ( .A(n_694), .B(n_775), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_699), .B(n_705), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_696), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_704), .Y(n_700) );
INVx2_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
OAI32xp33_ASAP7_75t_L g804 ( .A1(n_702), .A2(n_739), .A3(n_805), .B1(n_806), .B2(n_807), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_704), .B(n_871), .Y(n_893) );
OAI22xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B1(n_713), .B2(n_720), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_707), .B(n_808), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_707), .B(n_847), .Y(n_881) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR2x1_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx4_ASAP7_75t_L g749 ( .A(n_711), .Y(n_749) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_711), .Y(n_788) );
OR2x2_ASAP7_75t_L g828 ( .A(n_711), .B(n_744), .Y(n_828) );
INVx1_ASAP7_75t_L g726 ( .A(n_712), .Y(n_726) );
OR2x2_ASAP7_75t_L g805 ( .A(n_712), .B(n_761), .Y(n_805) );
OR2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
AND2x2_ASAP7_75t_L g833 ( .A(n_714), .B(n_717), .Y(n_833) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_715), .B(n_733), .Y(n_798) );
INVx1_ASAP7_75t_L g817 ( .A(n_715), .Y(n_817) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_717), .Y(n_725) );
AND2x2_ASAP7_75t_L g757 ( .A(n_717), .B(n_744), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_717), .B(n_817), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_717), .B(n_751), .Y(n_853) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
AND2x4_ASAP7_75t_SL g839 ( .A(n_718), .B(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g734 ( .A(n_719), .Y(n_734) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_727), .B1(n_731), .B2(n_736), .C1(n_738), .C2(n_743), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_726), .B(n_783), .Y(n_782) );
NOR4xp25_ASAP7_75t_L g885 ( .A(n_726), .B(n_809), .C(n_886), .D(n_887), .Y(n_885) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx2_ASAP7_75t_L g895 ( .A(n_730), .Y(n_895) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g826 ( .A(n_734), .Y(n_826) );
INVx2_ASAP7_75t_L g751 ( .A(n_735), .Y(n_751) );
INVx2_ASAP7_75t_L g795 ( .A(n_737), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_738), .A2(n_838), .B1(n_841), .B2(n_843), .Y(n_837) );
AND2x4_ASAP7_75t_SL g738 ( .A(n_739), .B(n_741), .Y(n_738) );
AND2x2_ASAP7_75t_L g843 ( .A(n_739), .B(n_767), .Y(n_843) );
INVx1_ASAP7_75t_L g846 ( .A(n_739), .Y(n_846) );
AND2x2_ASAP7_75t_L g821 ( .A(n_740), .B(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g858 ( .A(n_740), .Y(n_858) );
INVx1_ASAP7_75t_L g806 ( .A(n_741), .Y(n_806) );
AND2x2_ASAP7_75t_L g849 ( .A(n_741), .B(n_850), .Y(n_849) );
AND2x2_ASAP7_75t_L g867 ( .A(n_742), .B(n_868), .Y(n_867) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
HB1xp67_ASAP7_75t_L g883 ( .A(n_744), .Y(n_883) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g777 ( .A(n_745), .B(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g888 ( .A(n_746), .Y(n_888) );
AOI211xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_752), .B(n_755), .C(n_768), .Y(n_747) );
NOR2x1_ASAP7_75t_L g861 ( .A(n_748), .B(n_862), .Y(n_861) );
AOI322xp5_ASAP7_75t_L g877 ( .A1(n_748), .A2(n_749), .A3(n_814), .B1(n_878), .B2(n_880), .C1(n_882), .C2(n_911), .Y(n_877) );
AND2x4_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g838 ( .A(n_751), .B(n_839), .Y(n_838) );
OR2x2_ASAP7_75t_L g863 ( .A(n_751), .B(n_864), .Y(n_863) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_753), .Y(n_771) );
INVx2_ASAP7_75t_L g890 ( .A(n_753), .Y(n_890) );
INVx1_ASAP7_75t_L g831 ( .A(n_754), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_758), .B1(n_759), .B2(n_763), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g854 ( .A1(n_756), .A2(n_773), .B1(n_855), .B2(n_857), .Y(n_854) );
INVx2_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g871 ( .A(n_761), .Y(n_871) );
INVx4_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_767), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g772 ( .A(n_766), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_767), .B(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g873 ( .A(n_767), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_773), .B(n_776), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x4_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND4xp25_ASAP7_75t_L g779 ( .A(n_780), .B(n_796), .C(n_810), .D(n_823), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_788), .B(n_789), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_787), .B(n_793), .Y(n_792) );
INVx2_ASAP7_75t_L g829 ( .A(n_791), .Y(n_829) );
OR2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_795), .Y(n_791) );
INVxp67_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
BUFx3_ASAP7_75t_L g800 ( .A(n_794), .Y(n_800) );
AOI221xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_799), .B1(n_801), .B2(n_802), .C(n_804), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g808 ( .A(n_800), .Y(n_808) );
AND2x2_ASAP7_75t_L g820 ( .A(n_800), .B(n_821), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_800), .B(n_895), .Y(n_894) );
AND2x2_ASAP7_75t_L g813 ( .A(n_801), .B(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
O2A1O1Ixp33_ASAP7_75t_L g830 ( .A1(n_806), .A2(n_831), .B(n_832), .C(n_834), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_813), .B1(n_815), .B2(n_818), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g876 ( .A(n_821), .Y(n_876) );
O2A1O1Ixp33_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_827), .B(n_829), .C(n_830), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_829), .A2(n_838), .B1(n_893), .B2(n_894), .Y(n_892) );
INVxp67_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NOR3xp33_ASAP7_75t_L g835 ( .A(n_836), .B(n_874), .C(n_884), .Y(n_835) );
NAND3xp33_ASAP7_75t_SL g836 ( .A(n_837), .B(n_844), .C(n_859), .Y(n_836) );
INVx1_ASAP7_75t_L g864 ( .A(n_839), .Y(n_864) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_843), .A2(n_860), .B(n_865), .Y(n_859) );
AOI21xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_852), .B(n_854), .Y(n_844) );
OAI211xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_847), .B(n_848), .C(n_851), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_847), .B(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_869), .B1(n_871), .B2(n_872), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
OAI21xp33_ASAP7_75t_SL g874 ( .A1(n_875), .A2(n_876), .B(n_877), .Y(n_874) );
INVx2_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
OAI21xp33_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_889), .B(n_892), .Y(n_884) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
BUFx8_ASAP7_75t_SL g896 ( .A(n_897), .Y(n_896) );
OR2x6_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
BUFx8_ASAP7_75t_SL g900 ( .A(n_901), .Y(n_900) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_901), .Y(n_909) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx4_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
endmodule