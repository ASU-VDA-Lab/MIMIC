module fake_netlist_6_3576_n_2450 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2450);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2450;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_873;
wire n_461;
wire n_1285;
wire n_1371;
wire n_383;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_343;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_437;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_462;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_2442;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2301;
wire n_2209;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_374;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_137),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_98),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_23),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_30),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_69),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_232),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_87),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_116),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_32),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_78),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_101),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_5),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_32),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_87),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_56),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_42),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_19),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_48),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_121),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_176),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_115),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_154),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_221),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_62),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_224),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_78),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_33),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_201),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_37),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_85),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_97),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_129),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_159),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_14),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_17),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_86),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_46),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_14),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_160),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_114),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_72),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_165),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_75),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_199),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_95),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_211),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_169),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_43),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_226),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_185),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_84),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_94),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_147),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_158),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_179),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_101),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_16),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_80),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_118),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_106),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_132),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_23),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_33),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_80),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_84),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_58),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_153),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_122),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_89),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_143),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_18),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_202),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_123),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_53),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_141),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_131),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_48),
.Y(n_328)
);

INVxp33_ASAP7_75t_R g329 ( 
.A(n_42),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_229),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_44),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_220),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_37),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_69),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_93),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_26),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_112),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_227),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_184),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_151),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_168),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_28),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_108),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_150),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_83),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_117),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_198),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_10),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_4),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_124),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_106),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_13),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_81),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_99),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_130),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_3),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_52),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_61),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_4),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_100),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_16),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_79),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_149),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_92),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_218),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_40),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_163),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_88),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_13),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_128),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_71),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_51),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_90),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_89),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_222),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_205),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_146),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_210),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_171),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_53),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_27),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_83),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_90),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_17),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_34),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_54),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_138),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_91),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_43),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_135),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_30),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_77),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_81),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_206),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_61),
.Y(n_395)
);

BUFx2_ASAP7_75t_SL g396 ( 
.A(n_68),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_27),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_39),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_3),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_187),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_24),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_104),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_241),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_173),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_172),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_162),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_136),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_148),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_175),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_0),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_19),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_230),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_139),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_216),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_76),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_58),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_127),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_92),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_107),
.Y(n_419)
);

BUFx5_ASAP7_75t_L g420 ( 
.A(n_67),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_74),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_104),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_28),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_82),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_60),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_102),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_9),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_63),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_63),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_59),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_186),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_94),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_20),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_140),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_217),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_107),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_72),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_73),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_7),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_12),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_239),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_34),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_95),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_193),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_157),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_178),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_20),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_190),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_5),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_70),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_155),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_152),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_237),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_240),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_39),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_25),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_98),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_207),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_133),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_238),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_8),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_71),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_82),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_167),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_22),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_113),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_108),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_200),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_21),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_66),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_134),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_64),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_56),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_0),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_321),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_420),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_243),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_251),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_420),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_324),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_420),
.Y(n_481)
);

INVxp33_ASAP7_75t_SL g482 ( 
.A(n_272),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_355),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_420),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_420),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_420),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_420),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_290),
.B(n_1),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_413),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_R g491 ( 
.A(n_340),
.B(n_111),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_290),
.B(n_1),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_420),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_375),
.Y(n_494)
);

INVxp33_ASAP7_75t_SL g495 ( 
.A(n_447),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_356),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_420),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_320),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_320),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_320),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_320),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_R g502 ( 
.A(n_270),
.B(n_119),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_320),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_396),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_469),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_320),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_376),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_368),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_368),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_368),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_253),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_368),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_368),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_368),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_331),
.B(n_2),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_379),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g517 ( 
.A(n_331),
.B(n_2),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_408),
.B(n_6),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_265),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_342),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_467),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_394),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_266),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_269),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_281),
.Y(n_525)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_408),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_434),
.B(n_6),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_400),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_287),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_293),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_342),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_295),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_326),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_342),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_364),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_299),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_434),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_326),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_304),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_364),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_248),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_364),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_312),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_242),
.B(n_7),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_344),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_318),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_381),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_381),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_396),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_R g550 ( 
.A(n_319),
.B(n_327),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_381),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_242),
.B(n_8),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_391),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_344),
.B(n_9),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_391),
.B(n_10),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_391),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_421),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_244),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_L g559 ( 
.A(n_421),
.B(n_11),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_421),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_455),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_455),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_356),
.B(n_11),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_282),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_330),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_455),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_337),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_356),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_422),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_339),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_350),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_245),
.B(n_12),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_R g573 ( 
.A(n_367),
.B(n_120),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_422),
.Y(n_574)
);

NOR2xp67_ASAP7_75t_L g575 ( 
.A(n_470),
.B(n_15),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_370),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_422),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_440),
.B(n_15),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_390),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_404),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_344),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_405),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_406),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_260),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_244),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_414),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_431),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_245),
.B(n_18),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_440),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_441),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_R g591 ( 
.A(n_444),
.B(n_125),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_282),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_440),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_347),
.Y(n_594)
);

INVxp33_ASAP7_75t_L g595 ( 
.A(n_246),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_246),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_451),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_452),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_453),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_250),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_454),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_458),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_252),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_250),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_514),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_477),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_498),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_498),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_478),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_511),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_475),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_519),
.B(n_347),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_499),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_480),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_487),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_499),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_500),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_485),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_R g620 ( 
.A(n_543),
.B(n_460),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_500),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_523),
.B(n_347),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_501),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_R g624 ( 
.A(n_482),
.B(n_262),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_501),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_545),
.B(n_363),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_524),
.B(n_363),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_485),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_563),
.B(n_363),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_525),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_603),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_503),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_503),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_506),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_506),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_529),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_533),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_563),
.B(n_308),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_508),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_541),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_508),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_509),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_530),
.B(n_468),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_526),
.B(n_537),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_509),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_532),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_584),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_510),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_L g649 ( 
.A(n_491),
.B(n_264),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_510),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_512),
.Y(n_651)
);

AND3x2_ASAP7_75t_L g652 ( 
.A(n_489),
.B(n_518),
.C(n_492),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_505),
.B(n_296),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_483),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_536),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_512),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_539),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_513),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_567),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_513),
.Y(n_660)
);

BUFx8_ASAP7_75t_L g661 ( 
.A(n_496),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_570),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_594),
.B(n_255),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_560),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_494),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_560),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_476),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_496),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_571),
.B(n_308),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_579),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_495),
.A2(n_261),
.B1(n_317),
.B2(n_286),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_476),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_596),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_479),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_580),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_582),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_479),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_507),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_R g679 ( 
.A(n_546),
.B(n_273),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_481),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_596),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_600),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_600),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_583),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_604),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_604),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_516),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_481),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_484),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_484),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_586),
.Y(n_691)
);

BUFx8_ASAP7_75t_L g692 ( 
.A(n_578),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_486),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_522),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_587),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_486),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_599),
.B(n_602),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_488),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_550),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_538),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_488),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_493),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_565),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_620),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_638),
.A2(n_663),
.B1(n_629),
.B2(n_626),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_688),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_629),
.B(n_578),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_699),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_688),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_689),
.Y(n_710)
);

BUFx8_ASAP7_75t_SL g711 ( 
.A(n_611),
.Y(n_711)
);

INVxp33_ASAP7_75t_L g712 ( 
.A(n_631),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_606),
.B(n_505),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_628),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_664),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_664),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_609),
.B(n_564),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_672),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_689),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_669),
.B(n_490),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_644),
.A2(n_576),
.B1(n_597),
.B2(n_590),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_672),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_701),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_701),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_702),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_702),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_626),
.B(n_581),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_667),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_629),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_629),
.B(n_493),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_672),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_664),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_667),
.Y(n_733)
);

CKINVDCx16_ASAP7_75t_R g734 ( 
.A(n_679),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_667),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_610),
.B(n_564),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_638),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_672),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_674),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_638),
.B(n_247),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_630),
.B(n_592),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_638),
.B(n_497),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_624),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_636),
.B(n_592),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_646),
.B(n_655),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_637),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_664),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_668),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_703),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_612),
.B(n_497),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_674),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_622),
.B(n_581),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_674),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_663),
.B(n_568),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_627),
.B(n_288),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_673),
.B(n_568),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_677),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_628),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_628),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_673),
.B(n_569),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_628),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_677),
.Y(n_762)
);

NOR3xp33_ASAP7_75t_L g763 ( 
.A(n_616),
.B(n_521),
.C(n_527),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_697),
.B(n_575),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_692),
.A2(n_552),
.B1(n_572),
.B2(n_544),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_643),
.B(n_598),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_677),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_652),
.B(n_601),
.Y(n_768)
);

AND2x2_ASAP7_75t_SL g769 ( 
.A(n_649),
.B(n_308),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_681),
.B(n_569),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_680),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_680),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_664),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_653),
.B(n_575),
.Y(n_774)
);

AND2x6_ASAP7_75t_L g775 ( 
.A(n_680),
.B(n_445),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_672),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_664),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_619),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_619),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_672),
.Y(n_780)
);

AND2x2_ASAP7_75t_SL g781 ( 
.A(n_690),
.B(n_445),
.Y(n_781)
);

INVx6_ASAP7_75t_L g782 ( 
.A(n_628),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_680),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_628),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_690),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_693),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_635),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_SL g788 ( 
.A(n_657),
.B(n_521),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_681),
.B(n_247),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_637),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_693),
.Y(n_791)
);

OA22x2_ASAP7_75t_L g792 ( 
.A1(n_682),
.A2(n_577),
.B1(n_589),
.B2(n_574),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_682),
.B(n_254),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_640),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_693),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_661),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_615),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_683),
.B(n_574),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_693),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_696),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_696),
.B(n_303),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_619),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_690),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_690),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_635),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_659),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_696),
.B(n_323),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_696),
.B(n_346),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_607),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_605),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_605),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_607),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_608),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_662),
.B(n_502),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_683),
.B(n_577),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_605),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_690),
.B(n_459),
.Y(n_817)
);

AND2x6_ASAP7_75t_L g818 ( 
.A(n_690),
.B(n_445),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_608),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_613),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_635),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_613),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_617),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_617),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_618),
.Y(n_825)
);

OAI21xp33_ASAP7_75t_SL g826 ( 
.A1(n_685),
.A2(n_588),
.B(n_554),
.Y(n_826)
);

INVx6_ASAP7_75t_L g827 ( 
.A(n_698),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_698),
.B(n_589),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_618),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_698),
.B(n_593),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_698),
.B(n_593),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_621),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_698),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_698),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_621),
.B(n_309),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_623),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_635),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_623),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_635),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_614),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_692),
.A2(n_559),
.B1(n_555),
.B2(n_517),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_635),
.Y(n_842)
);

BUFx10_ASAP7_75t_L g843 ( 
.A(n_670),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_614),
.Y(n_844)
);

INVx4_ASAP7_75t_SL g845 ( 
.A(n_650),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_625),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_647),
.A2(n_549),
.B1(n_504),
.B2(n_528),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_692),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_675),
.B(n_595),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_676),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_661),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_625),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_632),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_614),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_685),
.B(n_520),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_L g856 ( 
.A(n_661),
.B(n_585),
.C(n_558),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_700),
.B(n_474),
.Y(n_857)
);

BUFx10_ASAP7_75t_L g858 ( 
.A(n_684),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_686),
.B(n_254),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_632),
.B(n_267),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_650),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_634),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_633),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_634),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_654),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_665),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_686),
.B(n_520),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_737),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_849),
.B(n_691),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_706),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_L g871 ( 
.A(n_765),
.B(n_705),
.C(n_727),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_750),
.B(n_692),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_SL g873 ( 
.A(n_763),
.B(n_671),
.C(n_695),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_737),
.B(n_633),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_710),
.B(n_641),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_710),
.B(n_641),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_743),
.B(n_700),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_748),
.B(n_671),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_727),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_706),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_841),
.B(n_661),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_769),
.A2(n_464),
.B1(n_446),
.B2(n_267),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_755),
.B(n_678),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_725),
.B(n_648),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_725),
.B(n_648),
.Y(n_885)
);

AND2x6_ASAP7_75t_SL g886 ( 
.A(n_768),
.B(n_329),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_769),
.A2(n_464),
.B1(n_446),
.B2(n_268),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_707),
.B(n_660),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_707),
.B(n_660),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_720),
.B(n_573),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_766),
.B(n_591),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_707),
.B(n_650),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_826),
.A2(n_382),
.B(n_256),
.C(n_259),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_709),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_709),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_711),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_707),
.B(n_752),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_730),
.A2(n_742),
.B(n_817),
.Y(n_898)
);

O2A1O1Ixp5_ASAP7_75t_L g899 ( 
.A1(n_740),
.A2(n_464),
.B(n_446),
.C(n_271),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_719),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_719),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_729),
.B(n_268),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_723),
.B(n_650),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_704),
.B(n_296),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_723),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_724),
.B(n_650),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_724),
.B(n_650),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_726),
.B(n_656),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_726),
.B(n_656),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_781),
.B(n_656),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_712),
.B(n_748),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_809),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_704),
.B(n_296),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_809),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_SL g915 ( 
.A(n_734),
.B(n_687),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_812),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_781),
.B(n_656),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_781),
.B(n_656),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_814),
.B(n_694),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_754),
.B(n_296),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_769),
.A2(n_271),
.B1(n_280),
.B2(n_275),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_801),
.B(n_656),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_807),
.B(n_666),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_740),
.A2(n_729),
.B1(n_754),
.B2(n_789),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_812),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_813),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_772),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_808),
.B(n_666),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_794),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_740),
.B(n_275),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_740),
.B(n_280),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_754),
.B(n_291),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_813),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_819),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_819),
.B(n_291),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_794),
.B(n_734),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_756),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_848),
.B(n_435),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_772),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_756),
.B(n_770),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_820),
.B(n_298),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_749),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_820),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_822),
.B(n_298),
.Y(n_944)
);

OAI22xp33_ASAP7_75t_L g945 ( 
.A1(n_774),
.A2(n_517),
.B1(n_515),
.B2(n_302),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_848),
.B(n_847),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_822),
.Y(n_947)
);

NAND2x1p5_ASAP7_75t_L g948 ( 
.A(n_791),
.B(n_302),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_756),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_791),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_823),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_823),
.B(n_311),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_824),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_824),
.B(n_311),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_789),
.A2(n_338),
.B1(n_341),
.B2(n_332),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_774),
.B(n_329),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_825),
.B(n_332),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_770),
.A2(n_559),
.B1(n_555),
.B2(n_515),
.Y(n_958)
);

BUFx6f_ASAP7_75t_SL g959 ( 
.A(n_806),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_774),
.B(n_258),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_825),
.B(n_338),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_770),
.A2(n_402),
.B1(n_365),
.B2(n_378),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_718),
.B(n_341),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_789),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_775),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_829),
.B(n_365),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_829),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_788),
.B(n_435),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_832),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_832),
.B(n_378),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_836),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_836),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_838),
.B(n_387),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_838),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_785),
.Y(n_975)
);

INVxp67_ASAP7_75t_SL g976 ( 
.A(n_785),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_846),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_846),
.B(n_387),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_789),
.A2(n_407),
.B1(n_409),
.B2(n_403),
.Y(n_979)
);

NOR3x1_ASAP7_75t_L g980 ( 
.A(n_856),
.B(n_256),
.C(n_255),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_852),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_793),
.A2(n_859),
.B1(n_798),
.B2(n_815),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_852),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_853),
.B(n_403),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_806),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_793),
.A2(n_409),
.B1(n_412),
.B2(n_407),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_793),
.A2(n_417),
.B1(n_448),
.B2(n_412),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_853),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_863),
.B(n_417),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_793),
.A2(n_466),
.B1(n_471),
.B2(n_448),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_863),
.B(n_466),
.Y(n_991)
);

O2A1O1Ixp5_ASAP7_75t_L g992 ( 
.A1(n_771),
.A2(n_471),
.B(n_639),
.C(n_634),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_764),
.A2(n_279),
.B1(n_377),
.B2(n_249),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_764),
.B(n_259),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_774),
.B(n_289),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_760),
.B(n_531),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_859),
.A2(n_279),
.B1(n_377),
.B2(n_249),
.Y(n_997)
);

OR2x6_ASAP7_75t_L g998 ( 
.A(n_764),
.B(n_263),
.Y(n_998)
);

O2A1O1Ixp5_ASAP7_75t_L g999 ( 
.A1(n_771),
.A2(n_642),
.B(n_645),
.C(n_639),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_783),
.B(n_658),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_783),
.B(n_658),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_859),
.A2(n_279),
.B1(n_377),
.B2(n_249),
.Y(n_1002)
);

NOR2x1p5_ASAP7_75t_L g1003 ( 
.A(n_749),
.B(n_263),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_786),
.B(n_639),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_721),
.B(n_435),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_786),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_795),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_859),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_795),
.B(n_658),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_760),
.B(n_531),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_799),
.B(n_651),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_708),
.B(n_435),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_799),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_861),
.A2(n_645),
.B(n_642),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_708),
.B(n_249),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_800),
.B(n_642),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_714),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_764),
.B(n_336),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_775),
.A2(n_279),
.B1(n_377),
.B2(n_249),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_746),
.B(n_257),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_800),
.B(n_645),
.Y(n_1021)
);

AND2x6_ASAP7_75t_SL g1022 ( 
.A(n_857),
.B(n_278),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_759),
.B(n_651),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_713),
.B(n_357),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_714),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_798),
.B(n_534),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_717),
.B(n_736),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_790),
.Y(n_1028)
);

NOR2xp67_ASAP7_75t_L g1029 ( 
.A(n_828),
.B(n_651),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_855),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_708),
.B(n_249),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_759),
.B(n_279),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_759),
.B(n_279),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_865),
.Y(n_1034)
);

AND2x6_ASAP7_75t_SL g1035 ( 
.A(n_857),
.B(n_278),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_784),
.B(n_377),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_775),
.A2(n_377),
.B1(n_473),
.B2(n_292),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_815),
.B(n_534),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_784),
.B(n_535),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_855),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_792),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_741),
.Y(n_1042)
);

AND2x2_ASAP7_75t_SL g1043 ( 
.A(n_830),
.B(n_284),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_940),
.B(n_879),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_870),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_1028),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_SL g1047 ( 
.A(n_873),
.B(n_866),
.C(n_865),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1006),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1006),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_940),
.B(n_879),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1007),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_870),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1030),
.B(n_792),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_880),
.B(n_835),
.Y(n_1054)
);

INVx3_ASAP7_75t_SL g1055 ( 
.A(n_942),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_SL g1056 ( 
.A(n_1024),
.B(n_866),
.C(n_797),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1007),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1013),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_965),
.Y(n_1059)
);

BUFx12f_ASAP7_75t_L g1060 ( 
.A(n_1022),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_897),
.A2(n_722),
.B(n_718),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_1028),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1013),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_985),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1030),
.B(n_792),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_985),
.Y(n_1066)
);

NAND2x1_ASAP7_75t_L g1067 ( 
.A(n_975),
.B(n_827),
.Y(n_1067)
);

NAND3xp33_ASAP7_75t_L g1068 ( 
.A(n_911),
.B(n_744),
.C(n_745),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_937),
.B(n_867),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_965),
.B(n_718),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_929),
.Y(n_1071)
);

NAND2x1_ASAP7_75t_L g1072 ( 
.A(n_975),
.B(n_827),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_900),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_R g1074 ( 
.A(n_942),
.B(n_806),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_950),
.Y(n_1075)
);

INVx6_ASAP7_75t_L g1076 ( 
.A(n_950),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_900),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_905),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_927),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_950),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_SL g1081 ( 
.A(n_956),
.B(n_276),
.C(n_274),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_869),
.B(n_843),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1040),
.B(n_867),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_937),
.B(n_843),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_880),
.B(n_831),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_927),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_905),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_916),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_L g1089 ( 
.A(n_921),
.B(n_775),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_916),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_894),
.B(n_728),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_925),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_927),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_1020),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_939),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_1020),
.Y(n_1096)
);

BUFx8_ASAP7_75t_SL g1097 ( 
.A(n_896),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_896),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_925),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_894),
.B(n_728),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_949),
.B(n_796),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_895),
.B(n_733),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_924),
.A2(n_857),
.B1(n_851),
.B2(n_796),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_871),
.A2(n_857),
.B1(n_775),
.B2(n_784),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_877),
.B(n_843),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_960),
.B(n_850),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_949),
.B(n_851),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_872),
.B(n_850),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_995),
.B(n_850),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_895),
.B(n_733),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_L g1111 ( 
.A(n_1018),
.B(n_860),
.C(n_283),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_878),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_943),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_943),
.Y(n_1114)
);

BUFx4_ASAP7_75t_SL g1115 ( 
.A(n_1022),
.Y(n_1115)
);

INVx5_ASAP7_75t_L g1116 ( 
.A(n_965),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_959),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_901),
.B(n_912),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_950),
.Y(n_1119)
);

BUFx12f_ASAP7_75t_L g1120 ( 
.A(n_1035),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_950),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_878),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_947),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1041),
.A2(n_775),
.B1(n_739),
.B2(n_751),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1041),
.B(n_715),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_947),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_901),
.B(n_735),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_893),
.A2(n_735),
.B(n_751),
.C(n_739),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_951),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_L g1130 ( 
.A(n_962),
.B(n_285),
.C(n_277),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_912),
.B(n_753),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_994),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_883),
.B(n_1042),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_R g1134 ( 
.A(n_915),
.B(n_858),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_945),
.B(n_858),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_891),
.B(n_1027),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_868),
.B(n_715),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_868),
.B(n_716),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_965),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_914),
.B(n_926),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_914),
.B(n_753),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_939),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_994),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_982),
.B(n_858),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1040),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_939),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_951),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_953),
.Y(n_1148)
);

NAND2x1p5_ASAP7_75t_L g1149 ( 
.A(n_965),
.B(n_722),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_902),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_953),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_996),
.B(n_757),
.Y(n_1152)
);

AND2x6_ASAP7_75t_L g1153 ( 
.A(n_982),
.B(n_716),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_969),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_969),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_1017),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_926),
.B(n_757),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_933),
.B(n_762),
.Y(n_1158)
);

NOR3xp33_ASAP7_75t_SL g1159 ( 
.A(n_1005),
.B(n_297),
.C(n_294),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_972),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_996),
.B(n_1010),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_R g1162 ( 
.A(n_959),
.B(n_775),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_933),
.B(n_762),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_972),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_934),
.B(n_767),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_902),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_959),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_974),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_890),
.B(n_785),
.Y(n_1169)
);

CKINVDCx8_ASAP7_75t_R g1170 ( 
.A(n_886),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_974),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_SL g1172 ( 
.A(n_946),
.B(n_305),
.C(n_301),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1010),
.B(n_767),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_902),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1003),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_975),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1026),
.B(n_1043),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1003),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_934),
.B(n_778),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_981),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1043),
.A2(n_818),
.B1(n_779),
.B2(n_802),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_964),
.A2(n_1008),
.B1(n_1043),
.B2(n_889),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_964),
.B(n_732),
.Y(n_1183)
);

BUFx4f_ASAP7_75t_L g1184 ( 
.A(n_948),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_994),
.B(n_827),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1008),
.B(n_732),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_981),
.Y(n_1187)
);

AOI211xp5_ASAP7_75t_L g1188 ( 
.A1(n_936),
.A2(n_372),
.B(n_385),
.C(n_257),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_967),
.Y(n_1189)
);

INVx5_ASAP7_75t_L g1190 ( 
.A(n_1017),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_962),
.A2(n_352),
.B1(n_316),
.B2(n_300),
.C(n_292),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_886),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1038),
.B(n_785),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_967),
.B(n_778),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1017),
.Y(n_1195)
);

NOR3xp33_ASAP7_75t_SL g1196 ( 
.A(n_904),
.B(n_307),
.C(n_306),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1038),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1038),
.B(n_747),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_971),
.Y(n_1199)
);

NOR2x1p5_ASAP7_75t_L g1200 ( 
.A(n_932),
.B(n_310),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_971),
.B(n_779),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_994),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_SL g1203 ( 
.A(n_913),
.B(n_314),
.C(n_313),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1026),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_977),
.B(n_802),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_977),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1034),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1025),
.Y(n_1208)
);

NOR3xp33_ASAP7_75t_SL g1209 ( 
.A(n_968),
.B(n_322),
.C(n_315),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_998),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_983),
.Y(n_1211)
);

NAND2xp33_ASAP7_75t_SL g1212 ( 
.A(n_882),
.B(n_785),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_998),
.B(n_325),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_983),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_988),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_988),
.B(n_787),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_999),
.Y(n_1217)
);

BUFx10_ASAP7_75t_L g1218 ( 
.A(n_919),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_998),
.B(n_747),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_887),
.B(n_787),
.Y(n_1220)
);

AND2x4_ASAP7_75t_SL g1221 ( 
.A(n_998),
.B(n_282),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_923),
.B(n_787),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_888),
.B(n_773),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_R g1224 ( 
.A(n_1035),
.B(n_805),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_928),
.B(n_805),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1025),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_958),
.B(n_804),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_948),
.Y(n_1228)
);

OR2x2_ASAP7_75t_SL g1229 ( 
.A(n_881),
.B(n_284),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_874),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1039),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1025),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1000),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_875),
.Y(n_1234)
);

NOR3xp33_ASAP7_75t_SL g1235 ( 
.A(n_1012),
.B(n_335),
.C(n_334),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_892),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_876),
.B(n_805),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1001),
.Y(n_1238)
);

CKINVDCx6p67_ASAP7_75t_R g1239 ( 
.A(n_1055),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1136),
.A2(n_910),
.B1(n_918),
.B2(n_917),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1217),
.A2(n_1061),
.B(n_1236),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1080),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1059),
.A2(n_898),
.B(n_976),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1161),
.B(n_884),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1217),
.A2(n_1236),
.B(n_1072),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1059),
.A2(n_922),
.B(n_731),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1161),
.B(n_1234),
.Y(n_1247)
);

OA22x2_ASAP7_75t_L g1248 ( 
.A1(n_1112),
.A2(n_990),
.B1(n_958),
.B2(n_920),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1236),
.A2(n_1033),
.B(n_1032),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1133),
.B(n_938),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1176),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1220),
.A2(n_906),
.B(n_903),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1062),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1177),
.A2(n_1002),
.B1(n_997),
.B2(n_963),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1230),
.B(n_885),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1067),
.A2(n_1036),
.B(n_992),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1176),
.Y(n_1257)
);

O2A1O1Ixp5_ASAP7_75t_L g1258 ( 
.A1(n_1169),
.A2(n_1031),
.B(n_1015),
.C(n_1227),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1182),
.A2(n_1089),
.B(n_1104),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1067),
.A2(n_1072),
.B(n_1118),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1204),
.B(n_935),
.Y(n_1261)
);

NAND3x1_ASAP7_75t_L g1262 ( 
.A(n_1082),
.B(n_990),
.C(n_316),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1176),
.A2(n_963),
.B(n_993),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1177),
.B(n_980),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1140),
.A2(n_908),
.B(n_907),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1054),
.B(n_1083),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1083),
.B(n_941),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1152),
.B(n_944),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1214),
.A2(n_963),
.B1(n_1019),
.B2(n_948),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1176),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1176),
.A2(n_931),
.B(n_930),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1152),
.B(n_952),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1089),
.A2(n_909),
.B(n_1029),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1228),
.A2(n_731),
.B(n_722),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1125),
.A2(n_1029),
.B(n_899),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1173),
.B(n_954),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1206),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1096),
.B(n_957),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1106),
.B(n_1105),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1184),
.B(n_961),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1097),
.Y(n_1281)
);

AOI31xp67_ASAP7_75t_L g1282 ( 
.A1(n_1206),
.A2(n_970),
.A3(n_973),
.B(n_966),
.Y(n_1282)
);

NAND3x1_ASAP7_75t_L g1283 ( 
.A(n_1191),
.B(n_328),
.C(n_300),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1053),
.B(n_1065),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1057),
.Y(n_1285)
);

AOI21xp33_ASAP7_75t_L g1286 ( 
.A1(n_1094),
.A2(n_984),
.B(n_978),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1046),
.B(n_989),
.Y(n_1287)
);

AO32x2_ASAP7_75t_L g1288 ( 
.A1(n_1228),
.A2(n_1166),
.A3(n_1103),
.B1(n_1121),
.B2(n_1075),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1059),
.A2(n_738),
.B(n_731),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1128),
.A2(n_1009),
.B(n_1004),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1097),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_SL g1292 ( 
.A1(n_1211),
.A2(n_1215),
.B(n_1166),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1214),
.A2(n_955),
.B1(n_986),
.B2(n_979),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1216),
.A2(n_1016),
.B(n_1011),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1091),
.A2(n_1102),
.B(n_1100),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1062),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1057),
.Y(n_1297)
);

BUFx8_ASAP7_75t_L g1298 ( 
.A(n_1096),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1080),
.B(n_738),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1173),
.B(n_991),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1197),
.B(n_980),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1110),
.A2(n_1021),
.B(n_1023),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1058),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1071),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1127),
.A2(n_1014),
.B(n_777),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1122),
.B(n_343),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1059),
.A2(n_776),
.B(n_738),
.Y(n_1307)
);

BUFx4f_ASAP7_75t_SL g1308 ( 
.A(n_1055),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1184),
.B(n_987),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1233),
.B(n_1037),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1058),
.A2(n_777),
.B(n_773),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1131),
.A2(n_837),
.B(n_821),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1059),
.A2(n_780),
.B(n_776),
.Y(n_1313)
);

AO21x1_ASAP7_75t_L g1314 ( 
.A1(n_1212),
.A2(n_333),
.B(n_328),
.Y(n_1314)
);

AND3x4_ASAP7_75t_L g1315 ( 
.A(n_1047),
.B(n_353),
.C(n_282),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1141),
.A2(n_1158),
.B(n_1157),
.Y(n_1316)
);

AO32x2_ASAP7_75t_L g1317 ( 
.A1(n_1075),
.A2(n_776),
.A3(n_780),
.B1(n_803),
.B2(n_359),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1163),
.A2(n_837),
.B(n_821),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1116),
.A2(n_803),
.B(n_780),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1233),
.B(n_862),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1238),
.B(n_862),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1053),
.A2(n_428),
.B(n_352),
.C(n_354),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1080),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1211),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1080),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1070),
.A2(n_1149),
.B(n_1119),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_L g1327 ( 
.A(n_1188),
.B(n_348),
.C(n_345),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1080),
.Y(n_1328)
);

AO32x2_ASAP7_75t_L g1329 ( 
.A1(n_1121),
.A2(n_803),
.A3(n_354),
.B1(n_359),
.B2(n_333),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1215),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1071),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1064),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1122),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1238),
.B(n_864),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1184),
.B(n_804),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1165),
.A2(n_837),
.B(n_821),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1116),
.A2(n_758),
.B(n_714),
.Y(n_1337)
);

AOI221xp5_ASAP7_75t_L g1338 ( 
.A1(n_1130),
.A2(n_349),
.B1(n_351),
.B2(n_358),
.C(n_366),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1116),
.A2(n_758),
.B(n_714),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1179),
.A2(n_839),
.B(n_864),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1189),
.A2(n_782),
.B1(n_827),
.B2(n_761),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1125),
.A2(n_839),
.B(n_811),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1045),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1194),
.A2(n_1205),
.B(n_1201),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1199),
.A2(n_782),
.B1(n_758),
.B2(n_761),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1065),
.A2(n_461),
.B(n_360),
.C(n_361),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1207),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1056),
.B(n_369),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_SL g1349 ( 
.A1(n_1195),
.A2(n_361),
.B(n_360),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1125),
.B(n_810),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1087),
.A2(n_811),
.B(n_810),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1139),
.Y(n_1352)
);

AO32x2_ASAP7_75t_L g1353 ( 
.A1(n_1195),
.A2(n_1229),
.A3(n_1153),
.B1(n_1172),
.B2(n_1212),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1150),
.A2(n_782),
.B1(n_758),
.B2(n_761),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1074),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1079),
.A2(n_839),
.B(n_816),
.Y(n_1356)
);

AOI211x1_ASAP7_75t_L g1357 ( 
.A1(n_1048),
.A2(n_429),
.B(n_428),
.C(n_426),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1079),
.A2(n_840),
.B(n_816),
.Y(n_1358)
);

NOR2xp67_ASAP7_75t_L g1359 ( 
.A(n_1068),
.B(n_126),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1069),
.B(n_840),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1087),
.Y(n_1361)
);

AOI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1099),
.A2(n_854),
.B(n_844),
.Y(n_1362)
);

AOI221xp5_ASAP7_75t_L g1363 ( 
.A1(n_1145),
.A2(n_437),
.B1(n_392),
.B2(n_371),
.C(n_373),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1119),
.B(n_804),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1079),
.A2(n_854),
.B(n_844),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1069),
.B(n_714),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1116),
.A2(n_761),
.B(n_758),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1086),
.A2(n_540),
.B(n_535),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1044),
.B(n_804),
.Y(n_1369)
);

AO21x1_ASAP7_75t_L g1370 ( 
.A1(n_1099),
.A2(n_386),
.B(n_362),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1064),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1076),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1086),
.A2(n_1095),
.B(n_1093),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1237),
.A2(n_542),
.B(n_540),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1126),
.A2(n_547),
.B(n_542),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1086),
.A2(n_1095),
.B(n_1093),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1207),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1223),
.A2(n_818),
.B(n_386),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1222),
.A2(n_1225),
.B(n_1085),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1093),
.A2(n_1142),
.B(n_1095),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1045),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1175),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1116),
.A2(n_761),
.B(n_804),
.Y(n_1383)
);

NAND2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1119),
.B(n_833),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1142),
.A2(n_548),
.B(n_547),
.Y(n_1385)
);

NOR2x1_ASAP7_75t_L g1386 ( 
.A(n_1066),
.B(n_362),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1052),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1069),
.B(n_548),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1223),
.A2(n_818),
.B(n_398),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1044),
.B(n_782),
.Y(n_1390)
);

AO21x1_ASAP7_75t_L g1391 ( 
.A1(n_1126),
.A2(n_398),
.B(n_389),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1142),
.A2(n_553),
.B(n_551),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1070),
.A2(n_834),
.B(n_833),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1052),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1119),
.B(n_833),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1044),
.B(n_833),
.Y(n_1396)
);

AO21x1_ASAP7_75t_L g1397 ( 
.A1(n_1147),
.A2(n_1160),
.B(n_1151),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1139),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1049),
.A2(n_1051),
.B(n_1063),
.C(n_1147),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1050),
.B(n_833),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1050),
.B(n_834),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1139),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1050),
.B(n_834),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1146),
.A2(n_553),
.B(n_551),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1146),
.A2(n_1092),
.B(n_1088),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1146),
.A2(n_557),
.B(n_556),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_SL g1407 ( 
.A1(n_1195),
.A2(n_399),
.B(n_389),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1285),
.Y(n_1408)
);

AOI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1397),
.A2(n_1160),
.B(n_1151),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1245),
.A2(n_1092),
.B(n_1088),
.Y(n_1410)
);

AO31x2_ASAP7_75t_L g1411 ( 
.A1(n_1314),
.A2(n_1164),
.A3(n_1129),
.B(n_1155),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1245),
.A2(n_1129),
.B(n_1114),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1279),
.A2(n_1174),
.B1(n_1150),
.B2(n_1197),
.Y(n_1413)
);

CKINVDCx9p33_ASAP7_75t_R g1414 ( 
.A(n_1347),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1297),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1303),
.Y(n_1416)
);

AO21x2_ASAP7_75t_L g1417 ( 
.A1(n_1259),
.A2(n_1318),
.B(n_1312),
.Y(n_1417)
);

AOI222xp33_ASAP7_75t_L g1418 ( 
.A1(n_1250),
.A2(n_1109),
.B1(n_1135),
.B2(n_1060),
.C1(n_1120),
.C2(n_1221),
.Y(n_1418)
);

AO21x1_ASAP7_75t_L g1419 ( 
.A1(n_1240),
.A2(n_1164),
.B(n_1108),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1266),
.B(n_1247),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1405),
.A2(n_1155),
.B(n_1114),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1312),
.A2(n_1144),
.B(n_1077),
.Y(n_1422)
);

AO21x2_ASAP7_75t_L g1423 ( 
.A1(n_1318),
.A2(n_1078),
.B(n_1073),
.Y(n_1423)
);

AO31x2_ASAP7_75t_L g1424 ( 
.A1(n_1314),
.A2(n_1171),
.A3(n_1113),
.B(n_1123),
.Y(n_1424)
);

NAND2xp33_ASAP7_75t_R g1425 ( 
.A(n_1355),
.B(n_1134),
.Y(n_1425)
);

INVx3_ASAP7_75t_SL g1426 ( 
.A(n_1239),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_SL g1427 ( 
.A1(n_1397),
.A2(n_1171),
.B(n_1148),
.Y(n_1427)
);

NOR2xp67_ASAP7_75t_L g1428 ( 
.A(n_1355),
.B(n_1111),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1284),
.B(n_1174),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1405),
.A2(n_1154),
.B(n_1090),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_SL g1431 ( 
.A1(n_1292),
.A2(n_1180),
.B(n_1168),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1277),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1336),
.A2(n_1187),
.B(n_1231),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1336),
.A2(n_1231),
.B(n_1208),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1340),
.A2(n_1208),
.B(n_1156),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_SL g1436 ( 
.A1(n_1309),
.A2(n_1193),
.B(n_1084),
.C(n_1178),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1324),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1340),
.A2(n_1208),
.B(n_1156),
.Y(n_1438)
);

NOR2xp67_ASAP7_75t_L g1439 ( 
.A(n_1333),
.B(n_1117),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1296),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1258),
.A2(n_1244),
.B(n_1254),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_SL g1442 ( 
.A1(n_1309),
.A2(n_1232),
.B(n_1213),
.C(n_1156),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1255),
.B(n_1218),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1249),
.A2(n_1181),
.B(n_1223),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1241),
.A2(n_1232),
.B(n_1149),
.Y(n_1445)
);

INVxp67_ASAP7_75t_SL g1446 ( 
.A(n_1257),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1330),
.Y(n_1447)
);

NAND2xp33_ASAP7_75t_R g1448 ( 
.A(n_1281),
.B(n_1162),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1326),
.A2(n_1149),
.B(n_1070),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1348),
.B(n_1159),
.C(n_1209),
.Y(n_1450)
);

CKINVDCx6p67_ASAP7_75t_R g1451 ( 
.A(n_1239),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1326),
.A2(n_1139),
.B(n_1190),
.Y(n_1452)
);

AO21x2_ASAP7_75t_L g1453 ( 
.A1(n_1249),
.A2(n_1138),
.B(n_1137),
.Y(n_1453)
);

AOI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1280),
.A2(n_1241),
.B(n_1351),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1268),
.B(n_1229),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1304),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1273),
.A2(n_1138),
.B(n_1137),
.Y(n_1457)
);

OAI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1377),
.A2(n_1167),
.B1(n_1117),
.B2(n_1213),
.Y(n_1458)
);

O2A1O1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1286),
.A2(n_1081),
.B(n_1235),
.C(n_1196),
.Y(n_1459)
);

OR2x6_ASAP7_75t_L g1460 ( 
.A(n_1263),
.B(n_1185),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1272),
.A2(n_1185),
.B1(n_1107),
.B2(n_1101),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1358),
.A2(n_1124),
.B(n_1200),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1352),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1358),
.A2(n_557),
.B(n_556),
.Y(n_1464)
);

OAI222xp33_ASAP7_75t_L g1465 ( 
.A1(n_1248),
.A2(n_1170),
.B1(n_1185),
.B2(n_1132),
.C1(n_1143),
.C2(n_1210),
.Y(n_1465)
);

NAND3x1_ASAP7_75t_L g1466 ( 
.A(n_1264),
.B(n_401),
.C(n_399),
.Y(n_1466)
);

AO21x2_ASAP7_75t_L g1467 ( 
.A1(n_1374),
.A2(n_1138),
.B(n_1137),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1331),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1365),
.A2(n_562),
.B(n_561),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1284),
.B(n_1218),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1327),
.B(n_1203),
.C(n_1192),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1361),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1343),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1265),
.A2(n_562),
.B(n_561),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1296),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1365),
.A2(n_566),
.B(n_1153),
.Y(n_1476)
);

AO21x1_ASAP7_75t_L g1477 ( 
.A1(n_1280),
.A2(n_1335),
.B(n_1269),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1343),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1248),
.A2(n_1264),
.B1(n_1301),
.B2(n_1143),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1332),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1287),
.B(n_1218),
.Y(n_1481)
);

BUFx4f_ASAP7_75t_SL g1482 ( 
.A(n_1298),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1381),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1388),
.B(n_1350),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1381),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_SL g1486 ( 
.A1(n_1370),
.A2(n_1153),
.B(n_410),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1251),
.Y(n_1487)
);

INVx4_ASAP7_75t_L g1488 ( 
.A(n_1242),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1253),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1356),
.A2(n_566),
.B(n_1153),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1301),
.B(n_1219),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1356),
.A2(n_1260),
.B(n_1368),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1260),
.A2(n_1153),
.B(n_410),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1387),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1387),
.Y(n_1495)
);

AO21x2_ASAP7_75t_L g1496 ( 
.A1(n_1374),
.A2(n_1219),
.B(n_1186),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1368),
.A2(n_1153),
.B(n_426),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1306),
.B(n_1132),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1382),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1265),
.A2(n_1186),
.B(n_1183),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1394),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1359),
.A2(n_1221),
.B(n_1107),
.C(n_1101),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1394),
.Y(n_1503)
);

AOI222xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1315),
.A2(n_430),
.B1(n_401),
.B2(n_429),
.C1(n_473),
.C2(n_461),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1350),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1375),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1375),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1320),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1385),
.A2(n_432),
.B(n_430),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1332),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1243),
.A2(n_1139),
.B(n_1190),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1322),
.A2(n_1210),
.B(n_1202),
.C(n_1107),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1388),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1276),
.A2(n_1185),
.B1(n_1101),
.B2(n_1076),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1278),
.B(n_1202),
.Y(n_1515)
);

CKINVDCx6p67_ASAP7_75t_R g1516 ( 
.A(n_1371),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1375),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1399),
.Y(n_1518)
);

AO21x1_ASAP7_75t_L g1519 ( 
.A1(n_1335),
.A2(n_1186),
.B(n_1183),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1385),
.A2(n_432),
.B(n_1190),
.Y(n_1520)
);

AO21x1_ASAP7_75t_L g1521 ( 
.A1(n_1252),
.A2(n_1183),
.B(n_1198),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1300),
.B(n_1198),
.Y(n_1522)
);

INVx1_ASAP7_75t_SL g1523 ( 
.A(n_1308),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1392),
.A2(n_1190),
.B(n_1119),
.Y(n_1524)
);

AO21x2_ASAP7_75t_L g1525 ( 
.A1(n_1374),
.A2(n_1219),
.B(n_1198),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1321),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1267),
.B(n_1066),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1338),
.B(n_1192),
.C(n_1170),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1278),
.B(n_1098),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1362),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1316),
.A2(n_438),
.B(n_380),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1392),
.A2(n_1190),
.B(n_1076),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1334),
.Y(n_1533)
);

AO21x2_ASAP7_75t_L g1534 ( 
.A1(n_1275),
.A2(n_1224),
.B(n_1076),
.Y(n_1534)
);

AOI22x1_ASAP7_75t_L g1535 ( 
.A1(n_1349),
.A2(n_1167),
.B1(n_834),
.B2(n_842),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1404),
.A2(n_1226),
.B(n_818),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1404),
.A2(n_1226),
.B(n_818),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1242),
.Y(n_1538)
);

NAND2x1p5_ASAP7_75t_L g1539 ( 
.A(n_1251),
.B(n_834),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1406),
.A2(n_818),
.B(n_845),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1251),
.B(n_842),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1399),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1352),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1301),
.A2(n_1120),
.B1(n_1060),
.B2(n_1098),
.Y(n_1544)
);

CKINVDCx6p67_ASAP7_75t_R g1545 ( 
.A(n_1371),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1360),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1261),
.B(n_374),
.Y(n_1547)
);

BUFx2_ASAP7_75t_R g1548 ( 
.A(n_1281),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1316),
.A2(n_384),
.B(n_388),
.Y(n_1549)
);

AO221x2_ASAP7_75t_L g1550 ( 
.A1(n_1293),
.A2(n_353),
.B1(n_383),
.B2(n_24),
.C(n_25),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1262),
.A2(n_433),
.B1(n_393),
.B2(n_395),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1406),
.A2(n_818),
.B(n_845),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1373),
.A2(n_1380),
.B(n_1376),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1298),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1386),
.B(n_397),
.Y(n_1555)
);

OAI22x1_ASAP7_75t_L g1556 ( 
.A1(n_1315),
.A2(n_436),
.B1(n_472),
.B2(n_465),
.Y(n_1556)
);

AOI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1290),
.A2(n_845),
.B(n_842),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1366),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1311),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1298),
.A2(n_353),
.B1(n_383),
.B2(n_427),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1373),
.A2(n_845),
.B(n_842),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1311),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1263),
.A2(n_842),
.B(n_142),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1311),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1242),
.Y(n_1565)
);

NOR2xp67_ASAP7_75t_L g1566 ( 
.A(n_1291),
.B(n_144),
.Y(n_1566)
);

AOI21xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1291),
.A2(n_439),
.B(n_463),
.Y(n_1567)
);

BUFx2_ASAP7_75t_R g1568 ( 
.A(n_1369),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1376),
.A2(n_234),
.B(n_231),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1380),
.Y(n_1570)
);

OR2x6_ASAP7_75t_L g1571 ( 
.A(n_1271),
.B(n_1115),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1352),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1379),
.B(n_411),
.Y(n_1573)
);

AOI21xp33_ASAP7_75t_L g1574 ( 
.A1(n_1262),
.A2(n_462),
.B(n_457),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1271),
.A2(n_209),
.B(n_156),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1379),
.B(n_456),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1310),
.A2(n_450),
.B(n_443),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1322),
.B(n_353),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1270),
.B(n_145),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1390),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1305),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1256),
.A2(n_228),
.B(n_225),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1398),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1369),
.A2(n_383),
.B1(n_425),
.B2(n_424),
.Y(n_1584)
);

AO21x2_ASAP7_75t_L g1585 ( 
.A1(n_1379),
.A2(n_223),
.B(n_219),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1396),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1295),
.B(n_415),
.Y(n_1587)
);

BUFx5_ASAP7_75t_L g1588 ( 
.A(n_1282),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1400),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1407),
.A2(n_383),
.B1(n_423),
.B2(n_419),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1283),
.A2(n_442),
.B1(n_418),
.B2(n_416),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1242),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_SL g1593 ( 
.A1(n_1550),
.A2(n_1378),
.B1(n_1389),
.B2(n_1283),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1484),
.B(n_1346),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1548),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1491),
.B(n_1270),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1408),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1449),
.A2(n_1295),
.B(n_1274),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1488),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1550),
.A2(n_1370),
.B1(n_1391),
.B2(n_1363),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1480),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1457),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1452),
.A2(n_1295),
.B(n_1274),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1408),
.Y(n_1604)
);

NOR3xp33_ASAP7_75t_SL g1605 ( 
.A(n_1450),
.B(n_1346),
.C(n_1354),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1498),
.A2(n_1401),
.B1(n_1403),
.B2(n_1270),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1415),
.Y(n_1607)
);

AO221x2_ASAP7_75t_L g1608 ( 
.A1(n_1465),
.A2(n_1353),
.B1(n_1329),
.B2(n_1288),
.C(n_1391),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1425),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1504),
.A2(n_1372),
.B1(n_1323),
.B2(n_1341),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1443),
.A2(n_1323),
.B1(n_1357),
.B2(n_1372),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1484),
.B(n_1353),
.Y(n_1612)
);

NAND3xp33_ASAP7_75t_SL g1613 ( 
.A(n_1418),
.B(n_1342),
.C(n_1246),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1455),
.A2(n_1323),
.B1(n_1299),
.B2(n_1328),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1420),
.B(n_1344),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1455),
.A2(n_1325),
.B1(n_1328),
.B2(n_1353),
.Y(n_1616)
);

A2O1A1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1512),
.A2(n_1344),
.B(n_1290),
.C(n_1302),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1538),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1528),
.A2(n_1345),
.B1(n_1398),
.B2(n_1402),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1479),
.A2(n_1299),
.B1(n_1328),
.B2(n_1325),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1481),
.A2(n_1328),
.B1(n_1325),
.B2(n_1395),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1457),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1491),
.B(n_1398),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1502),
.A2(n_1325),
.B(n_1395),
.Y(n_1624)
);

OR2x6_ASAP7_75t_SL g1625 ( 
.A(n_1471),
.B(n_1529),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1429),
.B(n_1353),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1529),
.B(n_1364),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1491),
.B(n_1402),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1473),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1475),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_SL g1631 ( 
.A(n_1560),
.B(n_1384),
.C(n_1364),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1429),
.B(n_1288),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1473),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1550),
.A2(n_1402),
.B1(n_1302),
.B2(n_1294),
.Y(n_1634)
);

AOI21xp33_ASAP7_75t_L g1635 ( 
.A1(n_1577),
.A2(n_1294),
.B(n_1305),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1574),
.A2(n_1393),
.B1(n_1383),
.B2(n_1339),
.C(n_1367),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1489),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1550),
.A2(n_1256),
.B1(n_1384),
.B2(n_1288),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1513),
.B(n_21),
.Y(n_1639)
);

AOI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1556),
.A2(n_1337),
.B1(n_1319),
.B2(n_1313),
.C(n_1307),
.Y(n_1640)
);

OAI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1470),
.A2(n_1551),
.B1(n_1527),
.B2(n_1571),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1416),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1573),
.A2(n_1289),
.B(n_1288),
.Y(n_1643)
);

BUFx2_ASAP7_75t_SL g1644 ( 
.A(n_1440),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1472),
.Y(n_1645)
);

AND2x2_ASAP7_75t_SL g1646 ( 
.A(n_1578),
.B(n_1317),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1437),
.Y(n_1647)
);

NOR3xp33_ASAP7_75t_SL g1648 ( 
.A(n_1458),
.B(n_1448),
.C(n_1459),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1432),
.Y(n_1649)
);

NAND2xp33_ASAP7_75t_R g1650 ( 
.A(n_1460),
.B(n_1317),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1429),
.B(n_1329),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1556),
.A2(n_1329),
.B1(n_26),
.B2(n_29),
.C(n_31),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1488),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1488),
.Y(n_1654)
);

NAND2xp33_ASAP7_75t_SL g1655 ( 
.A(n_1426),
.B(n_1317),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1538),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1515),
.B(n_1329),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1578),
.A2(n_22),
.B1(n_29),
.B2(n_31),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1456),
.B(n_1468),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1457),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1460),
.A2(n_1441),
.B(n_1511),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1460),
.A2(n_1317),
.B(n_214),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1580),
.B(n_35),
.Y(n_1663)
);

BUFx6f_ASAP7_75t_L g1664 ( 
.A(n_1538),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1499),
.Y(n_1665)
);

OAI22xp33_ASAP7_75t_SL g1666 ( 
.A1(n_1571),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1568),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_1667)
);

INVx6_ASAP7_75t_L g1668 ( 
.A(n_1440),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1480),
.Y(n_1669)
);

NAND2xp33_ASAP7_75t_SL g1670 ( 
.A(n_1426),
.B(n_41),
.Y(n_1670)
);

INVx4_ASAP7_75t_L g1671 ( 
.A(n_1516),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1475),
.B(n_213),
.Y(n_1672)
);

AOI21xp33_ASAP7_75t_L g1673 ( 
.A1(n_1576),
.A2(n_41),
.B(n_44),
.Y(n_1673)
);

AND2x2_ASAP7_75t_SL g1674 ( 
.A(n_1444),
.B(n_45),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1483),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1483),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1522),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1460),
.A2(n_212),
.B(n_208),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1461),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1482),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1451),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1505),
.B(n_50),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1447),
.Y(n_1683)
);

NAND2x1_ASAP7_75t_L g1684 ( 
.A(n_1431),
.B(n_197),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1446),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1538),
.Y(n_1686)
);

INVx4_ASAP7_75t_L g1687 ( 
.A(n_1516),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1544),
.A2(n_1571),
.B1(n_1555),
.B2(n_1584),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1510),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1439),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1495),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1522),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1525),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1571),
.A2(n_55),
.B1(n_57),
.B2(n_60),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_SL g1695 ( 
.A(n_1591),
.B(n_62),
.C(n_64),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1554),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1505),
.B(n_65),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1451),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1414),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1428),
.B(n_196),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1545),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1477),
.A2(n_68),
.B1(n_70),
.B2(n_73),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1477),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1538),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1546),
.B(n_77),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_SL g1706 ( 
.A(n_1567),
.B(n_79),
.C(n_85),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1587),
.A2(n_86),
.B(n_88),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1518),
.A2(n_91),
.B1(n_93),
.B2(n_96),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1492),
.A2(n_170),
.B(n_194),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1576),
.B(n_96),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1545),
.Y(n_1711)
);

NAND2x1_ASAP7_75t_L g1712 ( 
.A(n_1431),
.B(n_164),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1546),
.B(n_97),
.Y(n_1713)
);

OAI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1547),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_1714)
);

OAI222xp33_ASAP7_75t_L g1715 ( 
.A1(n_1413),
.A2(n_103),
.B1(n_105),
.B2(n_109),
.C1(n_110),
.C2(n_161),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1542),
.A2(n_103),
.B1(n_105),
.B2(n_109),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1495),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_SL g1718 ( 
.A1(n_1486),
.A2(n_110),
.B1(n_174),
.B2(n_177),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1523),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1558),
.B(n_195),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_SL g1721 ( 
.A(n_1590),
.B(n_180),
.C(n_181),
.Y(n_1721)
);

NAND2xp33_ASAP7_75t_SL g1722 ( 
.A(n_1542),
.B(n_182),
.Y(n_1722)
);

BUFx3_ASAP7_75t_L g1723 ( 
.A(n_1565),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1566),
.B(n_188),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1478),
.Y(n_1725)
);

INVx5_ASAP7_75t_L g1726 ( 
.A(n_1463),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1565),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_SL g1728 ( 
.A(n_1419),
.B(n_191),
.C(n_192),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1436),
.A2(n_1486),
.B1(n_1442),
.B2(n_1514),
.C(n_1563),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1586),
.B(n_1589),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1558),
.A2(n_1419),
.B1(n_1589),
.B2(n_1586),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1579),
.B(n_1485),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1485),
.Y(n_1733)
);

OAI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1508),
.A2(n_1533),
.B1(n_1526),
.B2(n_1466),
.Y(n_1734)
);

OAI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1492),
.A2(n_1493),
.B(n_1434),
.Y(n_1735)
);

OAI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1508),
.A2(n_1533),
.B1(n_1526),
.B2(n_1466),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1592),
.Y(n_1737)
);

INVx6_ASAP7_75t_L g1738 ( 
.A(n_1579),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1521),
.A2(n_1534),
.B1(n_1575),
.B2(n_1585),
.Y(n_1739)
);

CKINVDCx16_ASAP7_75t_R g1740 ( 
.A(n_1579),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1494),
.B(n_1501),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1521),
.A2(n_1444),
.B(n_1581),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1534),
.A2(n_1585),
.B1(n_1427),
.B2(n_1519),
.Y(n_1743)
);

CKINVDCx6p67_ASAP7_75t_R g1744 ( 
.A(n_1503),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1534),
.A2(n_1585),
.B1(n_1427),
.B2(n_1519),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1487),
.A2(n_1444),
.B1(n_1583),
.B2(n_1572),
.Y(n_1746)
);

NAND3xp33_ASAP7_75t_SL g1747 ( 
.A(n_1539),
.B(n_1541),
.C(n_1581),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1463),
.B(n_1583),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1444),
.A2(n_1500),
.B(n_1532),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1535),
.A2(n_1525),
.B1(n_1467),
.B2(n_1496),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1463),
.B(n_1583),
.Y(n_1751)
);

O2A1O1Ixp33_ASAP7_75t_SL g1752 ( 
.A1(n_1592),
.A2(n_1530),
.B(n_1506),
.C(n_1517),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1543),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1543),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1543),
.B(n_1572),
.Y(n_1755)
);

CKINVDCx11_ASAP7_75t_R g1756 ( 
.A(n_1530),
.Y(n_1756)
);

BUFx4f_ASAP7_75t_L g1757 ( 
.A(n_1572),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1539),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1525),
.A2(n_1496),
.B1(n_1467),
.B2(n_1506),
.C(n_1507),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1424),
.B(n_1411),
.Y(n_1760)
);

CKINVDCx16_ASAP7_75t_R g1761 ( 
.A(n_1496),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1531),
.B(n_1549),
.Y(n_1762)
);

OAI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1409),
.A2(n_1517),
.B1(n_1507),
.B2(n_1535),
.Y(n_1763)
);

O2A1O1Ixp33_ASAP7_75t_SL g1764 ( 
.A1(n_1559),
.A2(n_1562),
.B(n_1564),
.C(n_1570),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1462),
.B(n_1409),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1467),
.A2(n_1422),
.B1(n_1462),
.B2(n_1531),
.Y(n_1766)
);

OAI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1559),
.A2(n_1562),
.B1(n_1564),
.B2(n_1570),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1421),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1500),
.A2(n_1532),
.B(n_1417),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1588),
.Y(n_1770)
);

OR2x4_ASAP7_75t_L g1771 ( 
.A(n_1539),
.B(n_1541),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1531),
.B(n_1549),
.Y(n_1772)
);

AO21x2_ASAP7_75t_L g1773 ( 
.A1(n_1557),
.A2(n_1493),
.B(n_1454),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1430),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1424),
.B(n_1411),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1531),
.B(n_1549),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1541),
.A2(n_1500),
.B1(n_1454),
.B2(n_1549),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1500),
.B(n_1474),
.C(n_1424),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1424),
.B(n_1411),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1424),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1422),
.A2(n_1453),
.B1(n_1588),
.B2(n_1417),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1474),
.A2(n_1569),
.B1(n_1582),
.B2(n_1411),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1411),
.B(n_1422),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1453),
.B(n_1430),
.Y(n_1784)
);

OAI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1434),
.A2(n_1557),
.B(n_1464),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_SL g1786 ( 
.A(n_1569),
.B(n_1582),
.C(n_1497),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1421),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1453),
.A2(n_1588),
.B1(n_1417),
.B2(n_1423),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1410),
.B(n_1412),
.Y(n_1789)
);

AO21x1_ASAP7_75t_L g1790 ( 
.A1(n_1497),
.A2(n_1509),
.B(n_1476),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1593),
.A2(n_1474),
.B1(n_1520),
.B2(n_1509),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1761),
.B(n_1423),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1695),
.A2(n_1423),
.B1(n_1588),
.B2(n_1490),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1707),
.B(n_1474),
.C(n_1588),
.Y(n_1794)
);

AOI221x1_ASAP7_75t_SL g1795 ( 
.A1(n_1714),
.A2(n_1588),
.B1(n_1433),
.B2(n_1412),
.C(n_1410),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_SL g1796 ( 
.A1(n_1688),
.A2(n_1476),
.B1(n_1490),
.B2(n_1520),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1597),
.B(n_1604),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1706),
.A2(n_1588),
.B1(n_1433),
.B2(n_1537),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1632),
.B(n_1588),
.Y(n_1799)
);

CKINVDCx20_ASAP7_75t_R g1800 ( 
.A(n_1680),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1787),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1714),
.A2(n_1464),
.B1(n_1469),
.B2(n_1435),
.C(n_1438),
.Y(n_1802)
);

INVxp67_ASAP7_75t_L g1803 ( 
.A(n_1659),
.Y(n_1803)
);

OAI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1667),
.A2(n_1524),
.B1(n_1537),
.B2(n_1536),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1609),
.B(n_1553),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1779),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1740),
.A2(n_1536),
.B1(n_1524),
.B2(n_1540),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1630),
.Y(n_1808)
);

AOI222xp33_ASAP7_75t_L g1809 ( 
.A1(n_1658),
.A2(n_1469),
.B1(n_1438),
.B2(n_1435),
.C1(n_1445),
.C2(n_1553),
.Y(n_1809)
);

INVx8_ASAP7_75t_L g1810 ( 
.A(n_1623),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_SL g1811 ( 
.A1(n_1666),
.A2(n_1445),
.B1(n_1561),
.B2(n_1552),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1625),
.A2(n_1540),
.B1(n_1552),
.B2(n_1561),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1730),
.B(n_1665),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1658),
.A2(n_1673),
.B1(n_1703),
.B2(n_1702),
.C(n_1679),
.Y(n_1814)
);

OAI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1694),
.A2(n_1703),
.B1(n_1702),
.B2(n_1708),
.C(n_1677),
.Y(n_1815)
);

AOI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1677),
.A2(n_1692),
.B1(n_1694),
.B2(n_1708),
.C(n_1716),
.Y(n_1816)
);

OAI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1692),
.A2(n_1716),
.B1(n_1670),
.B2(n_1696),
.C(n_1600),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1626),
.B(n_1612),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1648),
.A2(n_1600),
.B1(n_1699),
.B2(n_1610),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1721),
.A2(n_1641),
.B1(n_1722),
.B2(n_1652),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1648),
.A2(n_1690),
.B1(n_1744),
.B2(n_1738),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1607),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_SL g1823 ( 
.A1(n_1674),
.A2(n_1646),
.B1(n_1608),
.B2(n_1710),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1641),
.A2(n_1722),
.B1(n_1613),
.B2(n_1594),
.Y(n_1824)
);

OA21x2_ASAP7_75t_L g1825 ( 
.A1(n_1617),
.A2(n_1769),
.B(n_1778),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_SL g1826 ( 
.A1(n_1674),
.A2(n_1646),
.B1(n_1608),
.B2(n_1685),
.Y(n_1826)
);

BUFx3_ASAP7_75t_L g1827 ( 
.A(n_1668),
.Y(n_1827)
);

OAI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1661),
.A2(n_1728),
.B(n_1605),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_L g1829 ( 
.A(n_1605),
.B(n_1718),
.C(n_1729),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1738),
.A2(n_1637),
.B1(n_1619),
.B2(n_1698),
.Y(n_1830)
);

OAI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1663),
.A2(n_1705),
.B1(n_1713),
.B2(n_1687),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1700),
.A2(n_1631),
.B1(n_1756),
.B2(n_1608),
.Y(n_1832)
);

BUFx4f_ASAP7_75t_SL g1833 ( 
.A(n_1719),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1700),
.A2(n_1756),
.B1(n_1738),
.B2(n_1736),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1734),
.A2(n_1736),
.B1(n_1596),
.B2(n_1672),
.Y(n_1835)
);

AOI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1715),
.A2(n_1734),
.B1(n_1639),
.B2(n_1616),
.C(n_1662),
.Y(n_1836)
);

OAI21x1_ASAP7_75t_L g1837 ( 
.A1(n_1598),
.A2(n_1735),
.B(n_1785),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1697),
.B(n_1627),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1596),
.A2(n_1672),
.B1(n_1623),
.B2(n_1628),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1689),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1628),
.A2(n_1720),
.B1(n_1732),
.B2(n_1611),
.Y(n_1841)
);

AO31x2_ASAP7_75t_L g1842 ( 
.A1(n_1617),
.A2(n_1777),
.A3(n_1790),
.B(n_1742),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1618),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1642),
.Y(n_1844)
);

OAI33xp33_ASAP7_75t_L g1845 ( 
.A1(n_1645),
.A2(n_1647),
.A3(n_1682),
.B1(n_1616),
.B2(n_1606),
.B3(n_1775),
.Y(n_1845)
);

AOI211xp5_ASAP7_75t_L g1846 ( 
.A1(n_1678),
.A2(n_1643),
.B(n_1724),
.C(n_1635),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1614),
.A2(n_1620),
.B1(n_1657),
.B2(n_1634),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1755),
.B(n_1753),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1651),
.B(n_1780),
.Y(n_1849)
);

OAI211xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1731),
.A2(n_1739),
.B(n_1745),
.C(n_1743),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1760),
.B(n_1693),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1644),
.A2(n_1601),
.B1(n_1711),
.B2(n_1671),
.Y(n_1852)
);

AO221x2_ASAP7_75t_L g1853 ( 
.A1(n_1763),
.A2(n_1746),
.B1(n_1650),
.B2(n_1621),
.C(n_1767),
.Y(n_1853)
);

OAI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1671),
.A2(n_1687),
.B1(n_1711),
.B2(n_1701),
.Y(n_1854)
);

OAI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1681),
.A2(n_1601),
.B1(n_1669),
.B2(n_1668),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1649),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1655),
.A2(n_1668),
.B1(n_1615),
.B2(n_1602),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_1770),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_SL g1859 ( 
.A1(n_1757),
.A2(n_1709),
.B1(n_1660),
.B2(n_1602),
.Y(n_1859)
);

OA21x2_ASAP7_75t_L g1860 ( 
.A1(n_1749),
.A2(n_1766),
.B(n_1745),
.Y(n_1860)
);

OAI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1595),
.A2(n_1650),
.B1(n_1757),
.B2(n_1684),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1615),
.A2(n_1660),
.B1(n_1622),
.B2(n_1739),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1741),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_SL g1864 ( 
.A1(n_1622),
.A2(n_1603),
.B1(n_1776),
.B2(n_1772),
.Y(n_1864)
);

INVx5_ASAP7_75t_SL g1865 ( 
.A(n_1773),
.Y(n_1865)
);

OAI222xp33_ASAP7_75t_L g1866 ( 
.A1(n_1638),
.A2(n_1731),
.B1(n_1743),
.B2(n_1712),
.C1(n_1683),
.C2(n_1733),
.Y(n_1866)
);

OAI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1771),
.A2(n_1723),
.B1(n_1727),
.B2(n_1726),
.Y(n_1867)
);

BUFx2_ASAP7_75t_L g1868 ( 
.A(n_1771),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1624),
.A2(n_1752),
.B(n_1764),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1723),
.B(n_1748),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1640),
.A2(n_1638),
.B1(n_1636),
.B2(n_1754),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1754),
.A2(n_1693),
.B1(n_1737),
.B2(n_1725),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1750),
.A2(n_1726),
.B1(n_1737),
.B2(n_1751),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1762),
.A2(n_1784),
.B1(n_1759),
.B2(n_1747),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1750),
.A2(n_1726),
.B1(n_1766),
.B2(n_1599),
.Y(n_1875)
);

AOI21x1_ASAP7_75t_L g1876 ( 
.A1(n_1765),
.A2(n_1774),
.B(n_1783),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1599),
.A2(n_1654),
.B1(n_1653),
.B2(n_1633),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1763),
.A2(n_1765),
.B1(n_1767),
.B2(n_1788),
.C(n_1752),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1726),
.A2(n_1654),
.B1(n_1653),
.B2(n_1788),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1629),
.A2(n_1633),
.B1(n_1717),
.B2(n_1691),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1618),
.A2(n_1656),
.B1(n_1664),
.B2(n_1704),
.Y(n_1881)
);

OAI211xp5_ASAP7_75t_SL g1882 ( 
.A1(n_1781),
.A2(n_1676),
.B(n_1691),
.C(n_1717),
.Y(n_1882)
);

AOI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1786),
.A2(n_1618),
.B1(n_1656),
.B2(n_1664),
.Y(n_1883)
);

OAI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1781),
.A2(n_1782),
.B(n_1675),
.Y(n_1884)
);

AOI21xp33_ASAP7_75t_L g1885 ( 
.A1(n_1676),
.A2(n_1773),
.B(n_1768),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1768),
.B(n_1789),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1789),
.B(n_1656),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1656),
.A2(n_1664),
.B1(n_1686),
.B2(n_1704),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1664),
.A2(n_1550),
.B1(n_1695),
.B2(n_1279),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1686),
.A2(n_1550),
.B1(n_1695),
.B2(n_1279),
.Y(n_1890)
);

INVx3_ASAP7_75t_L g1891 ( 
.A(n_1686),
.Y(n_1891)
);

AOI221xp5_ASAP7_75t_L g1892 ( 
.A1(n_1686),
.A2(n_1714),
.B1(n_1279),
.B2(n_492),
.C(n_527),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1704),
.Y(n_1893)
);

AOI222xp33_ASAP7_75t_L g1894 ( 
.A1(n_1704),
.A2(n_1191),
.B1(n_1005),
.B2(n_1658),
.C1(n_1695),
.C2(n_1688),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1630),
.Y(n_1895)
);

AOI21xp33_ASAP7_75t_L g1896 ( 
.A1(n_1641),
.A2(n_1279),
.B(n_1082),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1630),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1597),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1758),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1632),
.B(n_1626),
.Y(n_1900)
);

AOI221xp5_ASAP7_75t_L g1901 ( 
.A1(n_1714),
.A2(n_1279),
.B1(n_492),
.B2(n_527),
.C(n_518),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_SL g1902 ( 
.A1(n_1688),
.A2(n_1279),
.B1(n_1550),
.B2(n_1082),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1903)
);

OAI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1667),
.A2(n_1279),
.B1(n_1082),
.B2(n_788),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1597),
.Y(n_1908)
);

AOI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1593),
.A2(n_1279),
.B1(n_1082),
.B2(n_1106),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1593),
.A2(n_1279),
.B1(n_1082),
.B2(n_1106),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1761),
.B(n_1632),
.Y(n_1914)
);

OAI211xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1648),
.A2(n_1418),
.B(n_1081),
.C(n_1047),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1597),
.B(n_1604),
.Y(n_1917)
);

OAI211xp5_ASAP7_75t_L g1918 ( 
.A1(n_1658),
.A2(n_1279),
.B(n_1694),
.C(n_765),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1632),
.B(n_1626),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1761),
.B(n_1632),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1921)
);

AOI22xp33_ASAP7_75t_L g1922 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1922)
);

NOR2x1_ASAP7_75t_L g1923 ( 
.A(n_1671),
.B(n_1481),
.Y(n_1923)
);

BUFx4f_ASAP7_75t_L g1924 ( 
.A(n_1700),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_L g1925 ( 
.A(n_1618),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1593),
.A2(n_1279),
.B1(n_1082),
.B2(n_1106),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1597),
.B(n_1604),
.Y(n_1930)
);

OAI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1667),
.A2(n_1279),
.B1(n_1082),
.B2(n_788),
.Y(n_1931)
);

AOI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1932)
);

INVx2_ASAP7_75t_SL g1933 ( 
.A(n_1771),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1935)
);

AO221x2_ASAP7_75t_L g1936 ( 
.A1(n_1714),
.A2(n_1707),
.B1(n_1616),
.B2(n_1667),
.C(n_1715),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_SL g1937 ( 
.A1(n_1688),
.A2(n_1279),
.B1(n_1550),
.B2(n_1082),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1597),
.Y(n_1938)
);

AOI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1761),
.B(n_1632),
.Y(n_1940)
);

AOI21xp33_ASAP7_75t_SL g1941 ( 
.A1(n_1688),
.A2(n_734),
.B(n_1082),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1761),
.B(n_1632),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1761),
.B(n_1632),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1944)
);

AOI21xp33_ASAP7_75t_L g1945 ( 
.A1(n_1641),
.A2(n_1279),
.B(n_1082),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1597),
.Y(n_1946)
);

AO21x2_ASAP7_75t_L g1947 ( 
.A1(n_1786),
.A2(n_1598),
.B(n_1603),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1730),
.B(n_1279),
.Y(n_1948)
);

OA21x2_ASAP7_75t_L g1949 ( 
.A1(n_1617),
.A2(n_1769),
.B(n_1778),
.Y(n_1949)
);

OAI211xp5_ASAP7_75t_L g1950 ( 
.A1(n_1658),
.A2(n_1279),
.B(n_1694),
.C(n_765),
.Y(n_1950)
);

AOI221xp5_ASAP7_75t_L g1951 ( 
.A1(n_1714),
.A2(n_1279),
.B1(n_492),
.B2(n_527),
.C(n_518),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1761),
.B(n_1632),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1632),
.B(n_1626),
.Y(n_1955)
);

OR2x2_ASAP7_75t_SL g1956 ( 
.A(n_1695),
.B(n_1740),
.Y(n_1956)
);

AOI211xp5_ASAP7_75t_SL g1957 ( 
.A1(n_1715),
.A2(n_1279),
.B(n_1714),
.C(n_1666),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1958)
);

OAI21x1_ASAP7_75t_L g1959 ( 
.A1(n_1598),
.A2(n_1735),
.B(n_1785),
.Y(n_1959)
);

AOI22xp33_ASAP7_75t_L g1960 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1597),
.Y(n_1961)
);

BUFx5_ASAP7_75t_L g1962 ( 
.A(n_1787),
.Y(n_1962)
);

OAI221xp5_ASAP7_75t_L g1963 ( 
.A1(n_1707),
.A2(n_1279),
.B1(n_1082),
.B2(n_1106),
.C(n_1560),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1597),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1695),
.A2(n_1550),
.B1(n_1279),
.B2(n_1688),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1801),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1801),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1799),
.B(n_1806),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1799),
.B(n_1806),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1863),
.B(n_1856),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1876),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1962),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1822),
.Y(n_1973)
);

OAI211xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1901),
.A2(n_1951),
.B(n_1963),
.C(n_1892),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1900),
.B(n_1919),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1900),
.B(n_1919),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1962),
.Y(n_1977)
);

BUFx3_ASAP7_75t_L g1978 ( 
.A(n_1858),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1886),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1914),
.B(n_1920),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1887),
.B(n_1933),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1914),
.B(n_1920),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1844),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1955),
.B(n_1849),
.Y(n_1984)
);

OR2x2_ASAP7_75t_SL g1985 ( 
.A(n_1829),
.B(n_1794),
.Y(n_1985)
);

BUFx2_ASAP7_75t_L g1986 ( 
.A(n_1868),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1849),
.B(n_1818),
.Y(n_1987)
);

AOI22xp33_ASAP7_75t_L g1988 ( 
.A1(n_1936),
.A2(n_1902),
.B1(n_1937),
.B2(n_1816),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1940),
.B(n_1942),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1908),
.Y(n_1990)
);

INVx2_ASAP7_75t_SL g1991 ( 
.A(n_1797),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1851),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1808),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1851),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1860),
.Y(n_1995)
);

AND2x4_ASAP7_75t_L g1996 ( 
.A(n_1933),
.B(n_1868),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1938),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1940),
.B(n_1942),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1946),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1833),
.B(n_1948),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1936),
.A2(n_1815),
.B1(n_1960),
.B2(n_1928),
.Y(n_2001)
);

BUFx4f_ASAP7_75t_SL g2002 ( 
.A(n_1800),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1943),
.B(n_1952),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1943),
.B(n_1952),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1884),
.Y(n_2005)
);

BUFx3_ASAP7_75t_L g2006 ( 
.A(n_1827),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1860),
.B(n_1853),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1838),
.B(n_1803),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1860),
.B(n_1853),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1961),
.B(n_1797),
.Y(n_2010)
);

INVxp33_ASAP7_75t_L g2011 ( 
.A(n_1813),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1898),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1792),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1800),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1823),
.B(n_1792),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_1797),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1964),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1874),
.B(n_1862),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1853),
.B(n_1864),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1825),
.B(n_1949),
.Y(n_2020)
);

BUFx2_ASAP7_75t_L g2021 ( 
.A(n_1917),
.Y(n_2021)
);

BUFx3_ASAP7_75t_L g2022 ( 
.A(n_1827),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1825),
.B(n_1949),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1825),
.B(n_1949),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1842),
.B(n_1865),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1873),
.B(n_1842),
.Y(n_2026)
);

AND2x4_ASAP7_75t_SL g2027 ( 
.A(n_1848),
.B(n_1835),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1917),
.B(n_1930),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1930),
.Y(n_2029)
);

NOR2xp67_ASAP7_75t_R g2030 ( 
.A(n_1936),
.B(n_1910),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1930),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1795),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_1842),
.Y(n_2033)
);

OR2x2_ASAP7_75t_L g2034 ( 
.A(n_1842),
.B(n_1895),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1842),
.B(n_1897),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1865),
.B(n_1885),
.Y(n_2036)
);

HB1xp67_ASAP7_75t_L g2037 ( 
.A(n_1878),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1837),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1883),
.Y(n_2039)
);

OAI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1903),
.A2(n_1965),
.B1(n_1912),
.B2(n_1911),
.Y(n_2040)
);

NOR2xp67_ASAP7_75t_L g2041 ( 
.A(n_1869),
.B(n_1805),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1959),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1959),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1843),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1865),
.B(n_1871),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1947),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1865),
.B(n_1847),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1879),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1947),
.B(n_1826),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1967),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1968),
.B(n_1857),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1974),
.A2(n_1896),
.B1(n_1945),
.B2(n_1929),
.Y(n_2052)
);

BUFx10_ASAP7_75t_L g2053 ( 
.A(n_2014),
.Y(n_2053)
);

NAND2xp33_ASAP7_75t_SL g2054 ( 
.A(n_1988),
.B(n_1913),
.Y(n_2054)
);

AOI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1974),
.A2(n_2040),
.B1(n_2005),
.B2(n_2001),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_2030),
.A2(n_1828),
.B(n_1918),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1998),
.B(n_1840),
.Y(n_2057)
);

OAI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_2040),
.A2(n_1957),
.B1(n_1817),
.B2(n_1941),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1985),
.A2(n_1958),
.B1(n_1927),
.B2(n_1926),
.Y(n_2059)
);

BUFx2_ASAP7_75t_L g2060 ( 
.A(n_1986),
.Y(n_2060)
);

OAI221xp5_ASAP7_75t_L g2061 ( 
.A1(n_2037),
.A2(n_1916),
.B1(n_1906),
.B2(n_1907),
.C(n_1905),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_2013),
.Y(n_2062)
);

AO21x2_ASAP7_75t_L g2063 ( 
.A1(n_2046),
.A2(n_1947),
.B(n_1850),
.Y(n_2063)
);

OAI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_2037),
.A2(n_1819),
.B1(n_1814),
.B2(n_1904),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_1991),
.B(n_1899),
.Y(n_2065)
);

OR2x6_ASAP7_75t_L g2066 ( 
.A(n_2007),
.B(n_1875),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1967),
.Y(n_2067)
);

NAND3xp33_ASAP7_75t_L g2068 ( 
.A(n_2032),
.B(n_1935),
.C(n_1932),
.Y(n_2068)
);

NAND2xp33_ASAP7_75t_R g2069 ( 
.A(n_2005),
.B(n_1870),
.Y(n_2069)
);

INVx3_ASAP7_75t_L g2070 ( 
.A(n_2010),
.Y(n_2070)
);

AO21x2_ASAP7_75t_L g2071 ( 
.A1(n_2046),
.A2(n_1866),
.B(n_1812),
.Y(n_2071)
);

INVx4_ASAP7_75t_L g2072 ( 
.A(n_2044),
.Y(n_2072)
);

NOR2xp67_ASAP7_75t_L g2073 ( 
.A(n_1971),
.B(n_1899),
.Y(n_2073)
);

AOI221xp5_ASAP7_75t_L g2074 ( 
.A1(n_2032),
.A2(n_1931),
.B1(n_1831),
.B2(n_1921),
.C(n_1922),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1998),
.B(n_1824),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_SL g2076 ( 
.A1(n_2019),
.A2(n_1950),
.B1(n_1924),
.B2(n_1821),
.Y(n_2076)
);

OAI221xp5_ASAP7_75t_L g2077 ( 
.A1(n_2018),
.A2(n_1944),
.B1(n_1934),
.B2(n_1939),
.C(n_1909),
.Y(n_2077)
);

OAI22xp5_ASAP7_75t_SL g2078 ( 
.A1(n_1985),
.A2(n_1954),
.B1(n_1953),
.B2(n_1956),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1968),
.B(n_1832),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1966),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_2018),
.A2(n_1894),
.B1(n_1915),
.B2(n_1820),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2019),
.A2(n_1889),
.B1(n_1890),
.B2(n_1834),
.Y(n_2082)
);

AOI221xp5_ASAP7_75t_L g2083 ( 
.A1(n_2019),
.A2(n_1836),
.B1(n_1845),
.B2(n_1830),
.C(n_1854),
.Y(n_2083)
);

AND4x1_ASAP7_75t_L g2084 ( 
.A(n_2049),
.B(n_1852),
.C(n_1923),
.D(n_2009),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_2047),
.A2(n_1924),
.B1(n_1841),
.B2(n_1861),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1983),
.Y(n_2086)
);

NOR4xp25_ASAP7_75t_L g2087 ( 
.A(n_2049),
.B(n_1855),
.C(n_1867),
.D(n_1882),
.Y(n_2087)
);

AOI221xp5_ASAP7_75t_L g2088 ( 
.A1(n_2007),
.A2(n_1872),
.B1(n_1793),
.B2(n_1804),
.C(n_1846),
.Y(n_2088)
);

OAI33xp33_ASAP7_75t_L g2089 ( 
.A1(n_2034),
.A2(n_1881),
.A3(n_1791),
.B1(n_1807),
.B2(n_1956),
.B3(n_1859),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2047),
.A2(n_1924),
.B1(n_1810),
.B2(n_1796),
.Y(n_2090)
);

NAND5xp2_ASAP7_75t_SL g2091 ( 
.A(n_2030),
.B(n_1888),
.C(n_1798),
.D(n_1877),
.E(n_1839),
.Y(n_2091)
);

AOI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_2047),
.A2(n_1810),
.B1(n_1811),
.B2(n_1802),
.Y(n_2092)
);

OR2x2_ASAP7_75t_L g2093 ( 
.A(n_2013),
.B(n_1893),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1966),
.Y(n_2094)
);

AOI211xp5_ASAP7_75t_SL g2095 ( 
.A1(n_2049),
.A2(n_1891),
.B(n_1810),
.C(n_1809),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1990),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_1980),
.B(n_1880),
.Y(n_2097)
);

AOI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_2045),
.A2(n_2009),
.B1(n_2007),
.B2(n_2048),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_R g2099 ( 
.A(n_2002),
.B(n_1925),
.Y(n_2099)
);

NAND3xp33_ASAP7_75t_L g2100 ( 
.A(n_2039),
.B(n_1925),
.C(n_2048),
.Y(n_2100)
);

AOI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_2045),
.A2(n_2009),
.B1(n_2027),
.B2(n_2039),
.Y(n_2101)
);

AO21x2_ASAP7_75t_L g2102 ( 
.A1(n_2038),
.A2(n_2042),
.B(n_2043),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_2045),
.A2(n_2027),
.B1(n_2015),
.B2(n_2000),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1997),
.Y(n_2104)
);

INVxp67_ASAP7_75t_L g2105 ( 
.A(n_2008),
.Y(n_2105)
);

OA21x2_ASAP7_75t_L g2106 ( 
.A1(n_2020),
.A2(n_2024),
.B(n_2023),
.Y(n_2106)
);

NAND2xp33_ASAP7_75t_SL g2107 ( 
.A(n_2011),
.B(n_2021),
.Y(n_2107)
);

OAI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_2027),
.A2(n_2041),
.B1(n_1993),
.B2(n_1978),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_1968),
.B(n_1969),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1997),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1969),
.B(n_1989),
.Y(n_2111)
);

OA21x2_ASAP7_75t_L g2112 ( 
.A1(n_2020),
.A2(n_2023),
.B(n_2024),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1969),
.B(n_1989),
.Y(n_2113)
);

OAI221xp5_ASAP7_75t_L g2114 ( 
.A1(n_1993),
.A2(n_2026),
.B1(n_2035),
.B2(n_2034),
.C(n_1986),
.Y(n_2114)
);

NOR2x2_ASAP7_75t_L g2115 ( 
.A(n_1999),
.B(n_1972),
.Y(n_2115)
);

AOI33xp33_ASAP7_75t_L g2116 ( 
.A1(n_2015),
.A2(n_2024),
.A3(n_2023),
.B1(n_2020),
.B2(n_2012),
.B3(n_2017),
.Y(n_2116)
);

AOI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_1996),
.A2(n_1989),
.B1(n_2004),
.B2(n_2003),
.Y(n_2117)
);

AOI31xp33_ASAP7_75t_SL g2118 ( 
.A1(n_2026),
.A2(n_2035),
.A3(n_1980),
.B(n_1982),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1973),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2003),
.B(n_2004),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1973),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2106),
.B(n_1995),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2050),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_R g2124 ( 
.A(n_2069),
.B(n_2006),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2106),
.Y(n_2125)
);

BUFx2_ASAP7_75t_L g2126 ( 
.A(n_2115),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2050),
.Y(n_2127)
);

INVx6_ASAP7_75t_L g2128 ( 
.A(n_2053),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2067),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2116),
.B(n_1992),
.Y(n_2130)
);

OR2x2_ASAP7_75t_L g2131 ( 
.A(n_2106),
.B(n_1982),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2106),
.B(n_1995),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2112),
.Y(n_2133)
);

INVx2_ASAP7_75t_SL g2134 ( 
.A(n_2070),
.Y(n_2134)
);

AND2x2_ASAP7_75t_SL g2135 ( 
.A(n_2084),
.B(n_1995),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2062),
.B(n_1992),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2112),
.B(n_1995),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2112),
.B(n_1995),
.Y(n_2138)
);

NAND3xp33_ASAP7_75t_L g2139 ( 
.A(n_2054),
.B(n_2033),
.C(n_1995),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2112),
.B(n_1995),
.Y(n_2140)
);

OAI21xp33_ASAP7_75t_SL g2141 ( 
.A1(n_2066),
.A2(n_1991),
.B(n_2016),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2120),
.B(n_2093),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_2105),
.B(n_2028),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2109),
.B(n_2025),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2109),
.B(n_2025),
.Y(n_2145)
);

OR2x2_ASAP7_75t_L g2146 ( 
.A(n_2093),
.B(n_1994),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2111),
.B(n_2025),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2121),
.B(n_1994),
.Y(n_2148)
);

BUFx2_ASAP7_75t_L g2149 ( 
.A(n_2115),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2111),
.B(n_1975),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2113),
.B(n_1975),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2121),
.B(n_2003),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2113),
.B(n_1975),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2060),
.B(n_2033),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2070),
.B(n_2066),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2102),
.Y(n_2156)
);

AND2x4_ASAP7_75t_SL g2157 ( 
.A(n_2065),
.B(n_2010),
.Y(n_2157)
);

NOR3xp33_ASAP7_75t_L g2158 ( 
.A(n_2054),
.B(n_2036),
.C(n_1970),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2066),
.B(n_1976),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2102),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2080),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_2060),
.B(n_1979),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_2114),
.B(n_1979),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2066),
.B(n_1976),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2080),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2094),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2117),
.B(n_1987),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2094),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2051),
.B(n_1987),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2119),
.B(n_2096),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2104),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_2072),
.B(n_1977),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2110),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2051),
.B(n_1987),
.Y(n_2174)
);

BUFx2_ASAP7_75t_L g2175 ( 
.A(n_2107),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2071),
.B(n_1984),
.Y(n_2176)
);

BUFx2_ASAP7_75t_L g2177 ( 
.A(n_2107),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2086),
.B(n_1971),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2071),
.B(n_1984),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2119),
.B(n_2004),
.Y(n_2180)
);

INVx1_ASAP7_75t_SL g2181 ( 
.A(n_2124),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2126),
.B(n_2079),
.Y(n_2182)
);

INVx2_ASAP7_75t_SL g2183 ( 
.A(n_2157),
.Y(n_2183)
);

OR2x6_ASAP7_75t_L g2184 ( 
.A(n_2139),
.B(n_2056),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2130),
.B(n_2097),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2161),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2161),
.Y(n_2187)
);

INVxp67_ASAP7_75t_L g2188 ( 
.A(n_2143),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2126),
.B(n_2149),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2149),
.B(n_2159),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2165),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2165),
.Y(n_2192)
);

AOI221xp5_ASAP7_75t_L g2193 ( 
.A1(n_2158),
.A2(n_2058),
.B1(n_2059),
.B2(n_2055),
.C(n_2064),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2156),
.Y(n_2194)
);

OR2x2_ASAP7_75t_L g2195 ( 
.A(n_2130),
.B(n_2097),
.Y(n_2195)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2196 ( 
.A1(n_2135),
.A2(n_2061),
.B(n_2077),
.C(n_2082),
.D(n_2078),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2166),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2156),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_2157),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2158),
.B(n_2057),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2159),
.B(n_2079),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2169),
.B(n_2029),
.Y(n_2202)
);

INVxp33_ASAP7_75t_L g2203 ( 
.A(n_2152),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2156),
.Y(n_2204)
);

BUFx3_ASAP7_75t_L g2205 ( 
.A(n_2128),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2169),
.B(n_2029),
.Y(n_2206)
);

NOR2x1_ASAP7_75t_L g2207 ( 
.A(n_2175),
.B(n_2100),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2166),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2168),
.Y(n_2209)
);

INVxp33_ASAP7_75t_L g2210 ( 
.A(n_2152),
.Y(n_2210)
);

NAND3xp33_ASAP7_75t_L g2211 ( 
.A(n_2139),
.B(n_2052),
.C(n_2081),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2168),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_2131),
.B(n_2063),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2123),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2159),
.B(n_2072),
.Y(n_2215)
);

OR2x6_ASAP7_75t_L g2216 ( 
.A(n_2175),
.B(n_2108),
.Y(n_2216)
);

INVxp67_ASAP7_75t_L g2217 ( 
.A(n_2136),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2123),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2127),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2164),
.B(n_2176),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2131),
.B(n_2063),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_SL g2222 ( 
.A(n_2135),
.B(n_2091),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2127),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2129),
.Y(n_2224)
);

INVx2_ASAP7_75t_SL g2225 ( 
.A(n_2157),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_2128),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2160),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2164),
.B(n_2072),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2169),
.B(n_2031),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2129),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_2128),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2171),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2131),
.B(n_2063),
.Y(n_2233)
);

AOI32xp33_ASAP7_75t_L g2234 ( 
.A1(n_2177),
.A2(n_2095),
.A3(n_2074),
.B1(n_2076),
.B2(n_2098),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2187),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_2185),
.B(n_2195),
.Y(n_2236)
);

OR2x6_ASAP7_75t_L g2237 ( 
.A(n_2184),
.B(n_2128),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2187),
.Y(n_2238)
);

AND2x4_ASAP7_75t_SL g2239 ( 
.A(n_2184),
.B(n_2164),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2200),
.B(n_2174),
.Y(n_2240)
);

NOR3xp33_ASAP7_75t_SL g2241 ( 
.A(n_2211),
.B(n_2089),
.C(n_2068),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2189),
.B(n_2176),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2189),
.B(n_2176),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2194),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2182),
.B(n_2179),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2182),
.B(n_2179),
.Y(n_2246)
);

OR2x6_ASAP7_75t_L g2247 ( 
.A(n_2184),
.B(n_2128),
.Y(n_2247)
);

NOR2x1_ASAP7_75t_L g2248 ( 
.A(n_2207),
.B(n_2177),
.Y(n_2248)
);

NAND3xp33_ASAP7_75t_SL g2249 ( 
.A(n_2222),
.B(n_2087),
.C(n_2083),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2190),
.B(n_2179),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_2194),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2188),
.B(n_2174),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2190),
.B(n_2135),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2191),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2191),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2192),
.Y(n_2256)
);

BUFx2_ASAP7_75t_L g2257 ( 
.A(n_2184),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2185),
.B(n_2174),
.Y(n_2258)
);

NAND2xp33_ASAP7_75t_SL g2259 ( 
.A(n_2196),
.B(n_2099),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2192),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2198),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2198),
.Y(n_2262)
);

INVxp67_ASAP7_75t_L g2263 ( 
.A(n_2195),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2204),
.Y(n_2264)
);

BUFx3_ASAP7_75t_L g2265 ( 
.A(n_2205),
.Y(n_2265)
);

BUFx2_ASAP7_75t_L g2266 ( 
.A(n_2205),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2201),
.B(n_2155),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2204),
.Y(n_2268)
);

NAND2xp33_ASAP7_75t_SL g2269 ( 
.A(n_2183),
.B(n_2167),
.Y(n_2269)
);

OR2x2_ASAP7_75t_L g2270 ( 
.A(n_2217),
.B(n_2163),
.Y(n_2270)
);

OR2x2_ASAP7_75t_L g2271 ( 
.A(n_2202),
.B(n_2163),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2227),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2234),
.B(n_2150),
.Y(n_2273)
);

BUFx5_ASAP7_75t_L g2274 ( 
.A(n_2231),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2197),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2197),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2208),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2208),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_2206),
.B(n_2229),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_L g2280 ( 
.A(n_2181),
.B(n_2053),
.Y(n_2280)
);

OR2x6_ASAP7_75t_L g2281 ( 
.A(n_2216),
.B(n_2231),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2201),
.B(n_2155),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2193),
.B(n_2150),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2220),
.B(n_2155),
.Y(n_2284)
);

NOR2xp33_ASAP7_75t_R g2285 ( 
.A(n_2226),
.B(n_2053),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2283),
.B(n_2220),
.Y(n_2286)
);

INVxp67_ASAP7_75t_SL g2287 ( 
.A(n_2248),
.Y(n_2287)
);

AOI211xp5_ASAP7_75t_L g2288 ( 
.A1(n_2249),
.A2(n_2118),
.B(n_2088),
.C(n_2141),
.Y(n_2288)
);

OAI21xp5_ASAP7_75t_SL g2289 ( 
.A1(n_2273),
.A2(n_2103),
.B(n_2092),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2241),
.B(n_2150),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2235),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2236),
.B(n_2240),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2236),
.B(n_2142),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_2265),
.B(n_2266),
.Y(n_2294)
);

OAI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2248),
.A2(n_2216),
.B(n_2141),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2235),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2263),
.B(n_2151),
.Y(n_2297)
);

INVx1_ASAP7_75t_SL g2298 ( 
.A(n_2285),
.Y(n_2298)
);

OAI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2257),
.A2(n_2216),
.B1(n_2075),
.B2(n_2091),
.Y(n_2299)
);

AOI322xp5_ASAP7_75t_L g2300 ( 
.A1(n_2259),
.A2(n_2122),
.A3(n_2140),
.B1(n_2138),
.B2(n_2137),
.C1(n_2132),
.C2(n_2167),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2253),
.B(n_2215),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2257),
.B(n_2151),
.Y(n_2302)
);

INVxp67_ASAP7_75t_L g2303 ( 
.A(n_2266),
.Y(n_2303)
);

OAI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2253),
.A2(n_2216),
.B(n_2215),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2280),
.B(n_2203),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2281),
.A2(n_2101),
.B1(n_2183),
.B2(n_2225),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2238),
.Y(n_2307)
);

AOI21xp33_ASAP7_75t_L g2308 ( 
.A1(n_2237),
.A2(n_2210),
.B(n_2213),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2238),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2254),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2252),
.B(n_2151),
.Y(n_2311)
);

OAI21xp33_ASAP7_75t_SL g2312 ( 
.A1(n_2281),
.A2(n_2225),
.B(n_2228),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2267),
.B(n_2228),
.Y(n_2313)
);

AOI21xp5_ASAP7_75t_L g2314 ( 
.A1(n_2237),
.A2(n_2148),
.B(n_2136),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_SL g2315 ( 
.A(n_2281),
.B(n_2199),
.Y(n_2315)
);

AOI22xp5_ASAP7_75t_L g2316 ( 
.A1(n_2269),
.A2(n_2199),
.B1(n_2071),
.B2(n_2085),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2265),
.B(n_2153),
.Y(n_2317)
);

AOI22xp33_ASAP7_75t_L g2318 ( 
.A1(n_2237),
.A2(n_2090),
.B1(n_2140),
.B2(n_2132),
.Y(n_2318)
);

NAND4xp25_ASAP7_75t_L g2319 ( 
.A(n_2270),
.B(n_2233),
.C(n_2221),
.D(n_2213),
.Y(n_2319)
);

AOI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_2239),
.A2(n_2199),
.B1(n_1996),
.B2(n_2167),
.Y(n_2320)
);

OAI321xp33_ASAP7_75t_L g2321 ( 
.A1(n_2281),
.A2(n_2233),
.A3(n_2221),
.B1(n_2132),
.B2(n_2137),
.C(n_2138),
.Y(n_2321)
);

OAI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2237),
.A2(n_2137),
.B(n_2122),
.Y(n_2322)
);

AOI22xp5_ASAP7_75t_L g2323 ( 
.A1(n_2239),
.A2(n_1996),
.B1(n_2036),
.B2(n_1981),
.Y(n_2323)
);

AOI211x1_ASAP7_75t_SL g2324 ( 
.A1(n_2258),
.A2(n_2227),
.B(n_2073),
.C(n_2125),
.Y(n_2324)
);

INVx1_ASAP7_75t_SL g2325 ( 
.A(n_2265),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2267),
.B(n_2153),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2291),
.Y(n_2327)
);

OAI32xp33_ASAP7_75t_L g2328 ( 
.A1(n_2324),
.A2(n_2270),
.A3(n_2242),
.B1(n_2243),
.B2(n_2245),
.Y(n_2328)
);

HB1xp67_ASAP7_75t_L g2329 ( 
.A(n_2303),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2325),
.B(n_2242),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2296),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2307),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2294),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2303),
.B(n_2243),
.Y(n_2334)
);

OAI31xp33_ASAP7_75t_L g2335 ( 
.A1(n_2299),
.A2(n_2239),
.A3(n_2245),
.B(n_2246),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2301),
.B(n_2281),
.Y(n_2336)
);

AOI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2299),
.A2(n_2247),
.B(n_2237),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2309),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2310),
.Y(n_2339)
);

NOR3xp33_ASAP7_75t_L g2340 ( 
.A(n_2287),
.B(n_2271),
.C(n_2246),
.Y(n_2340)
);

OAI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2287),
.A2(n_2247),
.B1(n_2271),
.B2(n_2279),
.Y(n_2341)
);

AOI22xp5_ASAP7_75t_L g2342 ( 
.A1(n_2288),
.A2(n_2247),
.B1(n_2274),
.B2(n_2282),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2294),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2313),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2293),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2290),
.B(n_2282),
.Y(n_2346)
);

OAI21xp33_ASAP7_75t_SL g2347 ( 
.A1(n_2300),
.A2(n_2250),
.B(n_2247),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2289),
.B(n_2250),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2297),
.Y(n_2349)
);

OAI222xp33_ASAP7_75t_L g2350 ( 
.A1(n_2316),
.A2(n_2247),
.B1(n_2284),
.B2(n_2279),
.C1(n_2140),
.C2(n_2122),
.Y(n_2350)
);

AOI32xp33_ASAP7_75t_L g2351 ( 
.A1(n_2321),
.A2(n_2284),
.A3(n_2138),
.B1(n_2277),
.B2(n_2276),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2295),
.B(n_2274),
.Y(n_2352)
);

OAI21xp33_ASAP7_75t_L g2353 ( 
.A1(n_2286),
.A2(n_2255),
.B(n_2254),
.Y(n_2353)
);

OR2x2_ASAP7_75t_L g2354 ( 
.A(n_2292),
.B(n_2255),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2304),
.B(n_2298),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2317),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2305),
.B(n_2274),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2329),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_R g2359 ( 
.A(n_2355),
.B(n_2343),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_L g2360 ( 
.A(n_2355),
.B(n_2305),
.Y(n_2360)
);

AOI222xp33_ASAP7_75t_L g2361 ( 
.A1(n_2347),
.A2(n_2318),
.B1(n_2322),
.B2(n_2312),
.C1(n_2306),
.C2(n_2302),
.Y(n_2361)
);

OAI222xp33_ASAP7_75t_L g2362 ( 
.A1(n_2351),
.A2(n_2318),
.B1(n_2320),
.B2(n_2314),
.C1(n_2323),
.C2(n_2326),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2343),
.B(n_2311),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2345),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2345),
.Y(n_2365)
);

INVx1_ASAP7_75t_SL g2366 ( 
.A(n_2336),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2327),
.Y(n_2367)
);

XOR2xp5_ASAP7_75t_L g2368 ( 
.A(n_2342),
.B(n_2319),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2333),
.B(n_2315),
.Y(n_2369)
);

NOR3xp33_ASAP7_75t_L g2370 ( 
.A(n_2341),
.B(n_2308),
.C(n_2264),
.Y(n_2370)
);

NOR4xp25_ASAP7_75t_SL g2371 ( 
.A(n_2327),
.B(n_2278),
.C(n_2277),
.D(n_2276),
.Y(n_2371)
);

INVx3_ASAP7_75t_L g2372 ( 
.A(n_2333),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2331),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2336),
.B(n_2274),
.Y(n_2374)
);

INVxp67_ASAP7_75t_SL g2375 ( 
.A(n_2330),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_2335),
.B(n_2274),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2331),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2344),
.B(n_2274),
.Y(n_2378)
);

NOR2xp33_ASAP7_75t_R g2379 ( 
.A(n_2357),
.B(n_2274),
.Y(n_2379)
);

INVxp67_ASAP7_75t_L g2380 ( 
.A(n_2334),
.Y(n_2380)
);

NAND2xp33_ASAP7_75t_SL g2381 ( 
.A(n_2348),
.B(n_2256),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2332),
.Y(n_2382)
);

NOR3xp33_ASAP7_75t_L g2383 ( 
.A(n_2360),
.B(n_2337),
.C(n_2356),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2366),
.B(n_2344),
.Y(n_2384)
);

INVxp33_ASAP7_75t_L g2385 ( 
.A(n_2359),
.Y(n_2385)
);

INVxp67_ASAP7_75t_L g2386 ( 
.A(n_2369),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2372),
.B(n_2356),
.Y(n_2387)
);

OAI321xp33_ASAP7_75t_L g2388 ( 
.A1(n_2376),
.A2(n_2352),
.A3(n_2349),
.B1(n_2346),
.B2(n_2353),
.C(n_2354),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2369),
.B(n_2349),
.Y(n_2389)
);

NAND3xp33_ASAP7_75t_L g2390 ( 
.A(n_2361),
.B(n_2340),
.C(n_2339),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2372),
.B(n_2332),
.Y(n_2391)
);

AOI221xp5_ASAP7_75t_L g2392 ( 
.A1(n_2381),
.A2(n_2328),
.B1(n_2350),
.B2(n_2352),
.C(n_2338),
.Y(n_2392)
);

OAI221xp5_ASAP7_75t_L g2393 ( 
.A1(n_2368),
.A2(n_2354),
.B1(n_2338),
.B2(n_2328),
.C(n_2278),
.Y(n_2393)
);

AOI221xp5_ASAP7_75t_L g2394 ( 
.A1(n_2381),
.A2(n_2275),
.B1(n_2256),
.B2(n_2260),
.C(n_2264),
.Y(n_2394)
);

AOI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2368),
.A2(n_2274),
.B1(n_2275),
.B2(n_2260),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_2380),
.B(n_2274),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2372),
.B(n_2186),
.Y(n_2397)
);

INVx2_ASAP7_75t_SL g2398 ( 
.A(n_2374),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2385),
.B(n_2358),
.Y(n_2399)
);

AOI32xp33_ASAP7_75t_L g2400 ( 
.A1(n_2393),
.A2(n_2370),
.A3(n_2374),
.B1(n_2375),
.B2(n_2365),
.Y(n_2400)
);

A2O1A1Ixp33_ASAP7_75t_L g2401 ( 
.A1(n_2392),
.A2(n_2364),
.B(n_2365),
.C(n_2363),
.Y(n_2401)
);

OAI221xp5_ASAP7_75t_L g2402 ( 
.A1(n_2390),
.A2(n_2364),
.B1(n_2377),
.B2(n_2367),
.C(n_2373),
.Y(n_2402)
);

AOI221xp5_ASAP7_75t_L g2403 ( 
.A1(n_2388),
.A2(n_2362),
.B1(n_2382),
.B2(n_2378),
.C(n_2379),
.Y(n_2403)
);

AOI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2383),
.A2(n_2386),
.B1(n_2389),
.B2(n_2384),
.Y(n_2404)
);

NAND4xp25_ASAP7_75t_L g2405 ( 
.A(n_2395),
.B(n_2382),
.C(n_2378),
.D(n_2371),
.Y(n_2405)
);

AOI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2398),
.A2(n_2272),
.B1(n_2268),
.B2(n_2261),
.Y(n_2406)
);

AOI211xp5_ASAP7_75t_L g2407 ( 
.A1(n_2396),
.A2(n_2264),
.B(n_2251),
.C(n_2272),
.Y(n_2407)
);

OAI211xp5_ASAP7_75t_L g2408 ( 
.A1(n_2387),
.A2(n_2251),
.B(n_2262),
.C(n_2261),
.Y(n_2408)
);

OAI22xp33_ASAP7_75t_L g2409 ( 
.A1(n_2391),
.A2(n_2125),
.B1(n_2133),
.B2(n_2154),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_R g2410 ( 
.A(n_2397),
.B(n_2022),
.Y(n_2410)
);

NAND2x1_ASAP7_75t_L g2411 ( 
.A(n_2404),
.B(n_2244),
.Y(n_2411)
);

AOI221xp5_ASAP7_75t_L g2412 ( 
.A1(n_2400),
.A2(n_2394),
.B1(n_2251),
.B2(n_2262),
.C(n_2268),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_2399),
.B(n_2244),
.Y(n_2413)
);

AOI221xp5_ASAP7_75t_SL g2414 ( 
.A1(n_2401),
.A2(n_2125),
.B1(n_2133),
.B2(n_2224),
.C(n_2223),
.Y(n_2414)
);

BUFx2_ASAP7_75t_L g2415 ( 
.A(n_2410),
.Y(n_2415)
);

BUFx2_ASAP7_75t_L g2416 ( 
.A(n_2405),
.Y(n_2416)
);

AOI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_2403),
.A2(n_1996),
.B1(n_2230),
.B2(n_2224),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2415),
.B(n_2406),
.Y(n_2418)
);

NOR3xp33_ASAP7_75t_SL g2419 ( 
.A(n_2413),
.B(n_2402),
.C(n_2408),
.Y(n_2419)
);

NAND3x1_ASAP7_75t_L g2420 ( 
.A(n_2417),
.B(n_2407),
.C(n_2223),
.Y(n_2420)
);

INVx1_ASAP7_75t_SL g2421 ( 
.A(n_2411),
.Y(n_2421)
);

XNOR2xp5_ASAP7_75t_L g2422 ( 
.A(n_2416),
.B(n_2409),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_2412),
.Y(n_2423)
);

AO22x2_ASAP7_75t_L g2424 ( 
.A1(n_2414),
.A2(n_2133),
.B1(n_2230),
.B2(n_2219),
.Y(n_2424)
);

NOR2x1_ASAP7_75t_L g2425 ( 
.A(n_2415),
.B(n_2214),
.Y(n_2425)
);

NAND3xp33_ASAP7_75t_L g2426 ( 
.A(n_2419),
.B(n_2232),
.C(n_2219),
.Y(n_2426)
);

AOI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_2422),
.A2(n_2232),
.B1(n_2218),
.B2(n_2214),
.Y(n_2427)
);

AOI211xp5_ASAP7_75t_L g2428 ( 
.A1(n_2423),
.A2(n_2154),
.B(n_2212),
.C(n_2209),
.Y(n_2428)
);

OAI221xp5_ASAP7_75t_SL g2429 ( 
.A1(n_2421),
.A2(n_2154),
.B1(n_2162),
.B2(n_2146),
.C(n_2134),
.Y(n_2429)
);

NAND3xp33_ASAP7_75t_SL g2430 ( 
.A(n_2418),
.B(n_2162),
.C(n_2146),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2425),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2420),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2432),
.B(n_2431),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2427),
.B(n_2424),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2428),
.B(n_2424),
.Y(n_2435)
);

NAND3xp33_ASAP7_75t_SL g2436 ( 
.A(n_2426),
.B(n_2148),
.C(n_2178),
.Y(n_2436)
);

AOI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2435),
.A2(n_2430),
.B(n_2429),
.Y(n_2437)
);

AOI222xp33_ASAP7_75t_L g2438 ( 
.A1(n_2434),
.A2(n_2218),
.B1(n_2073),
.B2(n_2147),
.C1(n_2145),
.C2(n_2144),
.Y(n_2438)
);

INVx1_ASAP7_75t_SL g2439 ( 
.A(n_2437),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2438),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_L g2441 ( 
.A1(n_2439),
.A2(n_2436),
.B1(n_2433),
.B2(n_2160),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2440),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2439),
.Y(n_2443)
);

INVx4_ASAP7_75t_L g2444 ( 
.A(n_2443),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_2442),
.Y(n_2445)
);

AOI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2445),
.A2(n_2441),
.B1(n_2134),
.B2(n_2144),
.Y(n_2446)
);

AOI222xp33_ASAP7_75t_L g2447 ( 
.A1(n_2444),
.A2(n_2147),
.B1(n_2144),
.B2(n_2145),
.C1(n_2160),
.C2(n_2180),
.Y(n_2447)
);

AOI22xp5_ASAP7_75t_L g2448 ( 
.A1(n_2446),
.A2(n_2134),
.B1(n_2145),
.B2(n_2172),
.Y(n_2448)
);

OAI221xp5_ASAP7_75t_L g2449 ( 
.A1(n_2448),
.A2(n_2447),
.B1(n_2178),
.B2(n_2180),
.C(n_2170),
.Y(n_2449)
);

AOI211xp5_ASAP7_75t_L g2450 ( 
.A1(n_2449),
.A2(n_2178),
.B(n_2022),
.C(n_2173),
.Y(n_2450)
);


endmodule