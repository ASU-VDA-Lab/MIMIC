module fake_netlist_5_1828_n_1960 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1960);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1960;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_SL g195 ( 
.A(n_102),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_54),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_32),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_1),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_55),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_30),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_111),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_118),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_106),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_58),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

BUFx2_ASAP7_75t_SL g209 ( 
.A(n_1),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_3),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_38),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_63),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_181),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_105),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_86),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_114),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_135),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_38),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_33),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_127),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_101),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_52),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_64),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_144),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_75),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_73),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_94),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_92),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_104),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_17),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_96),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_63),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_7),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_145),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_52),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_93),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_158),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_41),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_13),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_4),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_64),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_82),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_91),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_20),
.Y(n_248)
);

BUFx8_ASAP7_75t_SL g249 ( 
.A(n_186),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_126),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_66),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_74),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_120),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_43),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_50),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_138),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_29),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_57),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_136),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_13),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_147),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_9),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_140),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_163),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_21),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_2),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_42),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_142),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_185),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_117),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_57),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_157),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_37),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_16),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_5),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_2),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_154),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_108),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_110),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_76),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_10),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_6),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_10),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_182),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_33),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_77),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_119),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_165),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_78),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_70),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_130),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_99),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_14),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_42),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_79),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_167),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_156),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_29),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_166),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_26),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_164),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_149),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_131),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_17),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_192),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_152),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_9),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_3),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_109),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_49),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_183),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_171),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_24),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_30),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_20),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_129),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_189),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_8),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_67),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_56),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_32),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_103),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_19),
.Y(n_325)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_132),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_100),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_60),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_71),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_62),
.Y(n_330)
);

BUFx5_ASAP7_75t_L g331 ( 
.A(n_115),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_116),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_59),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_133),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_153),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_39),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_155),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_28),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_21),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_62),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_8),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_24),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_124),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_71),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_27),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_45),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_35),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_12),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_58),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_18),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_148),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_18),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_146),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_180),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_122),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_69),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_68),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_143),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_87),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_151),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_162),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_6),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_56),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_98),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_176),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_95),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_36),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_161),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_141),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_46),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_11),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_150),
.Y(n_372)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_0),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_169),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_113),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_36),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_0),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_50),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_107),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_170),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_81),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_55),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_159),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_41),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_184),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_88),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_160),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_137),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_221),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_249),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_373),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_201),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_373),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_246),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_252),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_200),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_224),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_237),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_373),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_275),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_256),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_258),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_L g408 ( 
.A(n_238),
.B(n_4),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_337),
.B(n_5),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_231),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_264),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_265),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_251),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_287),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_251),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_278),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_327),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_285),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_369),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_202),
.B(n_7),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_316),
.B(n_11),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_288),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_250),
.B(n_12),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_250),
.B(n_14),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_223),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_290),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_263),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_296),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_263),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_298),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_198),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_268),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_280),
.B(n_15),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_196),
.B(n_15),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_301),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_305),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_268),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_307),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_222),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_308),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_330),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_358),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_359),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_357),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_360),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_361),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_231),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_367),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_198),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_199),
.B(n_16),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_364),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_210),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_233),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_365),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_368),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_372),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_235),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_374),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_241),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_243),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_326),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_245),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_244),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_239),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_204),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_248),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_254),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_255),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_196),
.B(n_19),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_272),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_277),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_283),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_284),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_204),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_291),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_362),
.B(n_22),
.Y(n_478)
);

BUFx6f_ASAP7_75t_SL g479 ( 
.A(n_239),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_294),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_257),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_295),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_260),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_299),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_302),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_320),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_266),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_R g488 ( 
.A(n_205),
.B(n_206),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_395),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_391),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_488),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_393),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_R g495 ( 
.A(n_461),
.B(n_205),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_396),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_394),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_405),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_259),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_410),
.B(n_362),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_462),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_397),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_448),
.B(n_280),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_423),
.B(n_424),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_399),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_399),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_411),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_259),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_402),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_412),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_416),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_418),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_464),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_R g517 ( 
.A(n_481),
.B(n_206),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_422),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_426),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_403),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_428),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_403),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_409),
.A2(n_215),
.B1(n_333),
.B2(n_356),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_450),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_430),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_438),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_463),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_407),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_442),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_463),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_433),
.B(n_466),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_459),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_404),
.A2(n_315),
.B1(n_226),
.B2(n_317),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_443),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_392),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_413),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_451),
.A2(n_323),
.B1(n_267),
.B2(n_382),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_466),
.B(n_355),
.Y(n_539)
);

BUFx8_ASAP7_75t_L g540 ( 
.A(n_479),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_459),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_465),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_465),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

AND2x6_ASAP7_75t_L g545 ( 
.A(n_420),
.B(n_214),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_468),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_447),
.Y(n_547)
);

AND3x2_ASAP7_75t_L g548 ( 
.A(n_421),
.B(n_398),
.C(n_389),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_453),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_468),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_456),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_413),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_415),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_457),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_483),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_415),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_455),
.B(n_213),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_469),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_427),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_469),
.B(n_355),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_427),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_470),
.B(n_213),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_429),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_429),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_400),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_432),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_470),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_441),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_492),
.B(n_460),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_489),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_506),
.B(n_487),
.C(n_439),
.Y(n_571)
);

NAND2x1p5_ASAP7_75t_L g572 ( 
.A(n_499),
.B(n_366),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_531),
.Y(n_573)
);

NOR3xp33_ASAP7_75t_L g574 ( 
.A(n_534),
.B(n_398),
.C(n_406),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_558),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_491),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_531),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_558),
.Y(n_579)
);

BUFx4f_ASAP7_75t_L g580 ( 
.A(n_545),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_493),
.Y(n_581)
);

NAND2x1p5_ASAP7_75t_L g582 ( 
.A(n_499),
.B(n_366),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_558),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_489),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_489),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_497),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_499),
.B(n_216),
.Y(n_587)
);

INVxp33_ASAP7_75t_L g588 ( 
.A(n_534),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_493),
.Y(n_589)
);

BUFx10_ASAP7_75t_L g590 ( 
.A(n_490),
.Y(n_590)
);

OA22x2_ASAP7_75t_L g591 ( 
.A1(n_506),
.A2(n_384),
.B1(n_350),
.B2(n_329),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_497),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_497),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_499),
.B(n_195),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_531),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_495),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_545),
.A2(n_451),
.B1(n_471),
.B2(n_434),
.Y(n_597)
);

AND2x2_ASAP7_75t_SL g598 ( 
.A(n_510),
.B(n_216),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_539),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_510),
.B(n_203),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_536),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_500),
.B(n_432),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_504),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_510),
.B(n_486),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_502),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_500),
.B(n_437),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_531),
.Y(n_607)
);

BUFx4f_ASAP7_75t_L g608 ( 
.A(n_545),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_523),
.B(n_401),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_504),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_510),
.B(n_232),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_532),
.B(n_240),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_502),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_531),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_492),
.B(n_431),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_494),
.Y(n_616)
);

AO21x1_ASAP7_75t_L g617 ( 
.A1(n_505),
.A2(n_340),
.B(n_339),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_524),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_507),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_532),
.B(n_435),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_504),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_507),
.B(n_292),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_545),
.B(n_247),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_531),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_560),
.B(n_437),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_545),
.A2(n_346),
.B1(n_341),
.B2(n_209),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_512),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_565),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_512),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_494),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_544),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_539),
.B(n_544),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_545),
.B(n_261),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_511),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_568),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_517),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_511),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_496),
.B(n_498),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_511),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_509),
.B(n_436),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_494),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_539),
.B(n_292),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_539),
.B(n_472),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_494),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_520),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_494),
.Y(n_646)
);

AO22x2_ASAP7_75t_L g647 ( 
.A1(n_538),
.A2(n_343),
.B1(n_208),
.B2(n_219),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_545),
.B(n_304),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_520),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_557),
.B(n_524),
.C(n_562),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_494),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_520),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_522),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_544),
.B(n_472),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_513),
.B(n_440),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_522),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_562),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_560),
.B(n_444),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_533),
.B(n_473),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_545),
.A2(n_408),
.B1(n_385),
.B2(n_335),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_503),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_522),
.Y(n_662)
);

AND2x2_ASAP7_75t_SL g663 ( 
.A(n_505),
.B(n_214),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_514),
.B(n_515),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_503),
.B(n_197),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_518),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_503),
.B(n_227),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_568),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_533),
.B(n_444),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_503),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_519),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_530),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_503),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_530),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_530),
.Y(n_675)
);

INVx6_ASAP7_75t_L g676 ( 
.A(n_503),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_557),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_508),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_508),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_508),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_508),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_559),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_521),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_541),
.B(n_445),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_548),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_508),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_528),
.Y(n_687)
);

OAI21xp33_ASAP7_75t_SL g688 ( 
.A1(n_567),
.A2(n_449),
.B(n_445),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_528),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_525),
.B(n_446),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_523),
.A2(n_345),
.B1(n_309),
.B2(n_306),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_559),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_538),
.A2(n_214),
.B1(n_297),
.B2(n_335),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_559),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_528),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_541),
.B(n_473),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_528),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_528),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_526),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_501),
.B(n_390),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_559),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_528),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_529),
.A2(n_458),
.B1(n_467),
.B2(n_476),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_542),
.B(n_486),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_559),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_559),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_527),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_542),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_543),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_535),
.B(n_547),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_527),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_549),
.B(n_425),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_551),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_554),
.B(n_479),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_543),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_516),
.B(n_474),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_SL g717 ( 
.A(n_540),
.B(n_414),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_546),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_546),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_552),
.Y(n_720)
);

O2A1O1Ixp5_ASAP7_75t_L g721 ( 
.A1(n_576),
.A2(n_581),
.B(n_589),
.C(n_578),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_632),
.B(n_550),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_618),
.B(n_555),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_618),
.B(n_417),
.Y(n_724)
);

BUFx8_ASAP7_75t_L g725 ( 
.A(n_685),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_657),
.B(n_552),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_677),
.B(n_217),
.Y(n_727)
);

BUFx8_ASAP7_75t_L g728 ( 
.A(n_685),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_677),
.B(n_217),
.Y(n_729)
);

BUFx4f_ASAP7_75t_L g730 ( 
.A(n_700),
.Y(n_730)
);

NOR3x1_ASAP7_75t_L g731 ( 
.A(n_571),
.B(n_475),
.C(n_474),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_663),
.B(n_552),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_718),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_598),
.B(n_214),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_663),
.B(n_552),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_598),
.B(n_580),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_612),
.B(n_556),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_576),
.B(n_556),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_716),
.B(n_650),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_620),
.B(n_596),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_578),
.B(n_556),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_716),
.B(n_218),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_594),
.B(n_218),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_718),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_591),
.A2(n_214),
.B1(n_297),
.B2(n_385),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_581),
.B(n_589),
.Y(n_746)
);

INVx8_ASAP7_75t_L g747 ( 
.A(n_587),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_580),
.B(n_297),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_605),
.B(n_556),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_605),
.B(n_242),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_580),
.B(n_297),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_613),
.B(n_253),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_613),
.B(n_262),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_632),
.A2(n_419),
.B1(n_228),
.B2(n_351),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_600),
.B(n_220),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_599),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_671),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_632),
.A2(n_353),
.B1(n_228),
.B2(n_229),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_619),
.B(n_269),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_599),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_720),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_627),
.B(n_629),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_597),
.B(n_271),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_596),
.B(n_550),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_591),
.A2(n_335),
.B1(n_385),
.B2(n_297),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_608),
.A2(n_527),
.B(n_537),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_575),
.B(n_273),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_635),
.B(n_567),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_608),
.B(n_335),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_579),
.B(n_279),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_636),
.B(n_540),
.Y(n_771)
);

NAND2x1p5_ASAP7_75t_L g772 ( 
.A(n_608),
.B(n_281),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_604),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_583),
.B(n_289),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_625),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_604),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_604),
.B(n_335),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_719),
.B(n_293),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_625),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_669),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_708),
.B(n_303),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_611),
.B(n_623),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_569),
.B(n_220),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_709),
.B(n_313),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_691),
.B(n_631),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_720),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_658),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_671),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_SL g789 ( 
.A(n_588),
.B(n_347),
.C(n_236),
.Y(n_789)
);

OAI221xp5_ASAP7_75t_L g790 ( 
.A1(n_693),
.A2(n_314),
.B1(n_380),
.B2(n_379),
.C(n_375),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_658),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_715),
.B(n_324),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_643),
.B(n_475),
.Y(n_793)
);

NOR2x1p5_ASAP7_75t_L g794 ( 
.A(n_636),
.B(n_207),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_669),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_602),
.B(n_354),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_668),
.B(n_477),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_615),
.B(n_229),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_587),
.B(n_326),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_643),
.B(n_477),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_602),
.B(n_606),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_643),
.B(n_230),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_633),
.A2(n_648),
.B(n_665),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_630),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_606),
.B(n_222),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_570),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_659),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_684),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_654),
.B(n_480),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_587),
.A2(n_230),
.B1(n_234),
.B2(n_270),
.Y(n_810)
);

NOR2x1p5_ASAP7_75t_L g811 ( 
.A(n_700),
.B(n_207),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_572),
.B(n_383),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_572),
.B(n_387),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_582),
.B(n_388),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_684),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_630),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_582),
.B(n_537),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_582),
.B(n_385),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_570),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_626),
.B(n_385),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_660),
.B(n_537),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_680),
.B(n_553),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_591),
.A2(n_334),
.B1(n_386),
.B2(n_234),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_617),
.A2(n_326),
.B1(n_331),
.B2(n_338),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_654),
.B(n_714),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_659),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_654),
.B(n_617),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_584),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_680),
.B(n_553),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_638),
.B(n_270),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_696),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_696),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_664),
.B(n_311),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_584),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_697),
.B(n_553),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_696),
.B(n_311),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_697),
.B(n_561),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_704),
.B(n_318),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_704),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_682),
.B(n_326),
.Y(n_841)
);

NOR3x1_ASAP7_75t_L g842 ( 
.A(n_690),
.B(n_485),
.C(n_484),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_682),
.B(n_326),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_641),
.B(n_561),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_683),
.B(n_222),
.Y(n_845)
);

AO22x1_ASAP7_75t_L g846 ( 
.A1(n_574),
.A2(n_212),
.B1(n_211),
.B2(n_225),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_647),
.A2(n_326),
.B1(n_331),
.B2(n_338),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_704),
.B(n_318),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_661),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_SL g850 ( 
.A(n_713),
.B(n_699),
.Y(n_850)
);

NAND3xp33_ASAP7_75t_L g851 ( 
.A(n_710),
.B(n_540),
.C(n_274),
.Y(n_851)
);

NOR2xp67_ASAP7_75t_L g852 ( 
.A(n_703),
.B(n_712),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_679),
.B(n_319),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_587),
.A2(n_386),
.B1(n_351),
.B2(n_332),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_641),
.B(n_678),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_667),
.A2(n_527),
.B(n_564),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_585),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_587),
.B(n_480),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_639),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_641),
.B(n_678),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_692),
.B(n_694),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_678),
.B(n_561),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_695),
.B(n_573),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_686),
.B(n_687),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_695),
.B(n_563),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_647),
.A2(n_326),
.B1(n_331),
.B2(n_211),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_695),
.B(n_563),
.Y(n_867)
);

NOR3xp33_ASAP7_75t_L g868 ( 
.A(n_640),
.B(n_484),
.C(n_482),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_585),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_573),
.B(n_563),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_647),
.A2(n_326),
.B1(n_331),
.B2(n_212),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_573),
.B(n_564),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_649),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_590),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_595),
.B(n_564),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_649),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_655),
.B(n_485),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_656),
.B(n_672),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_587),
.B(n_449),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_656),
.B(n_319),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_590),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_672),
.B(n_332),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_666),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_661),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_642),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_586),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_647),
.A2(n_331),
.B1(n_225),
.B2(n_344),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_776),
.B(n_642),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_806),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_773),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_757),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_806),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_723),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_SL g894 ( 
.A(n_736),
.B(n_699),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_SL g895 ( 
.A(n_798),
.B(n_609),
.C(n_601),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_722),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_817),
.A2(n_782),
.B(n_803),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_768),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_722),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_776),
.B(n_642),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_797),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_885),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_849),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_773),
.B(n_807),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_819),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_726),
.B(n_642),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_807),
.Y(n_907)
);

OAI21xp33_ASAP7_75t_SL g908 ( 
.A1(n_736),
.A2(n_675),
.B(n_674),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_739),
.B(n_666),
.Y(n_909)
);

INVxp67_ASAP7_75t_SL g910 ( 
.A(n_849),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_801),
.B(n_858),
.Y(n_911)
);

BUFx4f_ASAP7_75t_L g912 ( 
.A(n_874),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_SL g913 ( 
.A(n_798),
.B(n_609),
.C(n_628),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_743),
.B(n_642),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_724),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_743),
.B(n_642),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_819),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_733),
.Y(n_918)
);

BUFx10_ASAP7_75t_L g919 ( 
.A(n_788),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_R g920 ( 
.A(n_850),
.B(n_717),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_828),
.A2(n_688),
.B(n_674),
.C(n_322),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_744),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_730),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_764),
.B(n_452),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_756),
.B(n_673),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_SL g926 ( 
.A(n_789),
.B(n_325),
.C(n_236),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_740),
.B(n_673),
.Y(n_927)
);

NOR2x1_ASAP7_75t_L g928 ( 
.A(n_851),
.B(n_877),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_761),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_R g930 ( 
.A(n_881),
.B(n_540),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_825),
.A2(n_622),
.B1(n_331),
.B2(n_592),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_829),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_829),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_775),
.B(n_310),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_756),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_760),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_884),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_755),
.B(n_586),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_835),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_805),
.B(n_452),
.Y(n_940)
);

AND2x6_ASAP7_75t_SL g941 ( 
.A(n_831),
.B(n_310),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_755),
.B(n_592),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_779),
.B(n_312),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_760),
.B(n_681),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_725),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_823),
.B(n_681),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_835),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_761),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_857),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_884),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_730),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_L g952 ( 
.A(n_885),
.B(n_622),
.Y(n_952)
);

BUFx8_ASAP7_75t_L g953 ( 
.A(n_883),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_SL g954 ( 
.A(n_783),
.B(n_321),
.C(n_312),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_858),
.B(n_630),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_R g956 ( 
.A(n_725),
.B(n_334),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_737),
.B(n_593),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_786),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_885),
.B(n_630),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_879),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_857),
.Y(n_961)
);

NOR3xp33_ASAP7_75t_L g962 ( 
.A(n_831),
.B(n_381),
.C(n_353),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_746),
.B(n_787),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_SL g964 ( 
.A(n_783),
.B(n_754),
.C(n_834),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_791),
.B(n_593),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_727),
.B(n_321),
.Y(n_966)
);

BUFx4f_ASAP7_75t_L g967 ( 
.A(n_877),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_869),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_828),
.B(n_603),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_827),
.B(n_689),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_869),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_859),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_780),
.B(n_603),
.Y(n_973)
);

AND3x1_ASAP7_75t_SL g974 ( 
.A(n_794),
.B(n_811),
.C(n_790),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_795),
.B(n_610),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_727),
.B(n_322),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_808),
.B(n_610),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_815),
.B(n_621),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_728),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_762),
.B(n_621),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_825),
.A2(n_866),
.B1(n_871),
.B2(n_847),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_847),
.A2(n_871),
.B1(n_866),
.B2(n_887),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_873),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_729),
.B(n_634),
.Y(n_984)
);

CKINVDCx14_ASAP7_75t_R g985 ( 
.A(n_845),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_729),
.B(n_689),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_SL g987 ( 
.A(n_834),
.B(n_325),
.C(n_328),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_742),
.B(n_328),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_742),
.B(n_616),
.Y(n_989)
);

BUFx4f_ASAP7_75t_L g990 ( 
.A(n_877),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_728),
.B(n_381),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_SL g992 ( 
.A(n_852),
.B(n_479),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_SL g993 ( 
.A(n_785),
.B(n_336),
.Y(n_993)
);

INVx5_ASAP7_75t_L g994 ( 
.A(n_747),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_833),
.B(n_634),
.Y(n_995)
);

NOR3xp33_ASAP7_75t_SL g996 ( 
.A(n_785),
.B(n_349),
.C(n_378),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_809),
.B(n_336),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_886),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_R g999 ( 
.A(n_747),
.B(n_342),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_876),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_809),
.B(n_342),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_840),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_886),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_832),
.B(n_637),
.Y(n_1004)
);

INVxp33_ASAP7_75t_SL g1005 ( 
.A(n_842),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_793),
.B(n_800),
.Y(n_1006)
);

INVx5_ASAP7_75t_L g1007 ( 
.A(n_747),
.Y(n_1007)
);

AND3x1_ASAP7_75t_SL g1008 ( 
.A(n_846),
.B(n_352),
.C(n_378),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_793),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_721),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_885),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_868),
.Y(n_1012)
);

OR2x6_ASAP7_75t_L g1013 ( 
.A(n_771),
.B(n_692),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_816),
.Y(n_1014)
);

BUFx10_ASAP7_75t_L g1015 ( 
.A(n_837),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_804),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_800),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_887),
.A2(n_622),
.B1(n_331),
.B2(n_652),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_758),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_738),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_879),
.B(n_694),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_837),
.B(n_344),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_763),
.B(n_637),
.Y(n_1023)
);

CKINVDCx8_ASAP7_75t_R g1024 ( 
.A(n_839),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_826),
.B(n_616),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_SL g1026 ( 
.A(n_839),
.B(n_347),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_822),
.Y(n_1027)
);

AND3x2_ASAP7_75t_SL g1028 ( 
.A(n_745),
.B(n_348),
.C(n_349),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_796),
.B(n_348),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_816),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_880),
.B(n_645),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_759),
.Y(n_1032)
);

AOI211xp5_ASAP7_75t_L g1033 ( 
.A1(n_824),
.A2(n_376),
.B(n_382),
.C(n_352),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_741),
.Y(n_1034)
);

INVx5_ASAP7_75t_L g1035 ( 
.A(n_799),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_732),
.B(n_630),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_863),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_830),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_848),
.B(n_376),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_731),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_749),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_848),
.B(n_377),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_802),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_735),
.B(n_646),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_836),
.Y(n_1045)
);

AOI22x1_ASAP7_75t_L g1046 ( 
.A1(n_772),
.A2(n_701),
.B1(n_645),
.B2(n_652),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_838),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_812),
.B(n_646),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_781),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_813),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_814),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_864),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_864),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_844),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_870),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_855),
.Y(n_1056)
);

BUFx12f_ASAP7_75t_L g1057 ( 
.A(n_772),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_860),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_862),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_818),
.A2(n_670),
.B(n_644),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_872),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_802),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_767),
.B(n_377),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_865),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_880),
.B(n_882),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_SL g1066 ( 
.A(n_777),
.B(n_276),
.C(n_282),
.Y(n_1066)
);

AND2x6_ASAP7_75t_L g1067 ( 
.A(n_821),
.B(n_701),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_861),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_734),
.B(n_676),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_882),
.B(n_286),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_861),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_745),
.B(n_300),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_750),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_765),
.B(n_853),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_878),
.Y(n_1075)
);

AO31x2_ASAP7_75t_L g1076 ( 
.A1(n_921),
.A2(n_1010),
.A3(n_897),
.B(n_969),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_918),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1075),
.B(n_765),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_922),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_914),
.A2(n_734),
.B(n_818),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_902),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_981),
.B(n_1065),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_891),
.Y(n_1083)
);

NOR2xp67_ASAP7_75t_L g1084 ( 
.A(n_891),
.B(n_770),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1074),
.B(n_752),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_898),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_889),
.Y(n_1087)
);

NOR3xp33_ASAP7_75t_L g1088 ( 
.A(n_964),
.B(n_792),
.C(n_784),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_916),
.A2(n_769),
.B(n_748),
.Y(n_1089)
);

BUFx8_ASAP7_75t_SL g1090 ( 
.A(n_945),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_906),
.A2(n_748),
.B(n_751),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_902),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1046),
.A2(n_875),
.B(n_867),
.Y(n_1093)
);

AO31x2_ASAP7_75t_L g1094 ( 
.A1(n_921),
.A2(n_878),
.A3(n_753),
.B(n_778),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1060),
.A2(n_892),
.B(n_889),
.Y(n_1095)
);

BUFx8_ASAP7_75t_L g1096 ( 
.A(n_979),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_963),
.B(n_853),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1035),
.A2(n_751),
.B(n_769),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_892),
.A2(n_843),
.B(n_841),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_898),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_902),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_905),
.A2(n_843),
.B(n_841),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_SL g1103 ( 
.A(n_994),
.B(n_820),
.Y(n_1103)
);

AO21x1_ASAP7_75t_L g1104 ( 
.A1(n_989),
.A2(n_774),
.B(n_777),
.Y(n_1104)
);

INVx5_ASAP7_75t_L g1105 ( 
.A(n_902),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_905),
.A2(n_766),
.B(n_856),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_986),
.B(n_810),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_986),
.B(n_854),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_917),
.A2(n_933),
.B(n_932),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_1011),
.Y(n_1110)
);

O2A1O1Ixp5_ASAP7_75t_L g1111 ( 
.A1(n_989),
.A2(n_820),
.B(n_662),
.C(n_653),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1035),
.A2(n_644),
.B(n_616),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_908),
.A2(n_653),
.B(n_662),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_924),
.B(n_1052),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_1025),
.A2(n_670),
.A3(n_644),
.B(n_698),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1036),
.A2(n_698),
.B(n_670),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_972),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_993),
.B(n_363),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_932),
.A2(n_711),
.B(n_707),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_893),
.B(n_370),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_933),
.A2(n_711),
.B(n_707),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1035),
.A2(n_1023),
.B(n_1031),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1053),
.B(n_622),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_983),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_1011),
.Y(n_1125)
);

AOI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1044),
.A2(n_1048),
.B(n_942),
.Y(n_1126)
);

NOR2x1_ASAP7_75t_SL g1127 ( 
.A(n_994),
.B(n_646),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_1011),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_939),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_939),
.A2(n_711),
.B(n_707),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_940),
.B(n_622),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1044),
.A2(n_566),
.B(n_527),
.Y(n_1132)
);

AOI221x1_ASAP7_75t_L g1133 ( 
.A1(n_894),
.A2(n_706),
.B1(n_705),
.B2(n_702),
.C(n_651),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_981),
.A2(n_676),
.B1(n_577),
.B2(n_624),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1035),
.A2(n_624),
.B(n_577),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_982),
.B(n_646),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1032),
.B(n_577),
.Y(n_1137)
);

NOR2x1_ASAP7_75t_SL g1138 ( 
.A(n_994),
.B(n_646),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1011),
.Y(n_1139)
);

HB1xp67_ASAP7_75t_L g1140 ( 
.A(n_901),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_911),
.A2(n_527),
.B(n_371),
.Y(n_1141)
);

AO21x1_ASAP7_75t_L g1142 ( 
.A1(n_894),
.A2(n_331),
.B(n_23),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_966),
.B(n_23),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1062),
.A2(n_676),
.B1(n_577),
.B2(n_624),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1048),
.A2(n_676),
.B(n_577),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1049),
.B(n_624),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_SL g1147 ( 
.A1(n_982),
.A2(n_72),
.B(n_194),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1006),
.B(n_624),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1073),
.B(n_614),
.Y(n_1149)
);

AOI221x1_ASAP7_75t_L g1150 ( 
.A1(n_962),
.A2(n_987),
.B1(n_954),
.B2(n_927),
.C(n_938),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_947),
.A2(n_614),
.B(n_607),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1040),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_911),
.A2(n_614),
.B(n_607),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_947),
.A2(n_614),
.B(n_607),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1025),
.A2(n_706),
.A3(n_705),
.B(n_702),
.Y(n_1155)
);

OR2x6_ASAP7_75t_L g1156 ( 
.A(n_1006),
.B(n_702),
.Y(n_1156)
);

AO21x1_ASAP7_75t_L g1157 ( 
.A1(n_1033),
.A2(n_25),
.B(n_26),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_957),
.A2(n_614),
.B(n_607),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1070),
.B(n_607),
.Y(n_1159)
);

INVx5_ASAP7_75t_L g1160 ( 
.A(n_994),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1040),
.Y(n_1161)
);

AO21x1_ASAP7_75t_L g1162 ( 
.A1(n_984),
.A2(n_27),
.B(n_31),
.Y(n_1162)
);

AOI21x1_ASAP7_75t_SL g1163 ( 
.A1(n_1043),
.A2(n_706),
.B(n_705),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_888),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_888),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_L g1166 ( 
.A1(n_904),
.A2(n_702),
.B(n_651),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1072),
.A2(n_702),
.B(n_651),
.C(n_706),
.Y(n_1167)
);

AO32x2_ASAP7_75t_L g1168 ( 
.A1(n_1068),
.A2(n_31),
.A3(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_988),
.B(n_34),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1045),
.B(n_651),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1000),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1047),
.B(n_651),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_888),
.Y(n_1173)
);

OA22x2_ASAP7_75t_L g1174 ( 
.A1(n_1019),
.A2(n_1012),
.B1(n_1009),
.B2(n_1043),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_927),
.B(n_706),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1050),
.B(n_705),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_949),
.A2(n_128),
.B(n_190),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_909),
.A2(n_39),
.B(n_40),
.C(n_43),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_929),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1020),
.A2(n_40),
.A3(n_44),
.B(n_45),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_948),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1051),
.B(n_44),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1007),
.A2(n_527),
.B1(n_83),
.B2(n_84),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_980),
.A2(n_134),
.B(n_187),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_952),
.A2(n_125),
.B(n_179),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_919),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_949),
.A2(n_188),
.B(n_178),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1034),
.A2(n_46),
.A3(n_47),
.B(n_48),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_952),
.A2(n_1016),
.B(n_1038),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1022),
.B(n_47),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1068),
.A2(n_48),
.A3(n_49),
.B(n_51),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_961),
.A2(n_177),
.B(n_175),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_961),
.A2(n_174),
.B(n_121),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1039),
.B(n_51),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_968),
.A2(n_97),
.B(n_90),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1042),
.B(n_53),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1007),
.A2(n_89),
.B1(n_85),
.B2(n_80),
.Y(n_1197)
);

INVx4_ASAP7_75t_L g1198 ( 
.A(n_925),
.Y(n_1198)
);

CKINVDCx11_ASAP7_75t_R g1199 ( 
.A(n_919),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_915),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1027),
.B(n_53),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_958),
.Y(n_1202)
);

AOI31xp67_ASAP7_75t_L g1203 ( 
.A1(n_1055),
.A2(n_54),
.A3(n_59),
.B(n_60),
.Y(n_1203)
);

NOR3xp33_ASAP7_75t_L g1204 ( 
.A(n_895),
.B(n_61),
.C(n_65),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1027),
.A2(n_61),
.A3(n_65),
.B(n_66),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1038),
.B(n_67),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_909),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1054),
.A2(n_1059),
.B(n_1064),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_968),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_900),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_903),
.A2(n_910),
.B(n_937),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1041),
.B(n_1002),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1055),
.A2(n_1061),
.B(n_931),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_904),
.A2(n_1061),
.B(n_959),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1041),
.B(n_935),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_971),
.A2(n_998),
.B(n_959),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1007),
.A2(n_935),
.B1(n_1069),
.B2(n_1024),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1006),
.B(n_936),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_931),
.A2(n_995),
.B(n_1067),
.Y(n_1219)
);

BUFx12f_ASAP7_75t_L g1220 ( 
.A(n_953),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1018),
.A2(n_1003),
.B(n_971),
.Y(n_1221)
);

AOI21x1_ASAP7_75t_L g1222 ( 
.A1(n_973),
.A2(n_975),
.B(n_977),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_998),
.A2(n_978),
.B(n_955),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_955),
.A2(n_950),
.B(n_1004),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_936),
.B(n_896),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_925),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_965),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_950),
.A2(n_907),
.B(n_890),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_907),
.A2(n_890),
.B(n_960),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_976),
.B(n_1029),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1007),
.A2(n_1069),
.B1(n_1019),
.B2(n_960),
.Y(n_1231)
);

INVx3_ASAP7_75t_SL g1232 ( 
.A(n_923),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1160),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1100),
.Y(n_1234)
);

INVx4_ASAP7_75t_L g1235 ( 
.A(n_1105),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1118),
.A2(n_985),
.B1(n_1005),
.B2(n_951),
.Y(n_1236)
);

AOI221xp5_ASAP7_75t_L g1237 ( 
.A1(n_1118),
.A2(n_913),
.B1(n_1026),
.B2(n_996),
.C(n_920),
.Y(n_1237)
);

INVx6_ASAP7_75t_L g1238 ( 
.A(n_1186),
.Y(n_1238)
);

AND2x6_ASAP7_75t_L g1239 ( 
.A(n_1101),
.B(n_1071),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1145),
.A2(n_1018),
.B(n_928),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1204),
.A2(n_967),
.B1(n_990),
.B2(n_1015),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1122),
.A2(n_1080),
.B(n_1098),
.Y(n_1242)
);

OR2x6_ASAP7_75t_L g1243 ( 
.A(n_1231),
.B(n_1189),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1151),
.A2(n_1067),
.B(n_899),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1086),
.Y(n_1245)
);

AO21x2_ASAP7_75t_L g1246 ( 
.A1(n_1122),
.A2(n_1066),
.B(n_970),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1100),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1114),
.B(n_1015),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1140),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1208),
.B(n_926),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1107),
.A2(n_1067),
.B(n_946),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1154),
.A2(n_1067),
.B(n_1063),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1230),
.B(n_985),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1218),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1166),
.A2(n_1067),
.B(n_1001),
.Y(n_1255)
);

OAI21xp33_ASAP7_75t_L g1256 ( 
.A1(n_1120),
.A2(n_920),
.B(n_1005),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1077),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1095),
.A2(n_997),
.B(n_943),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1079),
.Y(n_1259)
);

AOI21xp33_ASAP7_75t_L g1260 ( 
.A1(n_1108),
.A2(n_934),
.B(n_967),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1097),
.B(n_1017),
.Y(n_1261)
);

CKINVDCx16_ASAP7_75t_R g1262 ( 
.A(n_1186),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1227),
.B(n_944),
.Y(n_1263)
);

INVx5_ASAP7_75t_L g1264 ( 
.A(n_1101),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1199),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1127),
.A2(n_900),
.B(n_1014),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1085),
.B(n_990),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1093),
.A2(n_1058),
.B(n_1037),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1083),
.Y(n_1269)
);

AOI221xp5_ASAP7_75t_L g1270 ( 
.A1(n_1204),
.A2(n_991),
.B1(n_956),
.B2(n_992),
.C(n_941),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1140),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1200),
.B(n_1013),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1105),
.B(n_1030),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1199),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_SL g1275 ( 
.A1(n_1147),
.A2(n_1057),
.B(n_1013),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1104),
.A2(n_1028),
.A3(n_1069),
.B(n_1008),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1169),
.B(n_999),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1133),
.A2(n_946),
.B(n_970),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1082),
.A2(n_946),
.B(n_970),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1167),
.A2(n_1219),
.B(n_1089),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1163),
.A2(n_1056),
.B(n_1037),
.Y(n_1281)
);

BUFx2_ASAP7_75t_R g1282 ( 
.A(n_1090),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1083),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1089),
.A2(n_1056),
.B(n_1058),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1167),
.A2(n_1021),
.B(n_925),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1143),
.B(n_1190),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1117),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_SL g1288 ( 
.A1(n_1185),
.A2(n_1057),
.B(n_1013),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1091),
.A2(n_1021),
.B(n_944),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1163),
.A2(n_1056),
.B(n_1037),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1124),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1164),
.B(n_944),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1129),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1194),
.B(n_1056),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1084),
.A2(n_974),
.B1(n_912),
.B2(n_1021),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1228),
.A2(n_1071),
.B(n_912),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1171),
.Y(n_1297)
);

AOI221xp5_ASAP7_75t_L g1298 ( 
.A1(n_1196),
.A2(n_1178),
.B1(n_1157),
.B2(n_1207),
.C(n_1161),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1179),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_SL g1300 ( 
.A1(n_1088),
.A2(n_1071),
.B(n_953),
.C(n_930),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1109),
.A2(n_1071),
.B(n_953),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1078),
.A2(n_930),
.B1(n_956),
.B2(n_991),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1129),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1212),
.A2(n_1189),
.B1(n_1215),
.B2(n_1198),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1174),
.A2(n_1152),
.B1(n_1220),
.B2(n_1182),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1229),
.A2(n_1113),
.B(n_1106),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1209),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1090),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1152),
.B(n_1161),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1209),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1214),
.A2(n_1216),
.B(n_1223),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1181),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1165),
.B(n_1173),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1198),
.A2(n_1226),
.B1(n_1217),
.B2(n_1213),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1174),
.A2(n_1088),
.B1(n_1225),
.B2(n_1232),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1214),
.A2(n_1195),
.B(n_1192),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1164),
.B(n_1210),
.Y(n_1317)
);

AND2x6_ASAP7_75t_L g1318 ( 
.A(n_1101),
.B(n_1165),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1202),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1150),
.B(n_1149),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1221),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1221),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1091),
.A2(n_1123),
.B(n_1159),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1225),
.A2(n_1232),
.B1(n_1173),
.B2(n_1131),
.Y(n_1324)
);

INVx3_ASAP7_75t_SL g1325 ( 
.A(n_1156),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1226),
.A2(n_1144),
.B1(n_1175),
.B2(n_1156),
.Y(n_1326)
);

AO21x2_ASAP7_75t_L g1327 ( 
.A1(n_1136),
.A2(n_1126),
.B(n_1116),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1177),
.A2(n_1193),
.B(n_1187),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1096),
.Y(n_1329)
);

CKINVDCx16_ASAP7_75t_R g1330 ( 
.A(n_1220),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1162),
.A2(n_1142),
.B1(n_1201),
.B2(n_1206),
.Y(n_1331)
);

NAND2x1_ASAP7_75t_L g1332 ( 
.A(n_1128),
.B(n_1101),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1176),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1096),
.A2(n_1160),
.B1(n_1197),
.B2(n_1141),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1184),
.A2(n_1185),
.B1(n_1136),
.B2(n_1183),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1137),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1221),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1164),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1158),
.A2(n_1153),
.B(n_1135),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1111),
.A2(n_1211),
.B(n_1224),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1148),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1158),
.A2(n_1153),
.B(n_1135),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1119),
.A2(n_1130),
.B(n_1121),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1111),
.A2(n_1211),
.B(n_1102),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1099),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1156),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1076),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1210),
.B(n_1148),
.Y(n_1348)
);

OAI222xp33_ASAP7_75t_L g1349 ( 
.A1(n_1103),
.A2(n_1184),
.B1(n_1178),
.B2(n_1172),
.C1(n_1170),
.C2(n_1146),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1210),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1148),
.B(n_1076),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_SL g1352 ( 
.A1(n_1134),
.A2(n_1168),
.B(n_1132),
.C(n_1092),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_SL g1353 ( 
.A(n_1128),
.B(n_1105),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1105),
.B(n_1160),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1081),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1168),
.A2(n_1081),
.B1(n_1092),
.B2(n_1139),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1112),
.A2(n_1222),
.B(n_1139),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1110),
.A2(n_1125),
.B(n_1203),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1168),
.A2(n_1110),
.B(n_1125),
.C(n_1094),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1155),
.A2(n_1076),
.B(n_1115),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1076),
.B(n_1094),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1155),
.A2(n_1115),
.B(n_1094),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1155),
.A2(n_1115),
.B(n_1094),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1138),
.A2(n_1115),
.B(n_1155),
.Y(n_1364)
);

INVxp67_ASAP7_75t_SL g1365 ( 
.A(n_1168),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1205),
.A2(n_1191),
.B(n_1180),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1205),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1191),
.A2(n_1180),
.B(n_1188),
.C(n_1205),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1191),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1205),
.A2(n_1191),
.B(n_1180),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1180),
.A2(n_993),
.B1(n_1118),
.B2(n_920),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1188),
.B(n_1164),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1188),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1188),
.A2(n_1145),
.B(n_1151),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1087),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1208),
.B(n_1085),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1114),
.B(n_1097),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1101),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1083),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1077),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_SL g1381 ( 
.A1(n_1178),
.A2(n_1082),
.B(n_964),
.C(n_921),
.Y(n_1381)
);

AO31x2_ASAP7_75t_L g1382 ( 
.A1(n_1104),
.A2(n_1133),
.A3(n_1167),
.B(n_1142),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1231),
.B(n_1189),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1164),
.B(n_1210),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1087),
.Y(n_1385)
);

NOR2x1_ASAP7_75t_SL g1386 ( 
.A(n_1160),
.B(n_1105),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1086),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1160),
.Y(n_1388)
);

NAND2xp33_ASAP7_75t_SL g1389 ( 
.A(n_1236),
.B(n_1325),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1277),
.B(n_1253),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1257),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1377),
.B(n_1376),
.Y(n_1392)
);

CKINVDCx16_ASAP7_75t_R g1393 ( 
.A(n_1262),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1376),
.B(n_1261),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1259),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1315),
.A2(n_1248),
.B1(n_1286),
.B2(n_1237),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1298),
.A2(n_1371),
.B1(n_1250),
.B2(n_1270),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1271),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_1241),
.B(n_1260),
.C(n_1250),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1256),
.A2(n_1267),
.B1(n_1241),
.B2(n_1302),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1381),
.A2(n_1267),
.B(n_1300),
.C(n_1349),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1249),
.B(n_1309),
.Y(n_1402)
);

NAND2xp33_ASAP7_75t_L g1403 ( 
.A(n_1338),
.B(n_1254),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1264),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1333),
.B(n_1263),
.Y(n_1405)
);

AO21x2_ASAP7_75t_L g1406 ( 
.A1(n_1344),
.A2(n_1340),
.B(n_1242),
.Y(n_1406)
);

INVx4_ASAP7_75t_L g1407 ( 
.A(n_1235),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1381),
.A2(n_1300),
.B(n_1320),
.C(n_1234),
.Y(n_1408)
);

BUFx4f_ASAP7_75t_L g1409 ( 
.A(n_1238),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1348),
.B(n_1292),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1295),
.A2(n_1272),
.B1(n_1324),
.B2(n_1305),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1348),
.B(n_1292),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1365),
.A2(n_1280),
.B1(n_1314),
.B2(n_1379),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1294),
.B(n_1247),
.Y(n_1414)
);

AOI221xp5_ASAP7_75t_L g1415 ( 
.A1(n_1331),
.A2(n_1352),
.B1(n_1335),
.B2(n_1368),
.C(n_1380),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1264),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1280),
.A2(n_1283),
.B1(n_1269),
.B2(n_1379),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1292),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1317),
.B(n_1384),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1247),
.B(n_1336),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1331),
.A2(n_1334),
.B1(n_1335),
.B2(n_1383),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1351),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1372),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1245),
.B(n_1387),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1269),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1243),
.A2(n_1383),
.B1(n_1291),
.B2(n_1287),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1297),
.A2(n_1319),
.B1(n_1312),
.B2(n_1299),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1328),
.A2(n_1316),
.B(n_1268),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1338),
.A2(n_1341),
.B1(n_1325),
.B2(n_1383),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1317),
.B(n_1384),
.Y(n_1430)
);

O2A1O1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1288),
.A2(n_1304),
.B(n_1326),
.C(n_1275),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1283),
.B(n_1350),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1243),
.A2(n_1383),
.B1(n_1369),
.B2(n_1279),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1293),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1317),
.B(n_1384),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1243),
.A2(n_1387),
.B1(n_1245),
.B2(n_1346),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1243),
.A2(n_1251),
.B1(n_1372),
.B2(n_1373),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1313),
.B(n_1235),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1303),
.B(n_1307),
.Y(n_1439)
);

AO31x2_ASAP7_75t_L g1440 ( 
.A1(n_1359),
.A2(n_1367),
.A3(n_1347),
.B(n_1361),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1310),
.B(n_1375),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1276),
.B(n_1355),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1372),
.A2(n_1246),
.B1(n_1289),
.B2(n_1238),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1375),
.B(n_1385),
.Y(n_1444)
);

OAI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1323),
.A2(n_1329),
.B1(n_1238),
.B2(n_1284),
.C(n_1265),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1385),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1276),
.B(n_1258),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1353),
.A2(n_1330),
.B1(n_1274),
.B2(n_1265),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1276),
.B(n_1258),
.Y(n_1449)
);

AO31x2_ASAP7_75t_L g1450 ( 
.A1(n_1359),
.A2(n_1347),
.A3(n_1345),
.B(n_1321),
.Y(n_1450)
);

NAND2xp33_ASAP7_75t_SL g1451 ( 
.A(n_1308),
.B(n_1274),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1308),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1233),
.Y(n_1453)
);

CKINVDCx14_ASAP7_75t_R g1454 ( 
.A(n_1282),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1255),
.A2(n_1252),
.B(n_1240),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1352),
.A2(n_1358),
.B(n_1246),
.C(n_1327),
.Y(n_1456)
);

NAND3xp33_ASAP7_75t_L g1457 ( 
.A(n_1356),
.B(n_1285),
.C(n_1345),
.Y(n_1457)
);

INVx3_ASAP7_75t_SL g1458 ( 
.A(n_1378),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1366),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1327),
.A2(n_1285),
.B1(n_1356),
.B2(n_1366),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1378),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1378),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1370),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1266),
.A2(n_1273),
.B1(n_1264),
.B2(n_1278),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1339),
.A2(n_1342),
.B(n_1285),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1328),
.A2(n_1316),
.B(n_1268),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1273),
.A2(n_1264),
.B1(n_1278),
.B2(n_1354),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1378),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1370),
.A2(n_1322),
.B1(n_1321),
.B2(n_1337),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1322),
.A2(n_1337),
.B1(n_1255),
.B2(n_1278),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1354),
.Y(n_1471)
);

OAI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1332),
.A2(n_1233),
.B1(n_1388),
.B2(n_1252),
.C(n_1240),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1318),
.A2(n_1239),
.B1(n_1364),
.B2(n_1363),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1239),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1239),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1318),
.Y(n_1476)
);

AOI222xp33_ASAP7_75t_L g1477 ( 
.A1(n_1318),
.A2(n_1239),
.B1(n_1386),
.B2(n_1388),
.C1(n_1233),
.C2(n_1363),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1239),
.A2(n_1318),
.B1(n_1388),
.B2(n_1296),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1362),
.A2(n_1360),
.B1(n_1301),
.B2(n_1296),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1244),
.A2(n_1357),
.B(n_1342),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1301),
.A2(n_1281),
.B1(n_1290),
.B2(n_1382),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1281),
.Y(n_1482)
);

AO32x2_ASAP7_75t_L g1483 ( 
.A1(n_1382),
.A2(n_1362),
.A3(n_1360),
.B1(n_1374),
.B2(n_1311),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1290),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1374),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1244),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1382),
.A2(n_1339),
.B1(n_1306),
.B2(n_1311),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1306),
.A2(n_964),
.B1(n_1118),
.B2(n_895),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1343),
.A2(n_964),
.B(n_1065),
.C(n_1118),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1382),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1343),
.A2(n_1242),
.B(n_1122),
.Y(n_1491)
);

AOI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1381),
.A2(n_588),
.B1(n_691),
.B2(n_964),
.C(n_1118),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1377),
.B(n_740),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1298),
.A2(n_964),
.B1(n_1204),
.B2(n_993),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1365),
.A2(n_993),
.B1(n_1118),
.B2(n_1074),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1234),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1377),
.A2(n_993),
.B1(n_1207),
.B2(n_1065),
.Y(n_1497)
);

AO21x2_ASAP7_75t_L g1498 ( 
.A1(n_1344),
.A2(n_1340),
.B(n_1242),
.Y(n_1498)
);

NAND3xp33_ASAP7_75t_SL g1499 ( 
.A(n_1237),
.B(n_993),
.C(n_1065),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1241),
.A2(n_981),
.B1(n_982),
.B2(n_1065),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1257),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1365),
.A2(n_993),
.B1(n_1118),
.B2(n_1074),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1298),
.A2(n_964),
.B1(n_1204),
.B2(n_993),
.Y(n_1503)
);

OAI221xp5_ASAP7_75t_L g1504 ( 
.A1(n_1237),
.A2(n_993),
.B1(n_1118),
.B2(n_620),
.C(n_964),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_R g1505 ( 
.A(n_1308),
.B(n_757),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1256),
.A2(n_964),
.B1(n_636),
.B2(n_596),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1348),
.B(n_1254),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1257),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1348),
.B(n_1254),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1377),
.B(n_740),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1257),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1298),
.A2(n_964),
.B1(n_1204),
.B2(n_993),
.Y(n_1512)
);

INVx8_ASAP7_75t_L g1513 ( 
.A(n_1264),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1256),
.A2(n_964),
.B1(n_636),
.B2(n_596),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1256),
.B(n_392),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1257),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1344),
.A2(n_1340),
.B(n_1242),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1262),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1269),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1308),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1241),
.A2(n_981),
.B1(n_982),
.B2(n_1065),
.Y(n_1521)
);

AOI21xp33_ASAP7_75t_L g1522 ( 
.A1(n_1376),
.A2(n_1065),
.B(n_993),
.Y(n_1522)
);

AND2x6_ASAP7_75t_L g1523 ( 
.A(n_1372),
.B(n_1233),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1256),
.A2(n_964),
.B1(n_636),
.B2(n_596),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1348),
.B(n_1254),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1328),
.A2(n_1316),
.B(n_1268),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1328),
.A2(n_1316),
.B(n_1268),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1409),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1504),
.A2(n_1492),
.B1(n_1500),
.B2(n_1521),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1391),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_SL g1531 ( 
.A1(n_1399),
.A2(n_1411),
.B1(n_1445),
.B2(n_1515),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1395),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1518),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1494),
.A2(n_1503),
.B1(n_1512),
.B2(n_1499),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1428),
.A2(n_1526),
.B(n_1466),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1397),
.A2(n_1497),
.B1(n_1502),
.B2(n_1495),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1397),
.A2(n_1497),
.B1(n_1502),
.B2(n_1495),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1430),
.B(n_1410),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1527),
.A2(n_1491),
.B(n_1480),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_L g1540 ( 
.A(n_1493),
.B(n_1510),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1392),
.B(n_1394),
.Y(n_1541)
);

BUFx4f_ASAP7_75t_SL g1542 ( 
.A(n_1425),
.Y(n_1542)
);

AO221x2_ASAP7_75t_L g1543 ( 
.A1(n_1396),
.A2(n_1436),
.B1(n_1429),
.B2(n_1427),
.C(n_1457),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1522),
.A2(n_1396),
.B1(n_1421),
.B2(n_1488),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1400),
.A2(n_1506),
.B1(n_1524),
.B2(n_1514),
.Y(n_1545)
);

NAND3xp33_ASAP7_75t_L g1546 ( 
.A(n_1489),
.B(n_1421),
.C(n_1415),
.Y(n_1546)
);

AOI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1401),
.A2(n_1427),
.B1(n_1431),
.B2(n_1433),
.C(n_1408),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1390),
.A2(n_1405),
.B1(n_1389),
.B2(n_1413),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1402),
.B(n_1496),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1412),
.B(n_1432),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1448),
.A2(n_1426),
.B1(n_1409),
.B2(n_1417),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1406),
.A2(n_1498),
.B(n_1517),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1419),
.B(n_1435),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1426),
.A2(n_1413),
.B1(n_1418),
.B2(n_1417),
.Y(n_1554)
);

AOI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1456),
.A2(n_1437),
.B1(n_1414),
.B2(n_1424),
.C(n_1508),
.Y(n_1555)
);

AOI221xp5_ASAP7_75t_L g1556 ( 
.A1(n_1456),
.A2(n_1437),
.B1(n_1511),
.B2(n_1516),
.C(n_1501),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1418),
.A2(n_1448),
.B1(n_1507),
.B2(n_1509),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1422),
.Y(n_1558)
);

OAI211xp5_ASAP7_75t_L g1559 ( 
.A1(n_1443),
.A2(n_1420),
.B(n_1447),
.C(n_1442),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1422),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1451),
.A2(n_1525),
.B1(n_1509),
.B2(n_1507),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1393),
.A2(n_1443),
.B1(n_1454),
.B2(n_1498),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1403),
.A2(n_1519),
.B(n_1472),
.C(n_1449),
.Y(n_1563)
);

AOI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1460),
.A2(n_1490),
.B1(n_1487),
.B2(n_1481),
.C(n_1464),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1406),
.A2(n_1517),
.B1(n_1438),
.B2(n_1446),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1461),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1452),
.A2(n_1520),
.B1(n_1462),
.B2(n_1468),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_SL g1568 ( 
.A1(n_1478),
.A2(n_1477),
.B(n_1460),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1423),
.B(n_1453),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1458),
.B(n_1471),
.Y(n_1570)
);

OAI221xp5_ASAP7_75t_L g1571 ( 
.A1(n_1505),
.A2(n_1478),
.B1(n_1455),
.B2(n_1476),
.C(n_1474),
.Y(n_1571)
);

AND2x2_ASAP7_75t_SL g1572 ( 
.A(n_1473),
.B(n_1475),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1470),
.A2(n_1467),
.B1(n_1469),
.B2(n_1463),
.C(n_1459),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1523),
.A2(n_1513),
.B1(n_1471),
.B2(n_1404),
.Y(n_1574)
);

OAI211xp5_ASAP7_75t_L g1575 ( 
.A1(n_1470),
.A2(n_1444),
.B(n_1441),
.C(n_1479),
.Y(n_1575)
);

AOI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1469),
.A2(n_1486),
.B1(n_1482),
.B2(n_1434),
.C(n_1479),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1471),
.Y(n_1577)
);

OAI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1404),
.A2(n_1416),
.B1(n_1513),
.B2(n_1407),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1473),
.A2(n_1404),
.B1(n_1416),
.B2(n_1513),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1450),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1440),
.B(n_1450),
.Y(n_1581)
);

INVx3_ASAP7_75t_SL g1582 ( 
.A(n_1523),
.Y(n_1582)
);

AOI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1484),
.A2(n_1485),
.B1(n_1440),
.B2(n_1450),
.C(n_1483),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1523),
.A2(n_1440),
.B1(n_1450),
.B2(n_1483),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1440),
.Y(n_1585)
);

AOI222xp33_ASAP7_75t_L g1586 ( 
.A1(n_1483),
.A2(n_1504),
.B1(n_1492),
.B2(n_964),
.C1(n_1118),
.C2(n_1503),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1503),
.B2(n_1494),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1503),
.B2(n_1494),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1439),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1503),
.B2(n_1494),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1419),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1492),
.B2(n_1494),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1492),
.B2(n_1494),
.Y(n_1593)
);

OAI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1504),
.A2(n_993),
.B1(n_1207),
.B2(n_1445),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1419),
.Y(n_1595)
);

OAI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1494),
.A2(n_1512),
.B(n_1503),
.C(n_1504),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1492),
.B2(n_1494),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1503),
.B2(n_1494),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1398),
.Y(n_1599)
);

INVx5_ASAP7_75t_SL g1600 ( 
.A(n_1404),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1504),
.A2(n_993),
.B1(n_1207),
.B2(n_1492),
.Y(n_1601)
);

AND2x6_ASAP7_75t_L g1602 ( 
.A(n_1474),
.B(n_1404),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1392),
.B(n_1394),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1391),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1391),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1391),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1503),
.B2(n_1494),
.Y(n_1607)
);

OAI211xp5_ASAP7_75t_L g1608 ( 
.A1(n_1494),
.A2(n_1512),
.B(n_1503),
.C(n_1504),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1493),
.B(n_1510),
.Y(n_1609)
);

AOI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1504),
.A2(n_1512),
.B1(n_1503),
.B2(n_1494),
.C(n_1497),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1503),
.B2(n_1494),
.Y(n_1611)
);

AO221x1_ASAP7_75t_L g1612 ( 
.A1(n_1396),
.A2(n_1497),
.B1(n_1288),
.B2(n_1464),
.C(n_1411),
.Y(n_1612)
);

OAI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1504),
.A2(n_993),
.B1(n_1207),
.B2(n_1492),
.Y(n_1613)
);

AOI222xp33_ASAP7_75t_L g1614 ( 
.A1(n_1504),
.A2(n_1492),
.B1(n_964),
.B2(n_1118),
.C1(n_1503),
.C2(n_1494),
.Y(n_1614)
);

OAI211xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1504),
.A2(n_1237),
.B(n_1270),
.C(n_1492),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1494),
.A2(n_1512),
.B1(n_1503),
.B2(n_1504),
.Y(n_1616)
);

CKINVDCx8_ASAP7_75t_R g1617 ( 
.A(n_1393),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1494),
.A2(n_1512),
.B1(n_1503),
.B2(n_1504),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1503),
.B2(n_1494),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1492),
.B2(n_993),
.Y(n_1620)
);

INVx5_ASAP7_75t_L g1621 ( 
.A(n_1513),
.Y(n_1621)
);

AO31x2_ASAP7_75t_L g1622 ( 
.A1(n_1487),
.A2(n_1481),
.A3(n_1133),
.B(n_1465),
.Y(n_1622)
);

AOI222xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1398),
.A2(n_534),
.B1(n_588),
.B2(n_267),
.C1(n_226),
.C2(n_323),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1402),
.B(n_1394),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1503),
.B2(n_1494),
.Y(n_1625)
);

AO31x2_ASAP7_75t_L g1626 ( 
.A1(n_1487),
.A2(n_1481),
.A3(n_1133),
.B(n_1465),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1494),
.A2(n_1512),
.B1(n_1503),
.B2(n_1504),
.Y(n_1627)
);

AOI221xp5_ASAP7_75t_L g1628 ( 
.A1(n_1504),
.A2(n_1512),
.B1(n_1503),
.B2(n_1494),
.C(n_1497),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1504),
.A2(n_964),
.B1(n_1503),
.B2(n_1494),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1504),
.A2(n_1512),
.B1(n_1503),
.B2(n_1494),
.C(n_1497),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1504),
.A2(n_1065),
.B(n_964),
.Y(n_1631)
);

INVx4_ASAP7_75t_L g1632 ( 
.A(n_1513),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1392),
.B(n_1394),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1494),
.A2(n_1512),
.B1(n_1503),
.B2(n_1504),
.Y(n_1634)
);

OA21x2_ASAP7_75t_L g1635 ( 
.A1(n_1552),
.A2(n_1583),
.B(n_1584),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1584),
.B(n_1580),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1581),
.B(n_1585),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1535),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1539),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1530),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1622),
.B(n_1626),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1622),
.B(n_1626),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1622),
.B(n_1626),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1565),
.B(n_1569),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_SL g1645 ( 
.A1(n_1616),
.A2(n_1634),
.B1(n_1618),
.B2(n_1627),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1602),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1558),
.B(n_1560),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1565),
.B(n_1549),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1532),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1568),
.B(n_1624),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1564),
.B(n_1572),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1543),
.B(n_1559),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1572),
.B(n_1573),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1543),
.B(n_1554),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1543),
.B(n_1604),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1605),
.B(n_1606),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1556),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_SL g1658 ( 
.A(n_1614),
.B(n_1620),
.C(n_1531),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1562),
.B(n_1547),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1589),
.Y(n_1660)
);

NOR2x1_ASAP7_75t_R g1661 ( 
.A(n_1621),
.B(n_1632),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1536),
.B(n_1537),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1536),
.B(n_1537),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_SL g1664 ( 
.A(n_1546),
.B(n_1579),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1540),
.B(n_1541),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1582),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1555),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1563),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1575),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1603),
.B(n_1633),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1602),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1612),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1576),
.B(n_1586),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1599),
.Y(n_1674)
);

OAI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1587),
.A2(n_1619),
.B1(n_1625),
.B2(n_1611),
.C(n_1590),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1544),
.B(n_1548),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1551),
.B(n_1544),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1548),
.B(n_1631),
.Y(n_1678)
);

OAI31xp33_ASAP7_75t_SL g1679 ( 
.A1(n_1596),
.A2(n_1608),
.A3(n_1613),
.B(n_1601),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1609),
.B(n_1529),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1529),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1534),
.B(n_1628),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1658),
.A2(n_1610),
.B1(n_1630),
.B2(n_1587),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1665),
.B(n_1534),
.Y(n_1684)
);

AOI33xp33_ASAP7_75t_L g1685 ( 
.A1(n_1645),
.A2(n_1590),
.A3(n_1629),
.B1(n_1625),
.B2(n_1598),
.B3(n_1607),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1649),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1644),
.B(n_1550),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1658),
.A2(n_1588),
.B1(n_1598),
.B2(n_1629),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1640),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1673),
.A2(n_1615),
.B1(n_1588),
.B2(n_1611),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1640),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_R g1692 ( 
.A(n_1666),
.B(n_1617),
.Y(n_1692)
);

OAI211xp5_ASAP7_75t_L g1693 ( 
.A1(n_1645),
.A2(n_1607),
.B(n_1619),
.C(n_1593),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1675),
.A2(n_1592),
.B1(n_1597),
.B2(n_1601),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1667),
.A2(n_1613),
.B1(n_1545),
.B2(n_1594),
.C(n_1571),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1644),
.B(n_1538),
.Y(n_1696)
);

AO21x2_ASAP7_75t_L g1697 ( 
.A1(n_1639),
.A2(n_1545),
.B(n_1578),
.Y(n_1697)
);

AOI221x1_ASAP7_75t_SL g1698 ( 
.A1(n_1682),
.A2(n_1623),
.B1(n_1578),
.B2(n_1570),
.C(n_1542),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1673),
.A2(n_1557),
.B1(n_1561),
.B2(n_1591),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1657),
.A2(n_1577),
.B1(n_1528),
.B2(n_1567),
.C(n_1595),
.Y(n_1700)
);

NAND4xp25_ASAP7_75t_L g1701 ( 
.A(n_1679),
.B(n_1566),
.C(n_1574),
.D(n_1553),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1656),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1640),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1673),
.A2(n_1595),
.B1(n_1542),
.B2(n_1533),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1675),
.A2(n_1600),
.B1(n_1676),
.B2(n_1678),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1644),
.B(n_1636),
.Y(n_1706)
);

AND2x6_ASAP7_75t_L g1707 ( 
.A(n_1646),
.B(n_1666),
.Y(n_1707)
);

INVxp67_ASAP7_75t_SL g1708 ( 
.A(n_1660),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1682),
.A2(n_1652),
.B1(n_1677),
.B2(n_1662),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1678),
.A2(n_1654),
.B1(n_1659),
.B2(n_1676),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1666),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1652),
.A2(n_1677),
.B1(n_1662),
.B2(n_1663),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1644),
.B(n_1636),
.Y(n_1713)
);

NAND4xp25_ASAP7_75t_L g1714 ( 
.A(n_1680),
.B(n_1677),
.C(n_1678),
.D(n_1669),
.Y(n_1714)
);

INVx5_ASAP7_75t_L g1715 ( 
.A(n_1666),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1648),
.B(n_1647),
.Y(n_1716)
);

NAND2xp33_ASAP7_75t_SL g1717 ( 
.A(n_1662),
.B(n_1663),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1670),
.B(n_1680),
.Y(n_1718)
);

NAND4xp75_ASAP7_75t_L g1719 ( 
.A(n_1678),
.B(n_1654),
.C(n_1659),
.D(n_1676),
.Y(n_1719)
);

OAI33xp33_ASAP7_75t_L g1720 ( 
.A1(n_1650),
.A2(n_1669),
.A3(n_1668),
.B1(n_1681),
.B2(n_1637),
.B3(n_1647),
.Y(n_1720)
);

NOR2x2_ASAP7_75t_L g1721 ( 
.A(n_1672),
.B(n_1671),
.Y(n_1721)
);

OAI211xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1657),
.A2(n_1669),
.B(n_1668),
.C(n_1681),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1644),
.B(n_1636),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1723),
.B(n_1635),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1686),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1706),
.B(n_1635),
.Y(n_1726)
);

NOR3xp33_ASAP7_75t_L g1727 ( 
.A(n_1693),
.B(n_1695),
.C(n_1694),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1706),
.B(n_1635),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1718),
.B(n_1656),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1721),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1709),
.B(n_1650),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1713),
.B(n_1635),
.Y(n_1732)
);

AND2x4_ASAP7_75t_SL g1733 ( 
.A(n_1711),
.B(n_1666),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1688),
.A2(n_1683),
.B1(n_1690),
.B2(n_1663),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1713),
.B(n_1723),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1707),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1702),
.B(n_1643),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1702),
.B(n_1643),
.Y(n_1738)
);

NOR2xp67_ASAP7_75t_L g1739 ( 
.A(n_1715),
.B(n_1638),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1716),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1689),
.Y(n_1741)
);

INVx6_ASAP7_75t_L g1742 ( 
.A(n_1715),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1708),
.B(n_1641),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1721),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1707),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1691),
.Y(n_1746)
);

BUFx2_ASAP7_75t_L g1747 ( 
.A(n_1707),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1703),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1696),
.B(n_1643),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1746),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1746),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1725),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1727),
.B(n_1685),
.C(n_1722),
.Y(n_1753)
);

OR2x6_ASAP7_75t_L g1754 ( 
.A(n_1742),
.B(n_1666),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1724),
.B(n_1697),
.Y(n_1755)
);

INVx5_ASAP7_75t_L g1756 ( 
.A(n_1742),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1731),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1724),
.B(n_1697),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1725),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1741),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1724),
.B(n_1697),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1741),
.Y(n_1762)
);

INVxp67_ASAP7_75t_SL g1763 ( 
.A(n_1725),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1741),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1748),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1730),
.B(n_1655),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1726),
.B(n_1687),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1748),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1748),
.Y(n_1769)
);

AOI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1727),
.A2(n_1698),
.B1(n_1712),
.B2(n_1710),
.C(n_1720),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1730),
.B(n_1655),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1731),
.B(n_1717),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1726),
.B(n_1642),
.Y(n_1773)
);

INVx2_ASAP7_75t_SL g1774 ( 
.A(n_1742),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1728),
.B(n_1732),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1740),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1744),
.B(n_1648),
.Y(n_1777)
);

OR2x6_ASAP7_75t_L g1778 ( 
.A(n_1742),
.B(n_1666),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1729),
.B(n_1674),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1760),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1753),
.A2(n_1734),
.B1(n_1714),
.B2(n_1705),
.C(n_1717),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1773),
.B(n_1744),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1757),
.B(n_1740),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1776),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1760),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1753),
.A2(n_1770),
.B(n_1664),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1756),
.B(n_1745),
.Y(n_1787)
);

INVxp67_ASAP7_75t_L g1788 ( 
.A(n_1772),
.Y(n_1788)
);

CKINVDCx16_ASAP7_75t_R g1789 ( 
.A(n_1754),
.Y(n_1789)
);

OR2x6_ASAP7_75t_L g1790 ( 
.A(n_1754),
.B(n_1742),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1777),
.B(n_1743),
.Y(n_1791)
);

NOR2x1_ASAP7_75t_L g1792 ( 
.A(n_1754),
.B(n_1719),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1776),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1752),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1762),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1752),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1762),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1764),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1752),
.Y(n_1799)
);

BUFx12f_ASAP7_75t_L g1800 ( 
.A(n_1756),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1770),
.A2(n_1734),
.B1(n_1654),
.B2(n_1662),
.C(n_1663),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1759),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1764),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1759),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1757),
.B(n_1749),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1775),
.B(n_1737),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1765),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1765),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1775),
.B(n_1737),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1768),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1759),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1775),
.B(n_1738),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1768),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1777),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1767),
.B(n_1738),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1750),
.B(n_1749),
.Y(n_1816)
);

NAND2x1_ASAP7_75t_L g1817 ( 
.A(n_1754),
.B(n_1742),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1756),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1756),
.B(n_1745),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1784),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1784),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1792),
.B(n_1756),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1814),
.B(n_1766),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1801),
.A2(n_1654),
.B1(n_1651),
.B2(n_1653),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_L g1825 ( 
.A1(n_1792),
.A2(n_1774),
.B(n_1754),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1793),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1806),
.Y(n_1827)
);

AND2x2_ASAP7_75t_SL g1828 ( 
.A(n_1801),
.B(n_1685),
.Y(n_1828)
);

OAI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1781),
.A2(n_1766),
.B1(n_1771),
.B2(n_1756),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_SL g1830 ( 
.A1(n_1781),
.A2(n_1664),
.B1(n_1676),
.B2(n_1659),
.Y(n_1830)
);

INVxp33_ASAP7_75t_L g1831 ( 
.A(n_1817),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1814),
.B(n_1771),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1789),
.B(n_1756),
.Y(n_1833)
);

NOR2xp67_ASAP7_75t_L g1834 ( 
.A(n_1800),
.B(n_1774),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1789),
.B(n_1774),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1786),
.B(n_1779),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1783),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1793),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1786),
.B(n_1735),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1803),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1800),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1788),
.B(n_1735),
.Y(n_1842)
);

AOI221x1_ASAP7_75t_L g1843 ( 
.A1(n_1783),
.A2(n_1750),
.B1(n_1751),
.B2(n_1769),
.C(n_1745),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1788),
.B(n_1735),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1805),
.B(n_1735),
.Y(n_1845)
);

O2A1O1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1818),
.A2(n_1672),
.B(n_1684),
.C(n_1778),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1800),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1803),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1805),
.B(n_1782),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1807),
.Y(n_1850)
);

OAI31xp33_ASAP7_75t_L g1851 ( 
.A1(n_1818),
.A2(n_1747),
.A3(n_1651),
.B(n_1653),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1817),
.A2(n_1664),
.B(n_1754),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1807),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1782),
.B(n_1767),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1780),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1818),
.B(n_1729),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1835),
.B(n_1782),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1855),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1830),
.A2(n_1651),
.B1(n_1681),
.B2(n_1653),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1836),
.B(n_1791),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1836),
.B(n_1828),
.Y(n_1861)
);

O2A1O1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_1822),
.A2(n_1668),
.B(n_1672),
.C(n_1650),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1849),
.B(n_1791),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1820),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1828),
.A2(n_1817),
.B(n_1790),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1829),
.A2(n_1761),
.B1(n_1758),
.B2(n_1755),
.C(n_1787),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1833),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1835),
.B(n_1787),
.Y(n_1868)
);

OAI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1824),
.A2(n_1672),
.B1(n_1715),
.B2(n_1778),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1837),
.B(n_1791),
.Y(n_1870)
);

NAND4xp25_ASAP7_75t_L g1871 ( 
.A(n_1851),
.B(n_1700),
.C(n_1704),
.D(n_1819),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1847),
.B(n_1787),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1821),
.B(n_1767),
.Y(n_1873)
);

INVx2_ASAP7_75t_SL g1874 ( 
.A(n_1833),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1822),
.A2(n_1790),
.B1(n_1651),
.B2(n_1778),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1826),
.Y(n_1876)
);

A2O1A1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1825),
.A2(n_1755),
.B(n_1761),
.C(n_1758),
.Y(n_1877)
);

OAI21xp33_ASAP7_75t_SL g1878 ( 
.A1(n_1834),
.A2(n_1790),
.B(n_1815),
.Y(n_1878)
);

AOI211xp5_ASAP7_75t_L g1879 ( 
.A1(n_1841),
.A2(n_1819),
.B(n_1787),
.C(n_1653),
.Y(n_1879)
);

OAI21xp33_ASAP7_75t_L g1880 ( 
.A1(n_1839),
.A2(n_1790),
.B(n_1816),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1842),
.B(n_1816),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1838),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1844),
.B(n_1787),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1860),
.B(n_1870),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1857),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1858),
.Y(n_1886)
);

NOR2x1_ASAP7_75t_L g1887 ( 
.A(n_1861),
.B(n_1840),
.Y(n_1887)
);

NAND2x1_ASAP7_75t_SL g1888 ( 
.A(n_1875),
.B(n_1819),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1864),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1876),
.Y(n_1890)
);

NAND2xp33_ASAP7_75t_R g1891 ( 
.A(n_1872),
.B(n_1692),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1882),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1874),
.B(n_1831),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1867),
.B(n_1831),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1873),
.Y(n_1895)
);

INVxp67_ASAP7_75t_SL g1896 ( 
.A(n_1862),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1859),
.A2(n_1843),
.B(n_1852),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1859),
.B(n_1856),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1863),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1868),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1872),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1881),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1883),
.Y(n_1903)
);

NAND4xp25_ASAP7_75t_L g1904 ( 
.A(n_1887),
.B(n_1865),
.C(n_1866),
.D(n_1879),
.Y(n_1904)
);

NAND4xp25_ASAP7_75t_SL g1905 ( 
.A(n_1897),
.B(n_1862),
.C(n_1878),
.D(n_1877),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1901),
.B(n_1871),
.Y(n_1906)
);

OAI221xp5_ASAP7_75t_SL g1907 ( 
.A1(n_1897),
.A2(n_1880),
.B1(n_1869),
.B2(n_1846),
.C(n_1832),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1885),
.B(n_1884),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1900),
.B(n_1856),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1894),
.B(n_1854),
.Y(n_1910)
);

NOR3xp33_ASAP7_75t_L g1911 ( 
.A(n_1893),
.B(n_1869),
.C(n_1850),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1898),
.B(n_1823),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1894),
.B(n_1823),
.Y(n_1913)
);

BUFx2_ASAP7_75t_L g1914 ( 
.A(n_1888),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1899),
.Y(n_1915)
);

NAND3xp33_ASAP7_75t_SL g1916 ( 
.A(n_1903),
.B(n_1832),
.C(n_1848),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1905),
.A2(n_1896),
.B1(n_1891),
.B2(n_1902),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1904),
.A2(n_1896),
.B1(n_1895),
.B2(n_1819),
.Y(n_1918)
);

OAI21xp33_ASAP7_75t_SL g1919 ( 
.A1(n_1912),
.A2(n_1890),
.B(n_1889),
.Y(n_1919)
);

OAI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1907),
.A2(n_1892),
.B1(n_1886),
.B2(n_1790),
.C(n_1853),
.Y(n_1920)
);

AOI211xp5_ASAP7_75t_L g1921 ( 
.A1(n_1916),
.A2(n_1906),
.B(n_1914),
.C(n_1913),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1908),
.Y(n_1922)
);

OAI211xp5_ASAP7_75t_SL g1923 ( 
.A1(n_1910),
.A2(n_1827),
.B(n_1845),
.C(n_1796),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1911),
.A2(n_1819),
.B1(n_1790),
.B2(n_1742),
.Y(n_1924)
);

AOI211xp5_ASAP7_75t_L g1925 ( 
.A1(n_1915),
.A2(n_1827),
.B(n_1747),
.C(n_1701),
.Y(n_1925)
);

AOI221xp5_ASAP7_75t_L g1926 ( 
.A1(n_1909),
.A2(n_1755),
.B1(n_1761),
.B2(n_1758),
.C(n_1785),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1922),
.Y(n_1927)
);

INVxp67_ASAP7_75t_L g1928 ( 
.A(n_1920),
.Y(n_1928)
);

AOI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1921),
.A2(n_1790),
.B1(n_1778),
.B2(n_1747),
.Y(n_1929)
);

A2O1A1Ixp33_ASAP7_75t_L g1930 ( 
.A1(n_1917),
.A2(n_1745),
.B(n_1736),
.C(n_1780),
.Y(n_1930)
);

O2A1O1Ixp5_ASAP7_75t_L g1931 ( 
.A1(n_1919),
.A2(n_1796),
.B(n_1794),
.C(n_1799),
.Y(n_1931)
);

OAI211xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1918),
.A2(n_1796),
.B(n_1802),
.C(n_1794),
.Y(n_1932)
);

OAI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1930),
.A2(n_1924),
.B(n_1925),
.Y(n_1933)
);

NOR2x1_ASAP7_75t_L g1934 ( 
.A(n_1927),
.B(n_1923),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1928),
.B(n_1926),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1929),
.B(n_1815),
.Y(n_1936)
);

NOR2x1p5_ASAP7_75t_L g1937 ( 
.A(n_1932),
.B(n_1745),
.Y(n_1937)
);

AND2x2_ASAP7_75t_SL g1938 ( 
.A(n_1931),
.B(n_1733),
.Y(n_1938)
);

XNOR2x1_ASAP7_75t_L g1939 ( 
.A(n_1927),
.B(n_1778),
.Y(n_1939)
);

NAND4xp25_ASAP7_75t_L g1940 ( 
.A(n_1935),
.B(n_1736),
.C(n_1745),
.D(n_1699),
.Y(n_1940)
);

OAI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1936),
.A2(n_1778),
.B1(n_1813),
.B2(n_1797),
.Y(n_1941)
);

NOR3xp33_ASAP7_75t_SL g1942 ( 
.A(n_1933),
.B(n_1795),
.C(n_1785),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1934),
.Y(n_1943)
);

NOR4xp25_ASAP7_75t_L g1944 ( 
.A(n_1939),
.B(n_1799),
.C(n_1794),
.D(n_1802),
.Y(n_1944)
);

OAI22x1_ASAP7_75t_L g1945 ( 
.A1(n_1937),
.A2(n_1795),
.B1(n_1813),
.B2(n_1798),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1943),
.B(n_1815),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1944),
.B(n_1938),
.Y(n_1947)
);

NOR4xp75_ASAP7_75t_L g1948 ( 
.A(n_1942),
.B(n_1812),
.C(n_1806),
.D(n_1809),
.Y(n_1948)
);

AOI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1940),
.A2(n_1804),
.B1(n_1811),
.B2(n_1799),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1946),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1950),
.Y(n_1951)
);

OAI22x1_ASAP7_75t_L g1952 ( 
.A1(n_1951),
.A2(n_1947),
.B1(n_1948),
.B2(n_1941),
.Y(n_1952)
);

CKINVDCx14_ASAP7_75t_R g1953 ( 
.A(n_1951),
.Y(n_1953)
);

AOI21x1_ASAP7_75t_L g1954 ( 
.A1(n_1952),
.A2(n_1945),
.B(n_1804),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1953),
.A2(n_1949),
.B1(n_1798),
.B2(n_1810),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1954),
.A2(n_1811),
.B1(n_1802),
.B2(n_1804),
.Y(n_1956)
);

AOI222xp33_ASAP7_75t_L g1957 ( 
.A1(n_1955),
.A2(n_1811),
.B1(n_1808),
.B2(n_1810),
.C1(n_1797),
.C2(n_1751),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1956),
.A2(n_1808),
.B1(n_1812),
.B2(n_1806),
.Y(n_1958)
);

OAI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1958),
.A2(n_1957),
.B1(n_1674),
.B2(n_1763),
.C(n_1736),
.Y(n_1959)
);

AOI211xp5_ASAP7_75t_L g1960 ( 
.A1(n_1959),
.A2(n_1661),
.B(n_1739),
.C(n_1692),
.Y(n_1960)
);


endmodule