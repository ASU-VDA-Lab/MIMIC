module fake_aes_10773_n_40 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
wire n_39;
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_6), .A2(n_5), .B1(n_3), .B2(n_8), .Y(n_12) );
CKINVDCx6p67_ASAP7_75t_R g13 ( .A(n_10), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_1), .B(n_11), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_17), .B(n_0), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_15), .A2(n_9), .B(n_2), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_14), .B(n_8), .Y(n_20) );
NAND2xp33_ASAP7_75t_L g21 ( .A(n_17), .B(n_1), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
OAI21x1_ASAP7_75t_L g23 ( .A1(n_18), .A2(n_15), .B(n_17), .Y(n_23) );
O2A1O1Ixp33_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_12), .B(n_16), .C(n_13), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_20), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_22), .A2(n_16), .B1(n_13), .B2(n_12), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_23), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_26), .B(n_24), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
AOI211x1_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_22), .B(n_27), .C(n_24), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_29), .B(n_23), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_29), .Y(n_33) );
OR2x2_ASAP7_75t_L g34 ( .A(n_33), .B(n_32), .Y(n_34) );
OAI21xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_2), .B(n_4), .Y(n_35) );
NAND3xp33_ASAP7_75t_L g36 ( .A(n_31), .B(n_4), .C(n_5), .Y(n_36) );
XNOR2xp5_ASAP7_75t_L g37 ( .A(n_36), .B(n_6), .Y(n_37) );
XNOR2x1_ASAP7_75t_L g38 ( .A(n_35), .B(n_7), .Y(n_38) );
AOI21xp33_ASAP7_75t_SL g39 ( .A1(n_38), .A2(n_34), .B(n_37), .Y(n_39) );
XNOR2xp5_ASAP7_75t_L g40 ( .A(n_39), .B(n_38), .Y(n_40) );
endmodule