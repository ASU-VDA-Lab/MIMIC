module real_aes_7361_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g269 ( .A1(n_0), .A2(n_270), .B(n_271), .C(n_274), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_1), .B(n_211), .Y(n_275) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_2), .B(n_91), .C(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g450 ( .A(n_2), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_3), .B(n_181), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_4), .A2(n_151), .B(n_154), .C(n_480), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_5), .A2(n_171), .B(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_6), .A2(n_171), .B(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_7), .B(n_211), .Y(n_526) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_8), .A2(n_138), .B(n_191), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_9), .A2(n_743), .B1(n_746), .B2(n_747), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_9), .Y(n_747) );
AND2x6_ASAP7_75t_L g151 ( .A(n_10), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_11), .A2(n_151), .B(n_154), .C(n_157), .Y(n_153) );
INVx1_ASAP7_75t_L g496 ( .A(n_12), .Y(n_496) );
INVx1_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_13), .B(n_41), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_14), .A2(n_45), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_14), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_15), .B(n_161), .Y(n_482) );
INVx1_ASAP7_75t_L g143 ( .A(n_16), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_17), .B(n_181), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_18), .A2(n_159), .B(n_504), .C(n_506), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_19), .B(n_211), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_20), .B(n_235), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_21), .A2(n_154), .B(n_198), .C(n_231), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_22), .A2(n_163), .B(n_273), .C(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_23), .B(n_161), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_24), .B(n_161), .Y(n_547) );
CKINVDCx16_ASAP7_75t_R g554 ( .A(n_25), .Y(n_554) );
INVx1_ASAP7_75t_L g546 ( .A(n_26), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_27), .A2(n_154), .B(n_194), .C(n_198), .Y(n_193) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_28), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_29), .Y(n_478) );
INVx1_ASAP7_75t_L g537 ( .A(n_30), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_31), .A2(n_171), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g149 ( .A(n_32), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_33), .A2(n_173), .B(n_184), .C(n_219), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_34), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_35), .A2(n_273), .B(n_523), .C(n_525), .Y(n_522) );
INVxp67_ASAP7_75t_L g538 ( .A(n_36), .Y(n_538) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_37), .A2(n_78), .B1(n_453), .B2(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_37), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_38), .B(n_196), .Y(n_195) );
CKINVDCx14_ASAP7_75t_R g521 ( .A(n_39), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_40), .A2(n_154), .B(n_198), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_41), .B(n_111), .Y(n_110) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_42), .A2(n_274), .B(n_494), .C(n_495), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_43), .B(n_229), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_44), .Y(n_166) );
INVx1_ASAP7_75t_L g745 ( .A(n_45), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_46), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_47), .B(n_171), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_48), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_49), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_50), .A2(n_173), .B(n_175), .C(n_184), .Y(n_172) );
INVx1_ASAP7_75t_L g272 ( .A(n_51), .Y(n_272) );
INVx1_ASAP7_75t_L g176 ( .A(n_52), .Y(n_176) );
AOI222xp33_ASAP7_75t_L g463 ( .A1(n_53), .A2(n_464), .B1(n_738), .B2(n_739), .C1(n_748), .C2(n_751), .Y(n_463) );
INVx1_ASAP7_75t_L g511 ( .A(n_54), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_55), .B(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_56), .A2(n_59), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_56), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_57), .Y(n_238) );
CKINVDCx14_ASAP7_75t_R g492 ( .A(n_58), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_59), .Y(n_126) );
INVx1_ASAP7_75t_L g152 ( .A(n_60), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_61), .B(n_171), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_62), .B(n_211), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_63), .A2(n_205), .B(n_207), .C(n_209), .Y(n_204) );
INVx1_ASAP7_75t_L g142 ( .A(n_64), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_65), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g524 ( .A(n_66), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_67), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_68), .B(n_181), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_69), .B(n_211), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_70), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g557 ( .A(n_71), .Y(n_557) );
CKINVDCx16_ASAP7_75t_R g268 ( .A(n_72), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_73), .B(n_178), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_74), .A2(n_154), .B(n_184), .C(n_245), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g203 ( .A(n_75), .Y(n_203) );
INVx1_ASAP7_75t_L g115 ( .A(n_76), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_77), .A2(n_171), .B(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_78), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_79), .A2(n_171), .B(n_501), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_80), .A2(n_229), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g502 ( .A(n_81), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_82), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_83), .B(n_177), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_84), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_85), .A2(n_171), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g505 ( .A(n_86), .Y(n_505) );
INVx2_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
INVx1_ASAP7_75t_L g481 ( .A(n_88), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_89), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_90), .B(n_161), .Y(n_160) );
OR2x2_ASAP7_75t_L g447 ( .A(n_91), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g467 ( .A(n_91), .B(n_449), .Y(n_467) );
INVx2_ASAP7_75t_L g737 ( .A(n_91), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_92), .A2(n_105), .B1(n_116), .B2(n_756), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_93), .A2(n_154), .B(n_184), .C(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_94), .B(n_171), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_95), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_95), .Y(n_740) );
INVx1_ASAP7_75t_L g220 ( .A(n_96), .Y(n_220) );
INVxp67_ASAP7_75t_L g208 ( .A(n_97), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_98), .B(n_138), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_99), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g145 ( .A(n_100), .Y(n_145) );
INVx1_ASAP7_75t_L g246 ( .A(n_101), .Y(n_246) );
INVx2_ASAP7_75t_L g514 ( .A(n_102), .Y(n_514) );
AND2x2_ASAP7_75t_L g187 ( .A(n_103), .B(n_186), .Y(n_187) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_108), .Y(n_757) );
CKINVDCx9p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_462), .Y(n_116) );
BUFx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g755 ( .A(n_120), .Y(n_755) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI321xp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_445), .A3(n_452), .B1(n_455), .B2(n_456), .C(n_459), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_123), .B(n_457), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_128), .B2(n_129), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22x1_ASAP7_75t_SL g464 ( .A1(n_128), .A2(n_465), .B1(n_468), .B2(n_734), .Y(n_464) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_129), .A2(n_469), .B1(n_749), .B2(n_750), .Y(n_748) );
OR3x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_343), .C(n_408), .Y(n_129) );
NAND4xp25_ASAP7_75t_SL g130 ( .A(n_131), .B(n_284), .C(n_310), .D(n_333), .Y(n_130) );
AOI221xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_212), .B1(n_253), .B2(n_260), .C(n_276), .Y(n_131) );
CKINVDCx14_ASAP7_75t_R g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_133), .A2(n_277), .B1(n_301), .B2(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_188), .Y(n_133) );
INVx1_ASAP7_75t_SL g337 ( .A(n_134), .Y(n_337) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_168), .Y(n_134) );
OR2x2_ASAP7_75t_L g258 ( .A(n_135), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g279 ( .A(n_135), .B(n_189), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_135), .B(n_199), .Y(n_292) );
AND2x2_ASAP7_75t_L g309 ( .A(n_135), .B(n_168), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_135), .B(n_256), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_135), .B(n_308), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_135), .B(n_188), .Y(n_430) );
AOI211xp5_ASAP7_75t_SL g441 ( .A1(n_135), .A2(n_347), .B(n_442), .C(n_443), .Y(n_441) );
INVx5_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_136), .B(n_189), .Y(n_313) );
AND2x2_ASAP7_75t_L g316 ( .A(n_136), .B(n_190), .Y(n_316) );
OR2x2_ASAP7_75t_L g361 ( .A(n_136), .B(n_189), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_136), .B(n_199), .Y(n_370) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_144), .B(n_165), .Y(n_136) );
INVx3_ASAP7_75t_L g211 ( .A(n_137), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_137), .B(n_223), .Y(n_222) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_137), .A2(n_243), .B(n_251), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_137), .B(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_137), .B(n_485), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_137), .B(n_549), .Y(n_548) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_137), .A2(n_553), .B(n_559), .Y(n_552) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_138), .A2(n_192), .B(n_193), .Y(n_191) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_138), .Y(n_200) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g186 ( .A(n_140), .B(n_141), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_153), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_146), .A2(n_478), .B(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_146), .A2(n_186), .B(n_543), .C(n_544), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_146), .A2(n_554), .B(n_555), .Y(n_553) );
NAND2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
AND2x4_ASAP7_75t_L g171 ( .A(n_147), .B(n_151), .Y(n_171) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
INVx1_ASAP7_75t_L g164 ( .A(n_149), .Y(n_164) );
INVx1_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx3_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
INVx1_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
INVx4_ASAP7_75t_SL g185 ( .A(n_151), .Y(n_185) );
BUFx3_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
INVx5_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx3_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_155), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B(n_162), .Y(n_157) );
INVx5_ASAP7_75t_L g181 ( .A(n_159), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_159), .B(n_496), .Y(n_495) );
INVx4_ASAP7_75t_L g273 ( .A(n_161), .Y(n_273) );
INVx2_ASAP7_75t_L g494 ( .A(n_161), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_162), .A2(n_195), .B(n_197), .Y(n_194) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx2_ASAP7_75t_L g531 ( .A(n_167), .Y(n_531) );
INVx5_ASAP7_75t_SL g259 ( .A(n_168), .Y(n_259) );
AND2x2_ASAP7_75t_L g278 ( .A(n_168), .B(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_168), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g364 ( .A(n_168), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g396 ( .A(n_168), .B(n_199), .Y(n_396) );
OR2x2_ASAP7_75t_L g402 ( .A(n_168), .B(n_292), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_168), .B(n_352), .Y(n_411) );
OR2x6_ASAP7_75t_L g168 ( .A(n_169), .B(n_187), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B(n_186), .Y(n_169) );
BUFx2_ASAP7_75t_L g229 ( .A(n_171), .Y(n_229) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_174), .A2(n_185), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_SL g267 ( .A1(n_174), .A2(n_185), .B(n_268), .C(n_269), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_SL g491 ( .A1(n_174), .A2(n_185), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g501 ( .A1(n_174), .A2(n_185), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_SL g510 ( .A1(n_174), .A2(n_185), .B(n_511), .C(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_174), .A2(n_185), .B(n_521), .C(n_522), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_174), .A2(n_185), .B(n_534), .C(n_535), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_180), .C(n_182), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_177), .A2(n_182), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp5_ASAP7_75t_L g480 ( .A1(n_177), .A2(n_481), .B(n_482), .C(n_483), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_177), .A2(n_483), .B(n_557), .C(n_558), .Y(n_556) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx4_ASAP7_75t_L g206 ( .A(n_179), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_181), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g270 ( .A(n_181), .Y(n_270) );
OAI22xp33_ASAP7_75t_L g536 ( .A1(n_181), .A2(n_206), .B1(n_537), .B2(n_538), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_181), .A2(n_234), .B(n_546), .C(n_547), .Y(n_545) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g274 ( .A(n_183), .Y(n_274) );
INVx1_ASAP7_75t_L g506 ( .A(n_183), .Y(n_506) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_186), .A2(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g236 ( .A(n_186), .Y(n_236) );
INVx1_ASAP7_75t_L g239 ( .A(n_186), .Y(n_239) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_186), .A2(n_490), .B(n_497), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_199), .Y(n_188) );
AND2x2_ASAP7_75t_L g293 ( .A(n_189), .B(n_259), .Y(n_293) );
INVx1_ASAP7_75t_SL g306 ( .A(n_189), .Y(n_306) );
OR2x2_ASAP7_75t_L g341 ( .A(n_189), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g347 ( .A(n_189), .B(n_199), .Y(n_347) );
AND2x2_ASAP7_75t_L g405 ( .A(n_189), .B(n_256), .Y(n_405) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_190), .B(n_259), .Y(n_332) );
INVx3_ASAP7_75t_L g256 ( .A(n_199), .Y(n_256) );
OR2x2_ASAP7_75t_L g298 ( .A(n_199), .B(n_259), .Y(n_298) );
AND2x2_ASAP7_75t_L g308 ( .A(n_199), .B(n_306), .Y(n_308) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_199), .Y(n_356) );
AND2x2_ASAP7_75t_L g365 ( .A(n_199), .B(n_279), .Y(n_365) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_210), .Y(n_199) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_200), .A2(n_500), .B(n_507), .Y(n_499) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_200), .A2(n_509), .B(n_515), .Y(n_508) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_200), .A2(n_519), .B(n_526), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_205), .A2(n_246), .B(n_247), .C(n_248), .Y(n_245) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_206), .B(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_206), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g234 ( .A(n_209), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_209), .B(n_536), .Y(n_535) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_211), .A2(n_266), .B(n_275), .Y(n_265) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_212), .A2(n_382), .B1(n_384), .B2(n_386), .C(n_389), .Y(n_381) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
AND2x2_ASAP7_75t_L g355 ( .A(n_214), .B(n_336), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_214), .B(n_414), .Y(n_418) );
OR2x2_ASAP7_75t_L g439 ( .A(n_214), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_214), .B(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx5_ASAP7_75t_L g286 ( .A(n_215), .Y(n_286) );
AND2x2_ASAP7_75t_L g363 ( .A(n_215), .B(n_226), .Y(n_363) );
AND2x2_ASAP7_75t_L g424 ( .A(n_215), .B(n_303), .Y(n_424) );
AND2x2_ASAP7_75t_L g437 ( .A(n_215), .B(n_256), .Y(n_437) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_222), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_240), .Y(n_224) );
AND2x4_ASAP7_75t_L g263 ( .A(n_225), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g282 ( .A(n_225), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g289 ( .A(n_225), .Y(n_289) );
AND2x2_ASAP7_75t_L g358 ( .A(n_225), .B(n_336), .Y(n_358) );
AND2x2_ASAP7_75t_L g368 ( .A(n_225), .B(n_286), .Y(n_368) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_225), .Y(n_376) );
AND2x2_ASAP7_75t_L g388 ( .A(n_225), .B(n_265), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_225), .B(n_320), .Y(n_392) );
AND2x2_ASAP7_75t_L g429 ( .A(n_225), .B(n_424), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_225), .B(n_303), .Y(n_440) );
OR2x2_ASAP7_75t_L g442 ( .A(n_225), .B(n_378), .Y(n_442) );
INVx5_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g328 ( .A(n_226), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g338 ( .A(n_226), .B(n_283), .Y(n_338) );
AND2x2_ASAP7_75t_L g350 ( .A(n_226), .B(n_265), .Y(n_350) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_226), .Y(n_380) );
AND2x4_ASAP7_75t_L g414 ( .A(n_226), .B(n_264), .Y(n_414) );
OR2x6_ASAP7_75t_L g226 ( .A(n_227), .B(n_237), .Y(n_226) );
AOI21xp5_ASAP7_75t_SL g227 ( .A1(n_228), .A2(n_230), .B(n_235), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_236), .B(n_454), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_239), .A2(n_477), .B(n_484), .Y(n_476) );
BUFx2_ASAP7_75t_L g262 ( .A(n_240), .Y(n_262) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g303 ( .A(n_241), .Y(n_303) );
AND2x2_ASAP7_75t_L g336 ( .A(n_241), .B(n_265), .Y(n_336) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g283 ( .A(n_242), .B(n_265), .Y(n_283) );
BUFx2_ASAP7_75t_L g329 ( .A(n_242), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_250), .Y(n_243) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g525 ( .A(n_249), .Y(n_525) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_255), .B(n_337), .Y(n_416) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_256), .B(n_279), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_256), .B(n_259), .Y(n_318) );
AND2x2_ASAP7_75t_L g373 ( .A(n_256), .B(n_309), .Y(n_373) );
AOI221xp5_ASAP7_75t_SL g310 ( .A1(n_257), .A2(n_311), .B1(n_319), .B2(n_321), .C(n_325), .Y(n_310) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g305 ( .A(n_258), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g346 ( .A(n_258), .B(n_347), .Y(n_346) );
OAI321xp33_ASAP7_75t_L g353 ( .A1(n_258), .A2(n_312), .A3(n_354), .B1(n_356), .B2(n_357), .C(n_359), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_259), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_262), .B(n_414), .Y(n_432) );
AND2x2_ASAP7_75t_L g319 ( .A(n_263), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_263), .B(n_323), .Y(n_322) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_264), .Y(n_295) );
AND2x2_ASAP7_75t_L g302 ( .A(n_264), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_264), .B(n_377), .Y(n_407) );
INVx1_ASAP7_75t_L g444 ( .A(n_264), .Y(n_444) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_273), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g483 ( .A(n_274), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B(n_281), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_278), .A2(n_388), .B(n_437), .C(n_438), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_279), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_279), .B(n_317), .Y(n_383) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g326 ( .A(n_283), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_283), .B(n_286), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_283), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_283), .B(n_368), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_287), .B1(n_299), .B2(n_304), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g300 ( .A(n_286), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g323 ( .A(n_286), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g335 ( .A(n_286), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_286), .B(n_329), .Y(n_371) );
OR2x2_ASAP7_75t_L g378 ( .A(n_286), .B(n_303), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_286), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g428 ( .A(n_286), .B(n_414), .Y(n_428) );
OAI22xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .B1(n_294), .B2(n_296), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g334 ( .A(n_289), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_292), .A2(n_307), .B1(n_375), .B2(n_379), .Y(n_374) );
INVx1_ASAP7_75t_L g422 ( .A(n_293), .Y(n_422) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_297), .A2(n_334), .B1(n_337), .B2(n_338), .C(n_339), .Y(n_333) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g312 ( .A(n_298), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_302), .B(n_368), .Y(n_400) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_303), .Y(n_320) );
INVx1_ASAP7_75t_L g324 ( .A(n_303), .Y(n_324) );
NAND2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g342 ( .A(n_309), .Y(n_342) );
AND2x2_ASAP7_75t_L g351 ( .A(n_309), .B(n_352), .Y(n_351) );
NAND2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx2_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g395 ( .A(n_316), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_319), .A2(n_345), .B1(n_348), .B2(n_351), .C(n_353), .Y(n_344) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_323), .B(n_380), .Y(n_379) );
AOI21xp33_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_327), .B(n_330), .Y(n_325) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g427 ( .A(n_330), .Y(n_427) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OR2x2_ASAP7_75t_L g369 ( .A(n_332), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g390 ( .A(n_335), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_335), .B(n_395), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_338), .B(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND4xp25_ASAP7_75t_L g343 ( .A(n_344), .B(n_362), .C(n_381), .D(n_394), .Y(n_343) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g352 ( .A(n_347), .Y(n_352) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g385 ( .A(n_356), .B(n_361), .Y(n_385) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI211xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B(n_366), .C(n_374), .Y(n_362) );
AOI211xp5_ASAP7_75t_L g433 ( .A1(n_364), .A2(n_406), .B(n_434), .C(n_441), .Y(n_433) );
INVx1_ASAP7_75t_SL g393 ( .A(n_365), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B1(n_371), .B2(n_372), .Y(n_366) );
INVx1_ASAP7_75t_L g397 ( .A(n_371), .Y(n_397) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_377), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_377), .B(n_388), .Y(n_421) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g398 ( .A(n_388), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B(n_393), .Y(n_389) );
INVxp33_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI322xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .A3(n_398), .B1(n_399), .B2(n_401), .C1(n_403), .C2(n_406), .Y(n_394) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND3xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_426), .C(n_433), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B1(n_415), .B2(n_417), .C(n_419), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g425 ( .A(n_414), .Y(n_425) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_429), .B2(n_430), .C(n_431), .Y(n_426) );
NAND2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVxp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g458 ( .A(n_447), .Y(n_458) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_447), .Y(n_461) );
NOR2x2_ASAP7_75t_L g753 ( .A(n_448), .B(n_737), .Y(n_753) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g736 ( .A(n_449), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g455 ( .A(n_452), .Y(n_455) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_459), .B(n_463), .C(n_754), .Y(n_462) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g749 ( .A(n_466), .Y(n_749) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_SL g469 ( .A(n_470), .B(n_689), .Y(n_469) );
NAND5xp2_ASAP7_75t_L g470 ( .A(n_471), .B(n_601), .C(n_639), .D(n_660), .E(n_677), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_573), .C(n_594), .Y(n_471) );
OAI221xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_516), .B1(n_540), .B2(n_560), .C(n_564), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_486), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_475), .B(n_562), .Y(n_581) );
OR2x2_ASAP7_75t_L g608 ( .A(n_475), .B(n_499), .Y(n_608) );
AND2x2_ASAP7_75t_L g622 ( .A(n_475), .B(n_499), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_475), .B(n_489), .Y(n_636) );
AND2x2_ASAP7_75t_L g674 ( .A(n_475), .B(n_638), .Y(n_674) );
AND2x2_ASAP7_75t_L g703 ( .A(n_475), .B(n_613), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_475), .B(n_585), .Y(n_720) );
INVx4_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g600 ( .A(n_476), .B(n_498), .Y(n_600) );
BUFx3_ASAP7_75t_L g625 ( .A(n_476), .Y(n_625) );
AND2x2_ASAP7_75t_L g654 ( .A(n_476), .B(n_499), .Y(n_654) );
AND3x2_ASAP7_75t_L g667 ( .A(n_476), .B(n_668), .C(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g590 ( .A(n_486), .Y(n_590) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
AOI32xp33_ASAP7_75t_L g645 ( .A1(n_487), .A2(n_597), .A3(n_646), .B1(n_649), .B2(n_650), .Y(n_645) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g572 ( .A(n_488), .B(n_498), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_488), .B(n_600), .Y(n_643) );
AND2x2_ASAP7_75t_L g650 ( .A(n_488), .B(n_622), .Y(n_650) );
OR2x2_ASAP7_75t_L g656 ( .A(n_488), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_488), .B(n_611), .Y(n_681) );
OR2x2_ASAP7_75t_L g699 ( .A(n_488), .B(n_528), .Y(n_699) );
BUFx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g563 ( .A(n_489), .B(n_508), .Y(n_563) );
INVx2_ASAP7_75t_L g585 ( .A(n_489), .Y(n_585) );
OR2x2_ASAP7_75t_L g607 ( .A(n_489), .B(n_508), .Y(n_607) );
AND2x2_ASAP7_75t_L g612 ( .A(n_489), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_489), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g668 ( .A(n_489), .B(n_562), .Y(n_668) );
INVx1_ASAP7_75t_SL g719 ( .A(n_498), .Y(n_719) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
INVx1_ASAP7_75t_SL g562 ( .A(n_499), .Y(n_562) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_499), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_499), .B(n_648), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_499), .B(n_585), .C(n_703), .Y(n_714) );
INVx2_ASAP7_75t_L g613 ( .A(n_508), .Y(n_613) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_508), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
INVx1_ASAP7_75t_L g649 ( .A(n_517), .Y(n_649) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g567 ( .A(n_518), .B(n_551), .Y(n_567) );
INVx2_ASAP7_75t_L g584 ( .A(n_518), .Y(n_584) );
AND2x2_ASAP7_75t_L g589 ( .A(n_518), .B(n_552), .Y(n_589) );
AND2x2_ASAP7_75t_L g604 ( .A(n_518), .B(n_541), .Y(n_604) );
AND2x2_ASAP7_75t_L g616 ( .A(n_518), .B(n_588), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_527), .B(n_632), .Y(n_631) );
NAND2x1p5_ASAP7_75t_L g688 ( .A(n_527), .B(n_589), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_527), .B(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_527), .B(n_583), .Y(n_711) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g550 ( .A(n_528), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_528), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g593 ( .A(n_528), .B(n_541), .Y(n_593) );
AND2x2_ASAP7_75t_L g619 ( .A(n_528), .B(n_551), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_528), .B(n_659), .Y(n_658) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_532), .B(n_539), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_530), .A2(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g578 ( .A(n_532), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_539), .Y(n_579) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_550), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_541), .B(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g583 ( .A(n_541), .B(n_584), .Y(n_583) );
INVx3_ASAP7_75t_SL g588 ( .A(n_541), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_541), .B(n_575), .Y(n_641) );
OR2x2_ASAP7_75t_L g651 ( .A(n_541), .B(n_577), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_541), .B(n_619), .Y(n_679) );
OR2x2_ASAP7_75t_L g709 ( .A(n_541), .B(n_551), .Y(n_709) );
AND2x2_ASAP7_75t_L g713 ( .A(n_541), .B(n_552), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_541), .B(n_589), .Y(n_726) );
AND2x2_ASAP7_75t_L g733 ( .A(n_541), .B(n_615), .Y(n_733) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_548), .Y(n_541) );
INVx1_ASAP7_75t_SL g676 ( .A(n_550), .Y(n_676) );
AND2x2_ASAP7_75t_L g615 ( .A(n_551), .B(n_577), .Y(n_615) );
AND2x2_ASAP7_75t_L g629 ( .A(n_551), .B(n_584), .Y(n_629) );
AND2x2_ASAP7_75t_L g632 ( .A(n_551), .B(n_588), .Y(n_632) );
INVx1_ASAP7_75t_L g659 ( .A(n_551), .Y(n_659) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
BUFx2_ASAP7_75t_L g571 ( .A(n_552), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g730 ( .A1(n_561), .A2(n_607), .B(n_731), .C(n_732), .Y(n_730) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g637 ( .A(n_562), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_563), .B(n_580), .Y(n_595) );
AND2x2_ASAP7_75t_L g621 ( .A(n_563), .B(n_622), .Y(n_621) );
OAI21xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_568), .B(n_572), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_566), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g592 ( .A(n_567), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_567), .B(n_588), .Y(n_633) );
AND2x2_ASAP7_75t_L g724 ( .A(n_567), .B(n_575), .Y(n_724) );
INVxp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g597 ( .A(n_571), .B(n_584), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_571), .B(n_582), .Y(n_598) );
OAI322xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_581), .A3(n_582), .B1(n_585), .B2(n_586), .C1(n_590), .C2(n_591), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_580), .Y(n_574) );
AND2x2_ASAP7_75t_L g685 ( .A(n_575), .B(n_597), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_575), .B(n_649), .Y(n_731) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g628 ( .A(n_577), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g694 ( .A(n_581), .B(n_607), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_582), .B(n_676), .Y(n_675) );
INVx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_583), .B(n_615), .Y(n_672) );
AND2x2_ASAP7_75t_L g618 ( .A(n_584), .B(n_588), .Y(n_618) );
AND2x2_ASAP7_75t_L g626 ( .A(n_585), .B(n_627), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g723 ( .A1(n_585), .A2(n_664), .B(n_724), .C(n_725), .Y(n_723) );
AOI21xp33_ASAP7_75t_L g696 ( .A1(n_586), .A2(n_599), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_588), .B(n_615), .Y(n_655) );
AND2x2_ASAP7_75t_L g661 ( .A(n_588), .B(n_629), .Y(n_661) );
AND2x2_ASAP7_75t_L g695 ( .A(n_588), .B(n_597), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_589), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g705 ( .A(n_589), .Y(n_705) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_593), .A2(n_621), .B1(n_623), .B2(n_628), .Y(n_620) );
OAI22xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_596), .B1(n_598), .B2(n_599), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g630 ( .A1(n_595), .A2(n_631), .B1(n_633), .B2(n_634), .Y(n_630) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_600), .A2(n_702), .B1(n_704), .B2(n_706), .C(n_710), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B(n_609), .C(n_630), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OR2x2_ASAP7_75t_L g671 ( .A(n_607), .B(n_624), .Y(n_671) );
INVx1_ASAP7_75t_L g722 ( .A(n_607), .Y(n_722) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_608), .A2(n_610), .B1(n_614), .B2(n_617), .C(n_620), .Y(n_609) );
INVx2_ASAP7_75t_SL g664 ( .A(n_608), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g729 ( .A(n_611), .Y(n_729) );
AND2x2_ASAP7_75t_L g653 ( .A(n_612), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g638 ( .A(n_613), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g700 ( .A(n_616), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_624), .B(n_726), .Y(n_725) );
CKINVDCx16_ASAP7_75t_R g624 ( .A(n_625), .Y(n_624) );
INVxp67_ASAP7_75t_L g669 ( .A(n_627), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_628), .A2(n_640), .B(n_642), .C(n_644), .Y(n_639) );
INVx1_ASAP7_75t_L g717 ( .A(n_631), .Y(n_717) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_635), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx2_ASAP7_75t_L g648 ( .A(n_638), .Y(n_648) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI222xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_651), .B1(n_652), .B2(n_655), .C1(n_656), .C2(n_658), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g684 ( .A(n_648), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_651), .B(n_705), .Y(n_704) );
NAND2xp33_ASAP7_75t_SL g682 ( .A(n_652), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g657 ( .A(n_654), .Y(n_657) );
AND2x2_ASAP7_75t_L g721 ( .A(n_654), .B(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g687 ( .A(n_657), .B(n_684), .Y(n_687) );
INVx1_ASAP7_75t_L g716 ( .A(n_658), .Y(n_716) );
AOI211xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B(n_665), .C(n_670), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_664), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AOI322xp5_ASAP7_75t_L g715 ( .A1(n_667), .A2(n_695), .A3(n_700), .B1(n_716), .B2(n_717), .C1(n_718), .C2(n_721), .Y(n_715) );
AND2x2_ASAP7_75t_L g702 ( .A(n_668), .B(n_703), .Y(n_702) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B1(n_673), .B2(n_675), .Y(n_670) );
INVxp33_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B1(n_682), .B2(n_685), .C(n_686), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NAND5xp2_ASAP7_75t_L g689 ( .A(n_690), .B(n_701), .C(n_715), .D(n_723), .E(n_727), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_695), .B(n_696), .Y(n_690) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVxp33_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_703), .A2(n_728), .B(n_729), .C(n_730), .Y(n_727) );
AOI31xp33_ASAP7_75t_L g710 ( .A1(n_705), .A2(n_711), .A3(n_712), .B(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVx1_ASAP7_75t_L g728 ( .A(n_726), .Y(n_728) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g750 ( .A(n_735), .Y(n_750) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_743), .Y(n_746) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx3_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
endmodule