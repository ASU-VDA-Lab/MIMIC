module fake_aes_12556_n_1142 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_137, n_277, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_210, n_184, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1142);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_210;
input n_184;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1142;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_1056;
wire n_802;
wire n_985;
wire n_856;
wire n_564;
wire n_353;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_971;
wire n_1128;
wire n_661;
wire n_850;
wire n_762;
wire n_904;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_599;
wire n_724;
wire n_857;
wire n_786;
wire n_360;
wire n_345;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1078;
wire n_1097;
wire n_572;
wire n_1017;
wire n_324;
wire n_1125;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_880;
wire n_1101;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_1018;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_910;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_415;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_990;
wire n_751;
wire n_800;
wire n_626;
wire n_941;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_601;
wire n_439;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_420;
wire n_446;
wire n_423;
wire n_621;
wire n_342;
wire n_666;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_597;
wire n_349;
wire n_723;
wire n_972;
wire n_1069;
wire n_1021;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_947;
wire n_924;
wire n_1043;
wire n_912;
wire n_582;
wire n_378;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_766;
wire n_602;
wire n_1007;
wire n_1027;
wire n_1117;
wire n_859;
wire n_831;
wire n_1040;
wire n_994;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_1016;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_695;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_405;
wire n_819;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_303), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_155), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_80), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_100), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_147), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_68), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_238), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_134), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_285), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_55), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_62), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_160), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_307), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_184), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_282), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_105), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_8), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_102), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_276), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_199), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_76), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_281), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_16), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_300), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_217), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_288), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_133), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_294), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_248), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_15), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_265), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_180), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_198), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_246), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_152), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_251), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_204), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_63), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_269), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_286), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_301), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_226), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_234), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_74), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_137), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_26), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_89), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_77), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_215), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_167), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g361 ( .A(n_73), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_87), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_299), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_119), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_195), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_86), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_90), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_260), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_72), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_197), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_240), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_241), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_212), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_57), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_111), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_5), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_37), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_187), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_4), .Y(n_379) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_235), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_283), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_297), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_209), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_53), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_51), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_185), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_88), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_5), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_278), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_158), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_41), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_161), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_196), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_255), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_18), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_19), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_284), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_65), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_59), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_44), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_75), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_46), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_275), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_42), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_23), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_33), .Y(n_406) );
BUFx10_ASAP7_75t_L g407 ( .A(n_183), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_279), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_7), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_150), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_273), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_290), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_10), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_70), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_54), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_289), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_39), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_302), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_213), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_14), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_218), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_47), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_121), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_205), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_140), .Y(n_425) );
BUFx5_ASAP7_75t_L g426 ( .A(n_280), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_23), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_113), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_210), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_263), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_229), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_12), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_6), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_206), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_308), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_103), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_48), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_262), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_291), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_159), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_201), .Y(n_441) );
CKINVDCx16_ASAP7_75t_R g442 ( .A(n_36), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_274), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_151), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_50), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_128), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_9), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_200), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_177), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_287), .Y(n_450) );
INVxp67_ASAP7_75t_L g451 ( .A(n_32), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_67), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_230), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_309), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_295), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_267), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_250), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_83), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_35), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_306), .Y(n_460) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_97), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_170), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_271), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_143), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_58), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_6), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_14), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_292), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_116), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_293), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_277), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_26), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_146), .Y(n_473) );
OAI21x1_ASAP7_75t_L g474 ( .A1(n_355), .A2(n_38), .B(n_34), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_321), .Y(n_475) );
INVx5_ASAP7_75t_L g476 ( .A(n_407), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_344), .B(n_0), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_357), .B(n_0), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_368), .B(n_1), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_453), .B(n_1), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_409), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_376), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_356), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_388), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_484) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_316), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_426), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_426), .Y(n_487) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_316), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_316), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_366), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_366), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_366), .Y(n_492) );
INVx5_ASAP7_75t_L g493 ( .A(n_407), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_361), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_432), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_455), .B(n_2), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_396), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_442), .B(n_3), .Y(n_498) );
OAI21x1_ASAP7_75t_L g499 ( .A1(n_369), .A2(n_43), .B(n_40), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_346), .Y(n_500) );
AND2x2_ASAP7_75t_SL g501 ( .A(n_311), .B(n_45), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_451), .B(n_7), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_494), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_494), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_498), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_481), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_476), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_481), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_483), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_476), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_482), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_486), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_495), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_476), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_476), .B(n_326), .Y(n_515) );
NOR2x1p5_ASAP7_75t_L g516 ( .A(n_475), .B(n_333), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_479), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_480), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_486), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_487), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_487), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_485), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_485), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_496), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_500), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_519), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_524), .B(n_480), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_518), .B(n_480), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_519), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_519), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_520), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_515), .B(n_493), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_507), .B(n_493), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_508), .B(n_477), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_506), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_514), .B(n_477), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_514), .B(n_501), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_507), .B(n_493), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_525), .B(n_493), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_510), .B(n_500), .Y(n_540) );
AND2x4_ASAP7_75t_SL g541 ( .A(n_509), .B(n_324), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_511), .B(n_478), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_505), .B(n_501), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_503), .B(n_502), .Y(n_544) );
INVx4_ASAP7_75t_L g545 ( .A(n_520), .Y(n_545) );
INVx4_ASAP7_75t_L g546 ( .A(n_520), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_513), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_516), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_512), .B(n_478), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_512), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_521), .B(n_310), .Y(n_551) );
NAND2xp33_ASAP7_75t_L g552 ( .A(n_521), .B(n_426), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_517), .B(n_312), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_504), .B(n_395), .Y(n_554) );
BUFx6f_ASAP7_75t_SL g555 ( .A(n_509), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_517), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_527), .B(n_420), .Y(n_557) );
O2A1O1Ixp5_ASAP7_75t_L g558 ( .A1(n_537), .A2(n_423), .B(n_398), .C(n_314), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_547), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_535), .B(n_427), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_543), .A2(n_484), .B1(n_413), .B2(n_433), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_535), .B(n_315), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_545), .B(n_474), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_542), .B(n_447), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_545), .Y(n_565) );
INVx3_ASAP7_75t_SL g566 ( .A(n_541), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_546), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_546), .B(n_317), .Y(n_568) );
AND2x2_ASAP7_75t_SL g569 ( .A(n_553), .B(n_338), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_542), .A2(n_410), .B1(n_441), .B2(n_435), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_526), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_549), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_528), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_529), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_544), .B(n_467), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_554), .B(n_484), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_548), .B(n_340), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_536), .B(n_466), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_534), .B(n_540), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_550), .Y(n_580) );
INVx5_ASAP7_75t_L g581 ( .A(n_530), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_553), .A2(n_472), .B1(n_322), .B2(n_327), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_551), .B(n_318), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_538), .A2(n_499), .B(n_329), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_531), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_SL g586 ( .A1(n_532), .A2(n_523), .B(n_522), .C(n_330), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_539), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_539), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_552), .A2(n_331), .B(n_313), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_556), .A2(n_470), .B1(n_473), .B2(n_458), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_572), .B(n_559), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_563), .A2(n_532), .B(n_533), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_576), .B(n_533), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_563), .A2(n_334), .B(n_332), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_590), .B(n_319), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_570), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_561), .B(n_379), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_584), .A2(n_337), .B(n_335), .Y(n_598) );
OAI22x1_ASAP7_75t_L g599 ( .A1(n_566), .A2(n_555), .B1(n_405), .B2(n_358), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_580), .A2(n_588), .B(n_557), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_573), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_569), .A2(n_555), .B1(n_359), .B2(n_360), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_569), .A2(n_371), .B1(n_373), .B2(n_345), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_579), .B(n_377), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_587), .A2(n_578), .B(n_583), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_571), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g607 ( .A1(n_558), .A2(n_381), .B(n_384), .C(n_382), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_577), .Y(n_608) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_565), .Y(n_609) );
BUFx2_ASAP7_75t_L g610 ( .A(n_566), .Y(n_610) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_567), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_561), .B(n_396), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_579), .B(n_396), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_564), .A2(n_574), .B(n_585), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_560), .B(n_320), .Y(n_615) );
BUFx12f_ASAP7_75t_L g616 ( .A(n_581), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_SL g617 ( .A1(n_586), .A2(n_391), .B(n_393), .C(n_386), .Y(n_617) );
O2A1O1Ixp33_ASAP7_75t_L g618 ( .A1(n_558), .A2(n_401), .B(n_421), .C(n_416), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_568), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_581), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_582), .B(n_497), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_581), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_581), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_582), .A2(n_462), .B1(n_325), .B2(n_328), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_575), .B(n_323), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_575), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_589), .A2(n_428), .B(n_430), .C(n_425), .Y(n_627) );
O2A1O1Ixp5_ASAP7_75t_SL g628 ( .A1(n_562), .A2(n_497), .B(n_437), .C(n_446), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_570), .B(n_8), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_620), .Y(n_630) );
AO21x2_ASAP7_75t_L g631 ( .A1(n_598), .A2(n_457), .B(n_440), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_616), .Y(n_632) );
AO21x2_ASAP7_75t_L g633 ( .A1(n_592), .A2(n_468), .B(n_522), .Y(n_633) );
BUFx2_ASAP7_75t_SL g634 ( .A(n_610), .Y(n_634) );
OAI21xp5_ASAP7_75t_L g635 ( .A1(n_600), .A2(n_523), .B(n_403), .Y(n_635) );
OAI21x1_ASAP7_75t_L g636 ( .A1(n_594), .A2(n_426), .B(n_385), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_596), .A2(n_426), .B1(n_436), .B2(n_362), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_591), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_620), .Y(n_639) );
BUFx2_ASAP7_75t_L g640 ( .A(n_620), .Y(n_640) );
OAI21x1_ASAP7_75t_L g641 ( .A1(n_628), .A2(n_426), .B(n_385), .Y(n_641) );
OAI21x1_ASAP7_75t_SL g642 ( .A1(n_605), .A2(n_9), .B(n_10), .Y(n_642) );
CKINVDCx16_ASAP7_75t_R g643 ( .A(n_602), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_626), .B(n_11), .Y(n_644) );
OAI21xp33_ASAP7_75t_SL g645 ( .A1(n_603), .A2(n_11), .B(n_12), .Y(n_645) );
INVx6_ASAP7_75t_SL g646 ( .A(n_613), .Y(n_646) );
CKINVDCx16_ASAP7_75t_R g647 ( .A(n_629), .Y(n_647) );
OAI21x1_ASAP7_75t_SL g648 ( .A1(n_614), .A2(n_13), .B(n_15), .Y(n_648) );
NAND2x1p5_ASAP7_75t_L g649 ( .A(n_595), .B(n_380), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_608), .B(n_13), .Y(n_650) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_623), .B(n_380), .Y(n_651) );
AO21x2_ASAP7_75t_L g652 ( .A1(n_617), .A2(n_492), .B(n_488), .Y(n_652) );
INVx4_ASAP7_75t_L g653 ( .A(n_622), .Y(n_653) );
INVx6_ASAP7_75t_L g654 ( .A(n_609), .Y(n_654) );
NAND2x1_ASAP7_75t_L g655 ( .A(n_606), .B(n_380), .Y(n_655) );
BUFx4f_ASAP7_75t_L g656 ( .A(n_619), .Y(n_656) );
OAI21x1_ASAP7_75t_L g657 ( .A1(n_618), .A2(n_461), .B(n_385), .Y(n_657) );
OAI21x1_ASAP7_75t_L g658 ( .A1(n_612), .A2(n_621), .B(n_601), .Y(n_658) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_599), .Y(n_659) );
INVx4_ASAP7_75t_L g660 ( .A(n_609), .Y(n_660) );
OA21x2_ASAP7_75t_L g661 ( .A1(n_607), .A2(n_627), .B(n_593), .Y(n_661) );
AO21x2_ASAP7_75t_L g662 ( .A1(n_597), .A2(n_492), .B(n_488), .Y(n_662) );
AO21x2_ASAP7_75t_L g663 ( .A1(n_604), .A2(n_492), .B(n_488), .Y(n_663) );
BUFx3_ASAP7_75t_L g664 ( .A(n_609), .Y(n_664) );
AO21x2_ASAP7_75t_L g665 ( .A1(n_604), .A2(n_492), .B(n_488), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_611), .Y(n_666) );
BUFx3_ASAP7_75t_L g667 ( .A(n_611), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_615), .B(n_17), .Y(n_668) );
AO21x2_ASAP7_75t_L g669 ( .A1(n_625), .A2(n_489), .B(n_485), .Y(n_669) );
INVx3_ASAP7_75t_L g670 ( .A(n_611), .Y(n_670) );
BUFx2_ASAP7_75t_SL g671 ( .A(n_624), .Y(n_671) );
NAND2x1_ASAP7_75t_L g672 ( .A(n_620), .B(n_461), .Y(n_672) );
BUFx6f_ASAP7_75t_SL g673 ( .A(n_604), .Y(n_673) );
AO21x2_ASAP7_75t_L g674 ( .A1(n_598), .A2(n_491), .B(n_489), .Y(n_674) );
INVx8_ASAP7_75t_L g675 ( .A(n_616), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_600), .A2(n_339), .B(n_336), .Y(n_676) );
BUFx12f_ASAP7_75t_L g677 ( .A(n_610), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_591), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_616), .Y(n_679) );
AO21x2_ASAP7_75t_L g680 ( .A1(n_598), .A2(n_491), .B(n_489), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_591), .B(n_17), .Y(n_681) );
INVx4_ASAP7_75t_L g682 ( .A(n_616), .Y(n_682) );
BUFx3_ASAP7_75t_L g683 ( .A(n_610), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_620), .B(n_341), .Y(n_684) );
OAI21x1_ASAP7_75t_L g685 ( .A1(n_592), .A2(n_489), .B(n_485), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_647), .B(n_18), .Y(n_686) );
AO21x2_ASAP7_75t_L g687 ( .A1(n_662), .A2(n_491), .B(n_490), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_638), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_638), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_647), .A2(n_343), .B1(n_347), .B2(n_342), .Y(n_690) );
CKINVDCx5p33_ASAP7_75t_R g691 ( .A(n_675), .Y(n_691) );
AO21x1_ASAP7_75t_L g692 ( .A1(n_644), .A2(n_19), .B(n_20), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_678), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_678), .Y(n_694) );
INVx2_ASAP7_75t_SL g695 ( .A(n_675), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_650), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_643), .B(n_20), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_644), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_643), .A2(n_349), .B1(n_350), .B2(n_348), .Y(n_699) );
INVx3_ASAP7_75t_L g700 ( .A(n_653), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_666), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_681), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_671), .A2(n_352), .B1(n_353), .B2(n_351), .Y(n_703) );
INVxp67_ASAP7_75t_L g704 ( .A(n_634), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_673), .A2(n_363), .B1(n_364), .B2(n_354), .Y(n_705) );
AOI21x1_ASAP7_75t_L g706 ( .A1(n_685), .A2(n_491), .B(n_490), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_666), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_683), .Y(n_708) );
INVx2_ASAP7_75t_SL g709 ( .A(n_679), .Y(n_709) );
INVx4_ASAP7_75t_L g710 ( .A(n_682), .Y(n_710) );
INVx3_ASAP7_75t_L g711 ( .A(n_653), .Y(n_711) );
BUFx3_ASAP7_75t_L g712 ( .A(n_677), .Y(n_712) );
OAI21xp5_ASAP7_75t_SL g713 ( .A1(n_668), .A2(n_676), .B(n_649), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_661), .B(n_21), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_642), .Y(n_715) );
INVx3_ASAP7_75t_L g716 ( .A(n_660), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_668), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_648), .Y(n_718) );
INVx2_ASAP7_75t_SL g719 ( .A(n_682), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g720 ( .A(n_632), .B(n_21), .Y(n_720) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_673), .A2(n_367), .B1(n_370), .B2(n_365), .Y(n_721) );
CKINVDCx11_ASAP7_75t_R g722 ( .A(n_639), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_656), .B(n_22), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_661), .A2(n_374), .B1(n_375), .B2(n_372), .Y(n_724) );
BUFx12f_ASAP7_75t_L g725 ( .A(n_659), .Y(n_725) );
INVx6_ASAP7_75t_L g726 ( .A(n_660), .Y(n_726) );
OA21x2_ASAP7_75t_L g727 ( .A1(n_658), .A2(n_383), .B(n_378), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_640), .Y(n_728) );
CKINVDCx11_ASAP7_75t_R g729 ( .A(n_664), .Y(n_729) );
BUFx2_ASAP7_75t_R g730 ( .A(n_667), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_645), .A2(n_389), .B1(n_390), .B2(n_387), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g732 ( .A1(n_645), .A2(n_394), .B1(n_397), .B2(n_392), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_656), .Y(n_733) );
OAI21x1_ASAP7_75t_L g734 ( .A1(n_657), .A2(n_490), .B(n_52), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_630), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_646), .A2(n_400), .B1(n_402), .B2(n_399), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_630), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_684), .Y(n_738) );
BUFx2_ASAP7_75t_SL g739 ( .A(n_670), .Y(n_739) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_654), .Y(n_740) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_676), .A2(n_406), .B1(n_408), .B2(n_404), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_663), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_646), .A2(n_631), .B1(n_637), .B2(n_635), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_663), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_665), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_651), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_665), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_670), .Y(n_748) );
INVx3_ASAP7_75t_L g749 ( .A(n_654), .Y(n_749) );
OR2x6_ASAP7_75t_L g750 ( .A(n_672), .B(n_490), .Y(n_750) );
INVx2_ASAP7_75t_SL g751 ( .A(n_655), .Y(n_751) );
BUFx2_ASAP7_75t_L g752 ( .A(n_669), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_635), .Y(n_753) );
INVx6_ASAP7_75t_L g754 ( .A(n_669), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_633), .B(n_22), .Y(n_755) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_662), .Y(n_756) );
CKINVDCx9p33_ASAP7_75t_R g757 ( .A(n_652), .Y(n_757) );
AO21x1_ASAP7_75t_SL g758 ( .A1(n_652), .A2(n_24), .B(n_25), .Y(n_758) );
AOI22xp33_ASAP7_75t_SL g759 ( .A1(n_633), .A2(n_471), .B1(n_412), .B2(n_414), .Y(n_759) );
INVx2_ASAP7_75t_SL g760 ( .A(n_674), .Y(n_760) );
NAND2x1p5_ASAP7_75t_L g761 ( .A(n_636), .B(n_24), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_641), .Y(n_762) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_674), .Y(n_763) );
CKINVDCx11_ASAP7_75t_R g764 ( .A(n_680), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_680), .Y(n_765) );
AO21x1_ASAP7_75t_SL g766 ( .A1(n_638), .A2(n_25), .B(n_27), .Y(n_766) );
INVxp67_ASAP7_75t_L g767 ( .A(n_634), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_647), .A2(n_415), .B1(n_417), .B2(n_411), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_647), .A2(n_469), .B1(n_465), .B2(n_464), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_647), .A2(n_463), .B1(n_460), .B2(n_459), .Y(n_770) );
AOI21x1_ASAP7_75t_L g771 ( .A1(n_685), .A2(n_419), .B(n_418), .Y(n_771) );
AOI21x1_ASAP7_75t_L g772 ( .A1(n_685), .A2(n_424), .B(n_422), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_638), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_638), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_647), .A2(n_456), .B1(n_454), .B2(n_452), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_638), .Y(n_776) );
AND2x4_ASAP7_75t_L g777 ( .A(n_700), .B(n_27), .Y(n_777) );
NAND3xp33_ASAP7_75t_SL g778 ( .A(n_720), .B(n_431), .C(n_429), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_688), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_694), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_773), .B(n_28), .Y(n_781) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_686), .A2(n_450), .B1(n_449), .B2(n_448), .Y(n_782) );
CKINVDCx16_ASAP7_75t_R g783 ( .A(n_712), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_776), .B(n_28), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_689), .Y(n_785) );
NOR2xp33_ASAP7_75t_R g786 ( .A(n_691), .B(n_29), .Y(n_786) );
NAND3xp33_ASAP7_75t_SL g787 ( .A(n_720), .B(n_438), .C(n_434), .Y(n_787) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_700), .Y(n_788) );
OA21x2_ASAP7_75t_L g789 ( .A1(n_765), .A2(n_443), .B(n_439), .Y(n_789) );
NOR3xp33_ASAP7_75t_SL g790 ( .A(n_713), .B(n_445), .C(n_444), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_695), .Y(n_791) );
INVx4_ASAP7_75t_L g792 ( .A(n_710), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_708), .B(n_29), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_693), .B(n_30), .Y(n_794) );
NOR2xp33_ASAP7_75t_R g795 ( .A(n_710), .B(n_30), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_711), .B(n_31), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_774), .Y(n_797) );
NOR2xp33_ASAP7_75t_R g798 ( .A(n_719), .B(n_31), .Y(n_798) );
NAND2xp33_ASAP7_75t_R g799 ( .A(n_711), .B(n_32), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_696), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_697), .B(n_49), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_728), .B(n_56), .Y(n_802) );
CKINVDCx6p67_ASAP7_75t_R g803 ( .A(n_722), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_698), .Y(n_804) );
BUFx6f_ASAP7_75t_L g805 ( .A(n_729), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_731), .A2(n_60), .B1(n_61), .B2(n_64), .Y(n_806) );
AO21x2_ASAP7_75t_L g807 ( .A1(n_687), .A2(n_66), .B(n_69), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_702), .B(n_71), .Y(n_808) );
AND2x4_ASAP7_75t_L g809 ( .A(n_716), .B(n_78), .Y(n_809) );
CKINVDCx16_ASAP7_75t_R g810 ( .A(n_709), .Y(n_810) );
NAND2xp33_ASAP7_75t_R g811 ( .A(n_723), .B(n_79), .Y(n_811) );
OAI22xp5_ASAP7_75t_SL g812 ( .A1(n_725), .A2(n_81), .B1(n_82), .B2(n_84), .Y(n_812) );
BUFx2_ASAP7_75t_L g813 ( .A(n_704), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_717), .Y(n_814) );
AO31x2_ASAP7_75t_L g815 ( .A1(n_752), .A2(n_85), .A3(n_91), .B(n_92), .Y(n_815) );
NOR3xp33_ASAP7_75t_SL g816 ( .A(n_713), .B(n_93), .C(n_94), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_701), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_707), .Y(n_818) );
NAND2xp33_ASAP7_75t_R g819 ( .A(n_716), .B(n_95), .Y(n_819) );
NOR2x1_ASAP7_75t_SL g820 ( .A(n_766), .B(n_96), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_767), .B(n_305), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_755), .Y(n_822) );
AND2x4_ASAP7_75t_L g823 ( .A(n_735), .B(n_98), .Y(n_823) );
INVx1_ASAP7_75t_SL g824 ( .A(n_730), .Y(n_824) );
A2O1A1Ixp33_ASAP7_75t_L g825 ( .A1(n_731), .A2(n_99), .B(n_101), .C(n_104), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_755), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_737), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_738), .B(n_106), .Y(n_828) );
INVx3_ASAP7_75t_SL g829 ( .A(n_726), .Y(n_829) );
NOR2xp33_ASAP7_75t_R g830 ( .A(n_726), .B(n_107), .Y(n_830) );
OAI211xp5_ASAP7_75t_L g831 ( .A1(n_699), .A2(n_108), .B(n_109), .C(n_110), .Y(n_831) );
INVx4_ASAP7_75t_L g832 ( .A(n_740), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_748), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_732), .A2(n_112), .B1(n_114), .B2(n_115), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_714), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_749), .B(n_117), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_749), .B(n_733), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_692), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_740), .Y(n_839) );
BUFx3_ASAP7_75t_L g840 ( .A(n_740), .Y(n_840) );
AO31x2_ASAP7_75t_L g841 ( .A1(n_742), .A2(n_118), .A3(n_120), .B(n_122), .Y(n_841) );
NOR2xp33_ASAP7_75t_R g842 ( .A(n_764), .B(n_123), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_714), .Y(n_843) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_739), .Y(n_844) );
OAI21xp5_ASAP7_75t_L g845 ( .A1(n_724), .A2(n_124), .B(n_125), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_730), .B(n_126), .Y(n_846) );
OR2x2_ASAP7_75t_L g847 ( .A(n_753), .B(n_127), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_718), .A2(n_129), .B1(n_130), .B2(n_131), .Y(n_848) );
NAND2xp33_ASAP7_75t_R g849 ( .A(n_727), .B(n_132), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_690), .B(n_304), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_715), .Y(n_851) );
NAND3xp33_ASAP7_75t_SL g852 ( .A(n_768), .B(n_135), .C(n_136), .Y(n_852) );
OR2x2_ASAP7_75t_L g853 ( .A(n_746), .B(n_138), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_756), .Y(n_854) );
NAND2xp33_ASAP7_75t_R g855 ( .A(n_727), .B(n_139), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_769), .B(n_141), .Y(n_856) );
AND2x4_ASAP7_75t_SL g857 ( .A(n_770), .B(n_142), .Y(n_857) );
NOR2xp33_ASAP7_75t_R g858 ( .A(n_775), .B(n_144), .Y(n_858) );
OR2x2_ASAP7_75t_L g859 ( .A(n_703), .B(n_298), .Y(n_859) );
NAND2xp33_ASAP7_75t_R g860 ( .A(n_750), .B(n_145), .Y(n_860) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_763), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_743), .A2(n_148), .B1(n_149), .B2(n_153), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_761), .Y(n_863) );
OR2x2_ASAP7_75t_L g864 ( .A(n_703), .B(n_154), .Y(n_864) );
NAND2xp33_ASAP7_75t_R g865 ( .A(n_750), .B(n_156), .Y(n_865) );
OR2x6_ASAP7_75t_L g866 ( .A(n_751), .B(n_157), .Y(n_866) );
BUFx6f_ASAP7_75t_L g867 ( .A(n_750), .Y(n_867) );
CKINVDCx5p33_ASAP7_75t_R g868 ( .A(n_721), .Y(n_868) );
INVxp67_ASAP7_75t_L g869 ( .A(n_758), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g870 ( .A(n_705), .Y(n_870) );
NOR3xp33_ASAP7_75t_SL g871 ( .A(n_762), .B(n_162), .C(n_163), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_759), .B(n_164), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_759), .B(n_165), .Y(n_873) );
NOR2xp33_ASAP7_75t_R g874 ( .A(n_736), .B(n_166), .Y(n_874) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_741), .Y(n_875) );
INVx3_ASAP7_75t_L g876 ( .A(n_754), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_754), .A2(n_168), .B1(n_169), .B2(n_171), .Y(n_877) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_744), .Y(n_878) );
NOR2xp33_ASAP7_75t_R g879 ( .A(n_771), .B(n_172), .Y(n_879) );
BUFx3_ASAP7_75t_L g880 ( .A(n_761), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_760), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_881) );
BUFx3_ASAP7_75t_L g882 ( .A(n_745), .Y(n_882) );
NOR2xp33_ASAP7_75t_R g883 ( .A(n_772), .B(n_176), .Y(n_883) );
INVx3_ASAP7_75t_L g884 ( .A(n_747), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_687), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_757), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_734), .B(n_178), .Y(n_887) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_706), .Y(n_888) );
BUFx2_ASAP7_75t_L g889 ( .A(n_700), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_800), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_779), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_889), .B(n_179), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_810), .B(n_785), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_788), .B(n_181), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_818), .Y(n_895) );
NOR2x1_ASAP7_75t_L g896 ( .A(n_792), .B(n_182), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_793), .B(n_186), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_797), .B(n_188), .Y(n_898) );
NAND3xp33_ASAP7_75t_L g899 ( .A(n_838), .B(n_189), .C(n_190), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_780), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_822), .B(n_191), .Y(n_901) );
BUFx2_ASAP7_75t_L g902 ( .A(n_844), .Y(n_902) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_861), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_817), .B(n_192), .Y(n_904) );
AO21x2_ASAP7_75t_L g905 ( .A1(n_885), .A2(n_193), .B(n_194), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_833), .B(n_813), .Y(n_906) );
OAI21xp33_ASAP7_75t_L g907 ( .A1(n_798), .A2(n_202), .B(n_203), .Y(n_907) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_799), .A2(n_207), .B1(n_208), .B2(n_211), .C(n_214), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_804), .Y(n_909) );
INVx1_ASAP7_75t_SL g910 ( .A(n_829), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_777), .B(n_216), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_826), .B(n_219), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_795), .A2(n_220), .B1(n_221), .B2(n_222), .C(n_223), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_814), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_839), .B(n_224), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_827), .B(n_225), .Y(n_916) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_878), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_854), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_837), .B(n_796), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_777), .B(n_227), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_781), .Y(n_921) );
OA21x2_ASAP7_75t_L g922 ( .A1(n_888), .A2(n_228), .B(n_231), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_784), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_824), .B(n_232), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_840), .B(n_233), .Y(n_925) );
OR2x2_ASAP7_75t_L g926 ( .A(n_783), .B(n_236), .Y(n_926) );
NOR2x1_ASAP7_75t_SL g927 ( .A(n_866), .B(n_237), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_851), .Y(n_928) );
NOR4xp25_ASAP7_75t_SL g929 ( .A(n_819), .B(n_239), .C(n_242), .D(n_243), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_801), .B(n_244), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_794), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_882), .Y(n_932) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_884), .Y(n_933) );
AND2x4_ASAP7_75t_SL g934 ( .A(n_809), .B(n_245), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_843), .Y(n_935) );
AND2x4_ASAP7_75t_SL g936 ( .A(n_809), .B(n_866), .Y(n_936) );
BUFx2_ASAP7_75t_L g937 ( .A(n_830), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_835), .Y(n_938) );
BUFx2_ASAP7_75t_L g939 ( .A(n_842), .Y(n_939) );
OAI21x1_ASAP7_75t_L g940 ( .A1(n_886), .A2(n_247), .B(n_249), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_802), .B(n_252), .Y(n_941) );
AND2x4_ASAP7_75t_L g942 ( .A(n_869), .B(n_253), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_863), .Y(n_943) );
BUFx6f_ASAP7_75t_L g944 ( .A(n_867), .Y(n_944) );
INVx2_ASAP7_75t_L g945 ( .A(n_876), .Y(n_945) );
INVxp67_ASAP7_75t_L g946 ( .A(n_860), .Y(n_946) );
BUFx2_ASAP7_75t_L g947 ( .A(n_832), .Y(n_947) );
BUFx6f_ASAP7_75t_L g948 ( .A(n_867), .Y(n_948) );
BUFx2_ASAP7_75t_L g949 ( .A(n_867), .Y(n_949) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_880), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_841), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_823), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_823), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_841), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_846), .B(n_254), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_816), .B(n_256), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_815), .Y(n_957) );
BUFx2_ASAP7_75t_L g958 ( .A(n_791), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_815), .Y(n_959) );
OR2x2_ASAP7_75t_L g960 ( .A(n_803), .B(n_257), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_828), .B(n_258), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_790), .B(n_259), .Y(n_962) );
OR2x2_ASAP7_75t_L g963 ( .A(n_805), .B(n_261), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_815), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_807), .Y(n_965) );
INVxp67_ASAP7_75t_SL g966 ( .A(n_865), .Y(n_966) );
BUFx3_ASAP7_75t_L g967 ( .A(n_805), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_847), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_853), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_858), .A2(n_264), .B1(n_266), .B2(n_268), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_849), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_808), .Y(n_972) );
INVx2_ASAP7_75t_L g973 ( .A(n_887), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_836), .B(n_270), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_906), .B(n_805), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_935), .B(n_789), .Y(n_976) );
INVx2_ASAP7_75t_L g977 ( .A(n_917), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_917), .B(n_789), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_919), .B(n_820), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_918), .Y(n_980) );
NAND2xp67_ASAP7_75t_L g981 ( .A(n_936), .B(n_857), .Y(n_981) );
AND2x4_ASAP7_75t_L g982 ( .A(n_933), .B(n_936), .Y(n_982) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_903), .Y(n_983) );
AND2x4_ASAP7_75t_L g984 ( .A(n_933), .B(n_871), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_890), .B(n_872), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_895), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_903), .B(n_873), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_932), .B(n_786), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_891), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_900), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_902), .B(n_821), .Y(n_991) );
OR2x2_ASAP7_75t_L g992 ( .A(n_893), .B(n_864), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_909), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_950), .B(n_870), .Y(n_994) );
OR2x2_ASAP7_75t_L g995 ( .A(n_914), .B(n_859), .Y(n_995) );
AND2x4_ASAP7_75t_L g996 ( .A(n_966), .B(n_949), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_938), .B(n_862), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_950), .B(n_874), .Y(n_998) );
OR2x2_ASAP7_75t_L g999 ( .A(n_928), .B(n_778), .Y(n_999) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_943), .B(n_787), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_943), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_971), .B(n_875), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_945), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_945), .B(n_845), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_947), .B(n_806), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_921), .Y(n_1006) );
OR2x2_ASAP7_75t_L g1007 ( .A(n_973), .B(n_868), .Y(n_1007) );
NAND3xp33_ASAP7_75t_L g1008 ( .A(n_913), .B(n_811), .C(n_855), .Y(n_1008) );
BUFx3_ASAP7_75t_L g1009 ( .A(n_958), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_952), .B(n_848), .Y(n_1010) );
INVx2_ASAP7_75t_L g1011 ( .A(n_944), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_923), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_953), .B(n_877), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_931), .Y(n_1014) );
NAND2x1p5_ASAP7_75t_L g1015 ( .A(n_937), .B(n_812), .Y(n_1015) );
INVx2_ASAP7_75t_L g1016 ( .A(n_944), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_969), .Y(n_1017) );
HB1xp67_ASAP7_75t_L g1018 ( .A(n_944), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_946), .B(n_856), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_968), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_973), .B(n_881), .Y(n_1021) );
CKINVDCx14_ASAP7_75t_R g1022 ( .A(n_967), .Y(n_1022) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_910), .B(n_825), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_966), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_967), .B(n_883), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_944), .Y(n_1026) );
OR2x2_ASAP7_75t_L g1027 ( .A(n_946), .B(n_852), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_971), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_983), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_983), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_989), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_982), .B(n_948), .Y(n_1032) );
INVxp67_ASAP7_75t_L g1033 ( .A(n_1028), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_977), .B(n_1020), .Y(n_1034) );
NOR2x1p5_ASAP7_75t_L g1035 ( .A(n_1008), .B(n_960), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_1017), .B(n_948), .Y(n_1036) );
INVx3_ASAP7_75t_L g1037 ( .A(n_982), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1003), .B(n_964), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1024), .B(n_986), .Y(n_1039) );
INVx4_ASAP7_75t_L g1040 ( .A(n_1015), .Y(n_1040) );
OR2x2_ASAP7_75t_L g1041 ( .A(n_987), .B(n_948), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_990), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_975), .B(n_948), .Y(n_1043) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_1009), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1006), .B(n_972), .Y(n_1045) );
AO21x1_ASAP7_75t_L g1046 ( .A1(n_1002), .A2(n_942), .B(n_934), .Y(n_1046) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1001), .Y(n_1047) );
AND2x4_ASAP7_75t_SL g1048 ( .A(n_998), .B(n_942), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1012), .B(n_964), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_993), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_994), .B(n_939), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_996), .B(n_924), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_980), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_1014), .B(n_957), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_987), .B(n_959), .Y(n_1055) );
NAND2xp5_ASAP7_75t_SL g1056 ( .A(n_1015), .B(n_907), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_976), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_1011), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_996), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_979), .B(n_951), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_1022), .B(n_951), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1029), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1057), .B(n_978), .Y(n_1063) );
AOI32xp33_ASAP7_75t_L g1064 ( .A1(n_1040), .A2(n_1002), .A3(n_1025), .B1(n_984), .B2(n_988), .Y(n_1064) );
OA222x2_ASAP7_75t_L g1065 ( .A1(n_1037), .A2(n_992), .B1(n_981), .B2(n_1007), .C1(n_978), .C2(n_995), .Y(n_1065) );
A2O1A1Ixp33_ASAP7_75t_L g1066 ( .A1(n_1056), .A2(n_1008), .B(n_934), .C(n_911), .Y(n_1066) );
NAND3xp33_ASAP7_75t_L g1067 ( .A(n_1040), .B(n_913), .C(n_999), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1030), .Y(n_1068) );
INVx2_ASAP7_75t_SL g1069 ( .A(n_1044), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1059), .B(n_991), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1031), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1042), .Y(n_1072) );
INVx2_ASAP7_75t_SL g1073 ( .A(n_1044), .Y(n_1073) );
NOR2xp67_ASAP7_75t_L g1074 ( .A(n_1040), .B(n_908), .Y(n_1074) );
NAND4xp75_ASAP7_75t_L g1075 ( .A(n_1056), .B(n_896), .C(n_1005), .D(n_1019), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1050), .Y(n_1076) );
O2A1O1Ixp5_ASAP7_75t_L g1077 ( .A1(n_1046), .A2(n_984), .B(n_1019), .C(n_1023), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1059), .B(n_1018), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1053), .Y(n_1079) );
INVx2_ASAP7_75t_SL g1080 ( .A(n_1037), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1058), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_1066), .A2(n_1035), .B1(n_1037), .B2(n_1048), .Y(n_1082) );
INVx1_ASAP7_75t_SL g1083 ( .A(n_1069), .Y(n_1083) );
AOI21xp33_ASAP7_75t_SL g1084 ( .A1(n_1064), .A2(n_926), .B(n_908), .Y(n_1084) );
NOR2xp33_ASAP7_75t_L g1085 ( .A(n_1073), .B(n_1051), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1062), .Y(n_1086) );
AOI31xp33_ASAP7_75t_L g1087 ( .A1(n_1067), .A2(n_1027), .A3(n_1000), .B(n_963), .Y(n_1087) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1081), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1063), .B(n_1033), .Y(n_1089) );
AOI21xp33_ASAP7_75t_SL g1090 ( .A1(n_1067), .A2(n_1033), .B(n_1052), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1065), .B(n_1043), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1068), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_1074), .A2(n_1048), .B1(n_1041), .B2(n_1034), .Y(n_1093) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_1075), .A2(n_1060), .B1(n_1021), .B2(n_1061), .Y(n_1094) );
AOI22xp5_ASAP7_75t_L g1095 ( .A1(n_1070), .A2(n_1055), .B1(n_1010), .B2(n_1013), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1086), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1088), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1091), .B(n_1078), .Y(n_1098) );
OAI22xp5_ASAP7_75t_SL g1099 ( .A1(n_1082), .A2(n_1083), .B1(n_1093), .B2(n_1094), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1083), .B(n_1080), .Y(n_1100) );
OAI211xp5_ASAP7_75t_L g1101 ( .A1(n_1084), .A2(n_1090), .B(n_1095), .C(n_1085), .Y(n_1101) );
CKINVDCx16_ASAP7_75t_R g1102 ( .A(n_1089), .Y(n_1102) );
AOI22xp5_ASAP7_75t_L g1103 ( .A1(n_1092), .A2(n_1045), .B1(n_985), .B2(n_911), .Y(n_1103) );
INVxp67_ASAP7_75t_L g1104 ( .A(n_1087), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1096), .Y(n_1105) );
OA22x2_ASAP7_75t_L g1106 ( .A1(n_1099), .A2(n_1077), .B1(n_1079), .B2(n_1076), .Y(n_1106) );
AOI21xp5_ASAP7_75t_L g1107 ( .A1(n_1104), .A2(n_1077), .B(n_927), .Y(n_1107) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_1102), .B(n_1063), .Y(n_1108) );
OA22x2_ASAP7_75t_L g1109 ( .A1(n_1101), .A2(n_1072), .B1(n_1071), .B2(n_1032), .Y(n_1109) );
AOI221xp5_ASAP7_75t_SL g1110 ( .A1(n_1098), .A2(n_985), .B1(n_1039), .B2(n_955), .C(n_1054), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1108), .Y(n_1111) );
AOI22xp5_ASAP7_75t_L g1112 ( .A1(n_1109), .A2(n_1100), .B1(n_1103), .B2(n_1097), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1110), .B(n_1103), .Y(n_1113) );
NOR2x1_ASAP7_75t_L g1114 ( .A(n_1107), .B(n_922), .Y(n_1114) );
OAI22xp33_ASAP7_75t_L g1115 ( .A1(n_1106), .A2(n_1036), .B1(n_1049), .B2(n_976), .Y(n_1115) );
NAND3xp33_ASAP7_75t_SL g1116 ( .A(n_1112), .B(n_1105), .C(n_929), .Y(n_1116) );
OAI211xp5_ASAP7_75t_L g1117 ( .A1(n_1111), .A2(n_970), .B(n_782), .C(n_962), .Y(n_1117) );
NAND3x1_ASAP7_75t_L g1118 ( .A(n_1114), .B(n_920), .C(n_897), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1113), .B(n_1039), .Y(n_1119) );
NOR2x1_ASAP7_75t_L g1120 ( .A(n_1116), .B(n_1115), .Y(n_1120) );
OA22x2_ASAP7_75t_L g1121 ( .A1(n_1119), .A2(n_1026), .B1(n_1018), .B2(n_1058), .Y(n_1121) );
AOI31xp33_ASAP7_75t_L g1122 ( .A1(n_1117), .A2(n_970), .A3(n_834), .B(n_930), .Y(n_1122) );
CKINVDCx5p33_ASAP7_75t_R g1123 ( .A(n_1121), .Y(n_1123) );
NAND4xp75_ASAP7_75t_L g1124 ( .A(n_1120), .B(n_1122), .C(n_1118), .D(n_925), .Y(n_1124) );
AND2x4_ASAP7_75t_L g1125 ( .A(n_1120), .B(n_1047), .Y(n_1125) );
CKINVDCx16_ASAP7_75t_R g1126 ( .A(n_1125), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1123), .Y(n_1127) );
NOR2xp33_ASAP7_75t_R g1128 ( .A(n_1124), .B(n_272), .Y(n_1128) );
OA22x2_ASAP7_75t_L g1129 ( .A1(n_1127), .A2(n_956), .B1(n_892), .B2(n_894), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1126), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_1128), .A2(n_956), .B1(n_1026), .B2(n_997), .Y(n_1131) );
NAND2x1_ASAP7_75t_L g1132 ( .A(n_1130), .B(n_915), .Y(n_1132) );
OAI31xp33_ASAP7_75t_SL g1133 ( .A1(n_1131), .A2(n_831), .A3(n_899), .B(n_940), .Y(n_1133) );
AOI22x1_ASAP7_75t_L g1134 ( .A1(n_1129), .A2(n_941), .B1(n_974), .B2(n_961), .Y(n_1134) );
AOI21xp5_ASAP7_75t_L g1135 ( .A1(n_1132), .A2(n_850), .B(n_901), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1134), .Y(n_1136) );
AOI32xp33_ASAP7_75t_L g1137 ( .A1(n_1133), .A2(n_916), .A3(n_904), .B1(n_898), .B2(n_912), .Y(n_1137) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_1136), .A2(n_1135), .B1(n_1137), .B2(n_905), .Y(n_1138) );
XNOR2xp5_ASAP7_75t_L g1139 ( .A(n_1138), .B(n_922), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_1139), .A2(n_1016), .B1(n_1004), .B2(n_1047), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1141 ( .A1(n_1140), .A2(n_879), .B1(n_1038), .B2(n_965), .C(n_954), .Y(n_1141) );
AOI22xp5_ASAP7_75t_L g1142 ( .A1(n_1141), .A2(n_922), .B1(n_1038), .B2(n_954), .Y(n_1142) );
endmodule