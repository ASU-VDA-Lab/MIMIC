module real_aes_9124_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_0), .Y(n_458) );
INVx1_ASAP7_75t_L g113 ( .A(n_1), .Y(n_113) );
INVx1_ASAP7_75t_L g485 ( .A(n_2), .Y(n_485) );
INVx1_ASAP7_75t_L g200 ( .A(n_3), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_4), .A2(n_39), .B1(n_161), .B2(n_515), .Y(n_530) );
AOI21xp33_ASAP7_75t_L g168 ( .A1(n_5), .A2(n_142), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_6), .B(n_135), .Y(n_498) );
AND2x6_ASAP7_75t_L g147 ( .A(n_7), .B(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_8), .A2(n_250), .B(n_251), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_9), .B(n_40), .Y(n_114) );
INVx1_ASAP7_75t_L g175 ( .A(n_10), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_11), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g140 ( .A(n_12), .Y(n_140) );
INVx1_ASAP7_75t_L g479 ( .A(n_13), .Y(n_479) );
INVx1_ASAP7_75t_L g256 ( .A(n_14), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_15), .B(n_183), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_16), .B(n_136), .Y(n_556) );
AO32x2_ASAP7_75t_L g528 ( .A1(n_17), .A2(n_135), .A3(n_180), .B1(n_507), .B2(n_529), .Y(n_528) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_18), .A2(n_63), .B1(n_124), .B2(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g125 ( .A(n_18), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_19), .B(n_161), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_20), .B(n_156), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_21), .B(n_136), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_22), .A2(n_51), .B1(n_161), .B2(n_515), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_23), .B(n_142), .Y(n_212) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_24), .A2(n_77), .B1(n_161), .B2(n_183), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_25), .B(n_161), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_26), .B(n_164), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_27), .A2(n_254), .B(n_255), .C(n_257), .Y(n_253) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_28), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_29), .B(n_177), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_30), .B(n_173), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_31), .A2(n_102), .B1(n_115), .B2(n_773), .Y(n_101) );
INVx1_ASAP7_75t_L g189 ( .A(n_32), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_33), .B(n_177), .Y(n_545) );
INVx2_ASAP7_75t_L g145 ( .A(n_34), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_35), .B(n_161), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_36), .B(n_177), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_37), .Y(n_770) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_38), .A2(n_147), .B(n_151), .C(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g187 ( .A(n_41), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_42), .B(n_173), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_43), .B(n_161), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_44), .A2(n_87), .B1(n_219), .B2(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_45), .B(n_161), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_46), .B(n_161), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_47), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_48), .A2(n_70), .B1(n_759), .B2(n_760), .Y(n_758) );
CKINVDCx16_ASAP7_75t_R g760 ( .A(n_48), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_49), .B(n_484), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_50), .B(n_142), .Y(n_244) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_52), .A2(n_61), .B1(n_161), .B2(n_183), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_53), .A2(n_151), .B1(n_183), .B2(n_185), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_54), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_55), .B(n_161), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g197 ( .A(n_56), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_57), .B(n_161), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_58), .A2(n_160), .B(n_172), .C(n_174), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_59), .Y(n_232) );
INVx1_ASAP7_75t_L g170 ( .A(n_60), .Y(n_170) );
INVx1_ASAP7_75t_L g148 ( .A(n_62), .Y(n_148) );
INVx1_ASAP7_75t_L g124 ( .A(n_63), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_64), .B(n_161), .Y(n_486) );
INVx1_ASAP7_75t_L g139 ( .A(n_65), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_66), .Y(n_119) );
AO32x2_ASAP7_75t_L g512 ( .A1(n_67), .A2(n_135), .A3(n_236), .B1(n_507), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g505 ( .A(n_68), .Y(n_505) );
INVx1_ASAP7_75t_L g540 ( .A(n_69), .Y(n_540) );
INVx1_ASAP7_75t_L g759 ( .A(n_70), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_SL g155 ( .A1(n_71), .A2(n_156), .B(n_157), .C(n_160), .Y(n_155) );
INVxp67_ASAP7_75t_L g158 ( .A(n_72), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_73), .B(n_183), .Y(n_541) );
INVx1_ASAP7_75t_L g107 ( .A(n_74), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_75), .Y(n_193) );
INVx1_ASAP7_75t_L g225 ( .A(n_76), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_78), .A2(n_147), .B(n_151), .C(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_79), .B(n_515), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_80), .B(n_183), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_81), .B(n_201), .Y(n_215) );
INVx2_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_83), .B(n_156), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_84), .B(n_183), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_85), .A2(n_147), .B(n_151), .C(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g110 ( .A(n_86), .Y(n_110) );
OR2x2_ASAP7_75t_L g455 ( .A(n_86), .B(n_111), .Y(n_455) );
OR2x2_ASAP7_75t_L g463 ( .A(n_86), .B(n_112), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_88), .A2(n_100), .B1(n_183), .B2(n_184), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_89), .B(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_90), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_91), .A2(n_147), .B(n_151), .C(n_239), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_92), .Y(n_246) );
INVx1_ASAP7_75t_L g154 ( .A(n_93), .Y(n_154) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_94), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_95), .B(n_201), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_96), .B(n_183), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_97), .B(n_135), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_98), .B(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_99), .A2(n_142), .B(n_149), .Y(n_141) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx12_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g774 ( .A(n_105), .Y(n_774) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g769 ( .A(n_109), .Y(n_769) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g466 ( .A(n_110), .B(n_112), .Y(n_466) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OAI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B(n_459), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g772 ( .A(n_118), .Y(n_772) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_452), .B(n_456), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_126), .B2(n_451), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g451 ( .A(n_126), .Y(n_451) );
INVx1_ASAP7_75t_SL g464 ( .A(n_126), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_126), .A2(n_762), .B1(n_764), .B2(n_765), .Y(n_761) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND4x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_369), .C(n_416), .D(n_436), .Y(n_127) );
NOR3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_299), .C(n_324), .Y(n_128) );
OAI211xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_207), .B(n_259), .C(n_289), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_178), .Y(n_131) );
INVx3_ASAP7_75t_SL g341 ( .A(n_132), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_132), .B(n_272), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_132), .B(n_194), .Y(n_422) );
AND2x2_ASAP7_75t_L g445 ( .A(n_132), .B(n_311), .Y(n_445) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_166), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g263 ( .A(n_134), .B(n_167), .Y(n_263) );
INVx3_ASAP7_75t_L g276 ( .A(n_134), .Y(n_276) );
AND2x2_ASAP7_75t_L g281 ( .A(n_134), .B(n_166), .Y(n_281) );
OR2x2_ASAP7_75t_L g332 ( .A(n_134), .B(n_273), .Y(n_332) );
BUFx2_ASAP7_75t_L g352 ( .A(n_134), .Y(n_352) );
AND2x2_ASAP7_75t_L g362 ( .A(n_134), .B(n_273), .Y(n_362) );
AND2x2_ASAP7_75t_L g368 ( .A(n_134), .B(n_179), .Y(n_368) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_141), .B(n_163), .Y(n_134) );
INVx4_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_135), .A2(n_491), .B(n_498), .Y(n_490) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_137), .B(n_138), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx2_ASAP7_75t_L g250 ( .A(n_142), .Y(n_250) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_147), .Y(n_142) );
NAND2x1p5_ASAP7_75t_L g191 ( .A(n_143), .B(n_147), .Y(n_191) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx1_ASAP7_75t_L g484 ( .A(n_144), .Y(n_484) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g152 ( .A(n_145), .Y(n_152) );
INVx1_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
INVx1_ASAP7_75t_L g153 ( .A(n_146), .Y(n_153) );
INVx1_ASAP7_75t_L g156 ( .A(n_146), .Y(n_156) );
INVx3_ASAP7_75t_L g159 ( .A(n_146), .Y(n_159) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_146), .Y(n_186) );
INVx4_ASAP7_75t_SL g162 ( .A(n_147), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_147), .A2(n_478), .B(n_482), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_147), .A2(n_492), .B(n_495), .Y(n_491) );
BUFx3_ASAP7_75t_L g507 ( .A(n_147), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_147), .A2(n_520), .B(n_524), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_147), .A2(n_539), .B(n_542), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_154), .B(n_155), .C(n_162), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_150), .A2(n_162), .B(n_170), .C(n_171), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_150), .A2(n_162), .B(n_252), .C(n_253), .Y(n_251) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_152), .Y(n_161) );
BUFx3_ASAP7_75t_L g219 ( .A(n_152), .Y(n_219) );
INVx1_ASAP7_75t_L g515 ( .A(n_152), .Y(n_515) );
INVx1_ASAP7_75t_L g523 ( .A(n_156), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_159), .B(n_175), .Y(n_174) );
INVx5_ASAP7_75t_L g201 ( .A(n_159), .Y(n_201) );
OAI22xp5_ASAP7_75t_SL g513 ( .A1(n_159), .A2(n_173), .B1(n_514), .B2(n_516), .Y(n_513) );
O2A1O1Ixp5_ASAP7_75t_SL g539 ( .A1(n_160), .A2(n_201), .B(n_540), .C(n_541), .Y(n_539) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_161), .Y(n_243) );
OAI22xp33_ASAP7_75t_L g181 ( .A1(n_162), .A2(n_182), .B1(n_190), .B2(n_191), .Y(n_181) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_164), .A2(n_168), .B(n_176), .Y(n_167) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_SL g221 ( .A(n_165), .B(n_222), .Y(n_221) );
AO21x1_ASAP7_75t_L g551 ( .A1(n_165), .A2(n_552), .B(n_555), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g570 ( .A(n_165), .B(n_507), .C(n_552), .Y(n_570) );
INVx1_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_167), .B(n_273), .Y(n_287) );
INVx2_ASAP7_75t_L g297 ( .A(n_167), .Y(n_297) );
AND2x2_ASAP7_75t_L g310 ( .A(n_167), .B(n_276), .Y(n_310) );
OR2x2_ASAP7_75t_L g321 ( .A(n_167), .B(n_273), .Y(n_321) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_167), .B(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g379 ( .A(n_167), .Y(n_379) );
AND2x2_ASAP7_75t_L g425 ( .A(n_167), .B(n_179), .Y(n_425) );
O2A1O1Ixp5_ASAP7_75t_L g504 ( .A1(n_172), .A2(n_483), .B(n_505), .C(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_172), .A2(n_525), .B(n_526), .Y(n_524) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g242 ( .A(n_173), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_173), .A2(n_487), .B1(n_530), .B2(n_531), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_173), .A2(n_487), .B1(n_553), .B2(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g206 ( .A(n_177), .Y(n_206) );
INVx2_ASAP7_75t_L g236 ( .A(n_177), .Y(n_236) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_177), .A2(n_249), .B(n_258), .Y(n_248) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_177), .A2(n_519), .B(n_527), .Y(n_518) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_177), .A2(n_538), .B(n_545), .Y(n_537) );
INVx3_ASAP7_75t_SL g298 ( .A(n_178), .Y(n_298) );
OR2x2_ASAP7_75t_L g351 ( .A(n_178), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_194), .Y(n_178) );
INVx3_ASAP7_75t_L g273 ( .A(n_179), .Y(n_273) );
AND2x2_ASAP7_75t_L g340 ( .A(n_179), .B(n_195), .Y(n_340) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_179), .Y(n_408) );
AOI33xp33_ASAP7_75t_L g412 ( .A1(n_179), .A2(n_341), .A3(n_348), .B1(n_357), .B2(n_413), .B3(n_414), .Y(n_412) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_192), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_180), .B(n_193), .Y(n_192) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_180), .A2(n_196), .B(n_204), .Y(n_195) );
INVx2_ASAP7_75t_L g220 ( .A(n_180), .Y(n_220) );
INVx2_ASAP7_75t_L g203 ( .A(n_183), .Y(n_203) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OAI22xp5_ASAP7_75t_SL g185 ( .A1(n_186), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_185) );
INVx2_ASAP7_75t_L g188 ( .A(n_186), .Y(n_188) );
INVx4_ASAP7_75t_L g254 ( .A(n_186), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g196 ( .A1(n_191), .A2(n_197), .B(n_198), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_191), .A2(n_225), .B(n_226), .Y(n_224) );
INVx1_ASAP7_75t_L g261 ( .A(n_194), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_194), .B(n_276), .Y(n_275) );
NOR3xp33_ASAP7_75t_L g335 ( .A(n_194), .B(n_336), .C(n_338), .Y(n_335) );
AND2x2_ASAP7_75t_L g361 ( .A(n_194), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_194), .B(n_368), .Y(n_371) );
AND2x2_ASAP7_75t_L g424 ( .A(n_194), .B(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g280 ( .A(n_195), .Y(n_280) );
OR2x2_ASAP7_75t_L g374 ( .A(n_195), .B(n_273), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_202), .C(n_203), .Y(n_199) );
INVx2_ASAP7_75t_L g487 ( .A(n_201), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_201), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_201), .A2(n_502), .B(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_203), .A2(n_479), .B(n_480), .C(n_481), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_206), .B(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_206), .B(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_233), .Y(n_207) );
AOI32xp33_ASAP7_75t_L g325 ( .A1(n_208), .A2(n_326), .A3(n_328), .B1(n_330), .B2(n_333), .Y(n_325) );
NOR2xp67_ASAP7_75t_L g398 ( .A(n_208), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g428 ( .A(n_208), .Y(n_428) );
INVx4_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g360 ( .A(n_209), .B(n_344), .Y(n_360) );
AND2x2_ASAP7_75t_L g380 ( .A(n_209), .B(n_306), .Y(n_380) );
AND2x2_ASAP7_75t_L g448 ( .A(n_209), .B(n_366), .Y(n_448) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_223), .Y(n_209) );
INVx3_ASAP7_75t_L g269 ( .A(n_210), .Y(n_269) );
AND2x2_ASAP7_75t_L g283 ( .A(n_210), .B(n_267), .Y(n_283) );
OR2x2_ASAP7_75t_L g288 ( .A(n_210), .B(n_266), .Y(n_288) );
INVx1_ASAP7_75t_L g295 ( .A(n_210), .Y(n_295) );
AND2x2_ASAP7_75t_L g303 ( .A(n_210), .B(n_277), .Y(n_303) );
AND2x2_ASAP7_75t_L g305 ( .A(n_210), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_210), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g358 ( .A(n_210), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_210), .B(n_443), .Y(n_442) );
OR2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_221), .Y(n_210) );
AOI21xp5_ASAP7_75t_SL g211 ( .A1(n_212), .A2(n_213), .B(n_220), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_217), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_217), .A2(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g257 ( .A(n_219), .Y(n_257) );
INVx1_ASAP7_75t_L g230 ( .A(n_220), .Y(n_230) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_220), .A2(n_477), .B(n_488), .Y(n_476) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_220), .A2(n_500), .B(n_508), .Y(n_499) );
INVx2_ASAP7_75t_L g267 ( .A(n_223), .Y(n_267) );
AND2x2_ASAP7_75t_L g313 ( .A(n_223), .B(n_234), .Y(n_313) );
AND2x2_ASAP7_75t_L g323 ( .A(n_223), .B(n_248), .Y(n_323) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_230), .B(n_231), .Y(n_223) );
INVx2_ASAP7_75t_L g443 ( .A(n_233), .Y(n_443) );
OR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_247), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_234), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g284 ( .A(n_234), .Y(n_284) );
AND2x2_ASAP7_75t_L g328 ( .A(n_234), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g344 ( .A(n_234), .B(n_307), .Y(n_344) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g292 ( .A(n_235), .Y(n_292) );
AND2x2_ASAP7_75t_L g306 ( .A(n_235), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g357 ( .A(n_235), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_235), .B(n_267), .Y(n_389) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_245), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_243), .Y(n_239) );
AND2x2_ASAP7_75t_L g268 ( .A(n_247), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g329 ( .A(n_247), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_247), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g366 ( .A(n_247), .Y(n_366) );
INVx1_ASAP7_75t_L g399 ( .A(n_247), .Y(n_399) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g277 ( .A(n_248), .B(n_267), .Y(n_277) );
INVx1_ASAP7_75t_L g307 ( .A(n_248), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_254), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g481 ( .A(n_254), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_254), .A2(n_543), .B(n_544), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_264), .B1(n_270), .B2(n_277), .C(n_278), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_261), .B(n_281), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_261), .B(n_344), .Y(n_421) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_263), .B(n_311), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_263), .B(n_272), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_263), .B(n_286), .Y(n_415) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g337 ( .A(n_267), .Y(n_337) );
AND2x2_ASAP7_75t_L g312 ( .A(n_268), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g390 ( .A(n_268), .Y(n_390) );
AND2x2_ASAP7_75t_L g322 ( .A(n_269), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_269), .B(n_292), .Y(n_338) );
AND2x2_ASAP7_75t_L g402 ( .A(n_269), .B(n_328), .Y(n_402) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g311 ( .A(n_273), .B(n_280), .Y(n_311) );
AND2x2_ASAP7_75t_L g407 ( .A(n_274), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_276), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_277), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_277), .B(n_284), .Y(n_372) );
AND2x2_ASAP7_75t_L g392 ( .A(n_277), .B(n_292), .Y(n_392) );
AND2x2_ASAP7_75t_L g413 ( .A(n_277), .B(n_357), .Y(n_413) );
OAI32xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_282), .A3(n_284), .B1(n_285), .B2(n_288), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_SL g286 ( .A(n_280), .Y(n_286) );
NAND2x1_ASAP7_75t_L g327 ( .A(n_280), .B(n_310), .Y(n_327) );
OR2x2_ASAP7_75t_L g331 ( .A(n_280), .B(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_280), .B(n_379), .Y(n_432) );
INVx1_ASAP7_75t_L g300 ( .A(n_281), .Y(n_300) );
OAI221xp5_ASAP7_75t_SL g418 ( .A1(n_282), .A2(n_373), .B1(n_419), .B2(n_422), .C(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g290 ( .A(n_283), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g333 ( .A(n_283), .B(n_306), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_283), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g411 ( .A(n_283), .B(n_344), .Y(n_411) );
INVxp67_ASAP7_75t_L g347 ( .A(n_284), .Y(n_347) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g417 ( .A(n_286), .B(n_404), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_286), .B(n_367), .Y(n_440) );
INVx1_ASAP7_75t_L g315 ( .A(n_288), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_288), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g433 ( .A(n_288), .B(n_434), .Y(n_433) );
OAI21xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_293), .B(n_296), .Y(n_289) );
AND2x2_ASAP7_75t_L g302 ( .A(n_291), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g386 ( .A(n_295), .B(n_306), .Y(n_386) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g404 ( .A(n_297), .B(n_362), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_297), .B(n_361), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_298), .B(n_310), .Y(n_384) );
OAI211xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B(n_304), .C(n_314), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_300), .A2(n_335), .B1(n_339), .B2(n_342), .C(n_345), .Y(n_334) );
AOI31xp33_ASAP7_75t_L g429 ( .A1(n_300), .A2(n_430), .A3(n_431), .B(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_308), .B1(n_310), .B2(n_312), .Y(n_304) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g430 ( .A(n_310), .Y(n_430) );
INVx1_ASAP7_75t_L g393 ( .A(n_311), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_L g436 ( .A1(n_313), .A2(n_437), .B(n_439), .C(n_441), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_318), .B2(n_322), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_319), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI221xp5_ASAP7_75t_SL g409 ( .A1(n_321), .A2(n_355), .B1(n_374), .B2(n_410), .C(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g405 ( .A(n_322), .Y(n_405) );
INVx1_ASAP7_75t_L g359 ( .A(n_323), .Y(n_359) );
NAND3xp33_ASAP7_75t_SL g324 ( .A(n_325), .B(n_334), .C(n_349), .Y(n_324) );
OAI21xp33_ASAP7_75t_L g375 ( .A1(n_326), .A2(n_376), .B(n_380), .Y(n_375) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_328), .B(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g435 ( .A(n_329), .Y(n_435) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g373 ( .A(n_336), .B(n_356), .Y(n_373) );
INVx1_ASAP7_75t_L g348 ( .A(n_337), .Y(n_348) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g346 ( .A(n_340), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_340), .B(n_378), .Y(n_377) );
NOR4xp25_ASAP7_75t_L g345 ( .A(n_341), .B(n_346), .C(n_347), .D(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI222xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_354), .B1(n_360), .B2(n_361), .C1(n_363), .C2(n_367), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g447 ( .A(n_351), .Y(n_447) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_359), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_363), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI21xp5_ASAP7_75t_SL g423 ( .A1(n_368), .A2(n_424), .B(n_426), .Y(n_423) );
NOR4xp25_ASAP7_75t_L g369 ( .A(n_370), .B(n_381), .C(n_394), .D(n_409), .Y(n_369) );
OAI221xp5_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_372), .B1(n_373), .B2(n_374), .C(n_375), .Y(n_370) );
INVx1_ASAP7_75t_L g450 ( .A(n_371), .Y(n_450) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_378), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
OAI222xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_385), .B1(n_387), .B2(n_388), .C1(n_391), .C2(n_393), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_386), .A2(n_417), .B(n_418), .C(n_429), .Y(n_416) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
OAI222xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_400), .B1(n_401), .B2(n_403), .C1(n_405), .C2(n_406), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_411), .A2(n_414), .B1(n_447), .B2(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI211xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_444), .B(n_446), .C(n_449), .Y(n_441) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g457 ( .A(n_455), .Y(n_457) );
OAI21xp5_ASAP7_75t_SL g459 ( .A1(n_456), .A2(n_460), .B(n_771), .Y(n_459) );
NOR2xp33_ASAP7_75t_SL g456 ( .A(n_457), .B(n_458), .Y(n_456) );
OAI222xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_758), .B1(n_761), .B2(n_766), .C1(n_767), .C2(n_770), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_464), .B1(n_465), .B2(n_467), .Y(n_461) );
INVx2_ASAP7_75t_L g763 ( .A(n_462), .Y(n_763) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx6_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g764 ( .A(n_466), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_467), .Y(n_765) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_468), .B(n_724), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_628), .C(n_712), .Y(n_468) );
NAND4xp25_ASAP7_75t_L g469 ( .A(n_470), .B(n_571), .C(n_593), .D(n_609), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_509), .B1(n_532), .B2(n_550), .C(n_557), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_489), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_473), .B(n_550), .Y(n_583) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_473), .B(n_611), .C(n_624), .D(n_626), .Y(n_623) );
INVxp67_ASAP7_75t_L g740 ( .A(n_473), .Y(n_740) );
INVx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g622 ( .A(n_474), .B(n_560), .Y(n_622) );
AND2x2_ASAP7_75t_L g646 ( .A(n_474), .B(n_489), .Y(n_646) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g613 ( .A(n_475), .B(n_549), .Y(n_613) );
AND2x2_ASAP7_75t_L g653 ( .A(n_475), .B(n_634), .Y(n_653) );
AND2x2_ASAP7_75t_L g670 ( .A(n_475), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_475), .B(n_490), .Y(n_694) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g548 ( .A(n_476), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g565 ( .A(n_476), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g577 ( .A(n_476), .B(n_490), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_476), .B(n_499), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B(n_486), .C(n_487), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_487), .A2(n_496), .B(n_497), .Y(n_495) );
AND2x2_ASAP7_75t_L g580 ( .A(n_489), .B(n_581), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_489), .A2(n_630), .B1(n_633), .B2(n_635), .C(n_639), .Y(n_629) );
AND2x2_ASAP7_75t_L g688 ( .A(n_489), .B(n_653), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_489), .B(n_670), .Y(n_722) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
INVx3_ASAP7_75t_L g549 ( .A(n_490), .Y(n_549) );
AND2x2_ASAP7_75t_L g597 ( .A(n_490), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g651 ( .A(n_490), .B(n_566), .Y(n_651) );
AND2x2_ASAP7_75t_L g709 ( .A(n_490), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g550 ( .A(n_499), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g566 ( .A(n_499), .Y(n_566) );
INVx1_ASAP7_75t_L g621 ( .A(n_499), .Y(n_621) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_499), .Y(n_627) );
AND2x2_ASAP7_75t_L g672 ( .A(n_499), .B(n_549), .Y(n_672) );
OR2x2_ASAP7_75t_L g711 ( .A(n_499), .B(n_551), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_504), .B(n_507), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_509), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_517), .Y(n_509) );
AND2x2_ASAP7_75t_L g707 ( .A(n_510), .B(n_704), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_510), .B(n_689), .Y(n_739) );
BUFx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g638 ( .A(n_511), .B(n_562), .Y(n_638) );
AND2x2_ASAP7_75t_L g687 ( .A(n_511), .B(n_535), .Y(n_687) );
INVx1_ASAP7_75t_L g733 ( .A(n_511), .Y(n_733) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_512), .Y(n_547) );
AND2x2_ASAP7_75t_L g588 ( .A(n_512), .B(n_562), .Y(n_588) );
INVx1_ASAP7_75t_L g605 ( .A(n_512), .Y(n_605) );
AND2x2_ASAP7_75t_L g611 ( .A(n_512), .B(n_528), .Y(n_611) );
AND2x2_ASAP7_75t_L g679 ( .A(n_517), .B(n_587), .Y(n_679) );
INVx2_ASAP7_75t_L g744 ( .A(n_517), .Y(n_744) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .Y(n_517) );
AND2x2_ASAP7_75t_L g561 ( .A(n_518), .B(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g574 ( .A(n_518), .B(n_536), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_518), .B(n_535), .Y(n_602) );
INVx1_ASAP7_75t_L g608 ( .A(n_518), .Y(n_608) );
INVx1_ASAP7_75t_L g625 ( .A(n_518), .Y(n_625) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_518), .Y(n_637) );
INVx2_ASAP7_75t_L g705 ( .A(n_518), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_523), .Y(n_520) );
INVx2_ASAP7_75t_L g562 ( .A(n_528), .Y(n_562) );
BUFx2_ASAP7_75t_L g659 ( .A(n_528), .Y(n_659) );
AND2x2_ASAP7_75t_L g704 ( .A(n_528), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_546), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_534), .B(n_641), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_534), .A2(n_703), .B(n_717), .Y(n_727) );
AND2x2_ASAP7_75t_L g752 ( .A(n_534), .B(n_638), .Y(n_752) );
BUFx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g674 ( .A(n_536), .Y(n_674) );
AND2x2_ASAP7_75t_L g703 ( .A(n_536), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_537), .Y(n_587) );
INVx2_ASAP7_75t_L g606 ( .A(n_537), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_537), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx2_ASAP7_75t_L g560 ( .A(n_547), .Y(n_560) );
OR2x2_ASAP7_75t_L g573 ( .A(n_547), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g641 ( .A(n_547), .B(n_637), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_547), .B(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g742 ( .A(n_547), .B(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_547), .B(n_679), .Y(n_754) );
AND2x2_ASAP7_75t_L g633 ( .A(n_548), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g656 ( .A(n_548), .B(n_550), .Y(n_656) );
INVx2_ASAP7_75t_L g568 ( .A(n_549), .Y(n_568) );
AND2x2_ASAP7_75t_L g596 ( .A(n_549), .B(n_569), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_549), .B(n_621), .Y(n_677) );
AND2x2_ASAP7_75t_L g591 ( .A(n_550), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g738 ( .A(n_550), .Y(n_738) );
AND2x2_ASAP7_75t_L g750 ( .A(n_550), .B(n_613), .Y(n_750) );
AND2x2_ASAP7_75t_L g576 ( .A(n_551), .B(n_566), .Y(n_576) );
INVx1_ASAP7_75t_L g671 ( .A(n_551), .Y(n_671) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_L g569 ( .A(n_556), .B(n_570), .Y(n_569) );
INVxp67_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_563), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_560), .B(n_607), .Y(n_616) );
OR2x2_ASAP7_75t_L g748 ( .A(n_560), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g665 ( .A(n_561), .B(n_606), .Y(n_665) );
AND2x2_ASAP7_75t_L g673 ( .A(n_561), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g732 ( .A(n_561), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g756 ( .A(n_561), .B(n_603), .Y(n_756) );
NOR2xp67_ASAP7_75t_L g714 ( .A(n_562), .B(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g743 ( .A(n_562), .B(n_606), .Y(n_743) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2x1p5_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
AND2x2_ASAP7_75t_L g595 ( .A(n_565), .B(n_596), .Y(n_595) );
INVxp67_ASAP7_75t_L g757 ( .A(n_565), .Y(n_757) );
NOR2x1_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g592 ( .A(n_568), .Y(n_592) );
AND2x2_ASAP7_75t_L g643 ( .A(n_568), .B(n_576), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_568), .B(n_711), .Y(n_737) );
INVx2_ASAP7_75t_L g582 ( .A(n_569), .Y(n_582) );
INVx3_ASAP7_75t_L g634 ( .A(n_569), .Y(n_634) );
OR2x2_ASAP7_75t_L g662 ( .A(n_569), .B(n_663), .Y(n_662) );
AOI311xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_575), .A3(n_577), .B(n_578), .C(n_589), .Y(n_571) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_572), .A2(n_610), .B(n_612), .C(n_614), .Y(n_609) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_SL g594 ( .A(n_574), .Y(n_594) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g612 ( .A(n_576), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_576), .B(n_592), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_576), .B(n_577), .Y(n_745) );
AND2x2_ASAP7_75t_L g667 ( .A(n_577), .B(n_581), .Y(n_667) );
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_583), .B(n_584), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g725 ( .A(n_581), .B(n_613), .Y(n_725) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_582), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g619 ( .A(n_582), .Y(n_619) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
AND2x2_ASAP7_75t_L g610 ( .A(n_586), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g655 ( .A(n_588), .Y(n_655) );
AND2x4_ASAP7_75t_L g717 ( .A(n_588), .B(n_686), .Y(n_717) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_591), .A2(n_657), .B1(n_669), .B2(n_673), .C1(n_675), .C2(n_679), .Y(n_668) );
A2O1A1Ixp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B(n_597), .C(n_600), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_594), .B(n_638), .Y(n_661) );
INVx1_ASAP7_75t_L g683 ( .A(n_596), .Y(n_683) );
INVx1_ASAP7_75t_L g617 ( .A(n_598), .Y(n_617) );
OR2x2_ASAP7_75t_L g682 ( .A(n_599), .B(n_683), .Y(n_682) );
OAI21xp33_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_603), .B(n_607), .Y(n_600) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_601), .B(n_619), .C(n_620), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_601), .A2(n_638), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_605), .Y(n_658) );
AND2x2_ASAP7_75t_SL g624 ( .A(n_606), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g715 ( .A(n_606), .Y(n_715) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_606), .Y(n_731) );
INVx2_ASAP7_75t_L g689 ( .A(n_607), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_611), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g663 ( .A(n_613), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_617), .B1(n_618), .B2(n_622), .C(n_623), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_617), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g751 ( .A(n_617), .Y(n_751) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g632 ( .A(n_624), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_624), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g690 ( .A(n_624), .B(n_638), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_624), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g723 ( .A(n_624), .B(n_658), .Y(n_723) );
BUFx3_ASAP7_75t_L g686 ( .A(n_625), .Y(n_686) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND5xp2_ASAP7_75t_L g628 ( .A(n_629), .B(n_647), .C(n_668), .D(n_680), .E(n_695), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI32xp33_ASAP7_75t_L g720 ( .A1(n_632), .A2(n_659), .A3(n_675), .B1(n_721), .B2(n_723), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_634), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g644 ( .A(n_638), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B1(n_644), .B2(n_645), .Y(n_639) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_654), .B1(n_656), .B2(n_657), .C(n_660), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g719 ( .A(n_651), .B(n_670), .Y(n_719) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_656), .A2(n_717), .B1(n_735), .B2(n_740), .C(n_741), .Y(n_734) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx2_ASAP7_75t_L g700 ( .A(n_659), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_664), .B2(n_666), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g678 ( .A(n_670), .Y(n_678) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B1(n_688), .B2(n_689), .C1(n_690), .C2(n_691), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI22xp33_ASAP7_75t_L g735 ( .A1(n_689), .A2(n_736), .B1(n_738), .B2(n_739), .Y(n_735) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B(n_701), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_706), .B(n_708), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g749 ( .A(n_704), .Y(n_749) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_716), .B(n_718), .C(n_720), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AOI211xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B(n_728), .C(n_753), .Y(n_724) );
CKINVDCx16_ASAP7_75t_R g729 ( .A(n_725), .Y(n_729) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI211xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B(n_734), .C(n_746), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
AOI21xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_744), .B(n_745), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AOI21xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B(n_757), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g766 ( .A(n_758), .Y(n_766) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
endmodule