module fake_jpeg_6386_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_15),
.B(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_14),
.B(n_0),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_20),
.A2(n_8),
.B1(n_10),
.B2(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_21),
.B(n_22),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_19),
.B(n_17),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_30),
.B1(n_9),
.B2(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_12),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_12),
.B1(n_17),
.B2(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_1),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_12),
.B1(n_20),
.B2(n_11),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_1),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_2),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_38),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_18),
.C(n_16),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_34),
.B(n_18),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_47),
.C(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

AOI322xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_41),
.A3(n_45),
.B1(n_40),
.B2(n_5),
.C1(n_7),
.C2(n_11),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_42),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_7),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_53),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_52),
.C(n_50),
.Y(n_56)
);

OAI321xp33_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_54),
.A3(n_27),
.B1(n_9),
.B2(n_3),
.C(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_9),
.Y(n_59)
);


endmodule