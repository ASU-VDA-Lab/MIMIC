module real_aes_17873_n_329 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_329);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_329;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1744;
wire n_1044;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_1745;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_1740;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_1749;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_1192;
wire n_518;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1280;
wire n_394;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI221xp5_ASAP7_75t_L g998 ( .A1(n_0), .A2(n_92), .B1(n_646), .B2(n_689), .C(n_999), .Y(n_998) );
AOI22xp33_ASAP7_75t_SL g1013 ( .A1(n_0), .A2(n_221), .B1(n_1014), .B2(n_1016), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_1), .A2(n_260), .B1(n_520), .B2(n_942), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1220 ( .A1(n_1), .A2(n_230), .B1(n_604), .B2(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g343 ( .A(n_2), .Y(n_343) );
AND2x2_ASAP7_75t_L g368 ( .A(n_2), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g404 ( .A(n_2), .B(n_236), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_2), .B(n_353), .Y(n_635) );
INVx1_ASAP7_75t_L g681 ( .A(n_3), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_3), .A2(n_67), .B1(n_545), .B2(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g891 ( .A(n_4), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_4), .A2(n_11), .B1(n_624), .B2(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g935 ( .A(n_5), .Y(n_935) );
OAI221xp5_ASAP7_75t_L g960 ( .A1(n_5), .A2(n_130), .B1(n_775), .B2(n_961), .C(n_963), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g1741 ( .A1(n_6), .A2(n_1742), .B1(n_1743), .B2(n_1744), .Y(n_1741) );
CKINVDCx5p33_ASAP7_75t_R g1744 ( .A(n_6), .Y(n_1744) );
INVx1_ASAP7_75t_L g1172 ( .A(n_7), .Y(n_1172) );
INVx1_ASAP7_75t_L g988 ( .A(n_8), .Y(n_988) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_8), .A2(n_79), .B1(n_947), .B2(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g661 ( .A(n_9), .Y(n_661) );
INVx1_ASAP7_75t_L g1051 ( .A(n_10), .Y(n_1051) );
OA222x2_ASAP7_75t_L g1064 ( .A1(n_10), .A2(n_132), .B1(n_156), .B2(n_617), .C1(n_664), .C2(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g902 ( .A(n_11), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g1502 ( .A1(n_12), .A2(n_180), .B1(n_1476), .B2(n_1490), .Y(n_1502) );
INVxp67_ASAP7_75t_SL g1160 ( .A(n_13), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_13), .A2(n_102), .B1(n_515), .B2(n_1040), .Y(n_1190) );
INVx1_ASAP7_75t_L g1158 ( .A(n_14), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_14), .A2(n_149), .B1(n_563), .B2(n_701), .Y(n_1191) );
AOI22xp33_ASAP7_75t_SL g1208 ( .A1(n_15), .A2(n_187), .B1(n_571), .B2(n_938), .Y(n_1208) );
AOI221xp5_ASAP7_75t_L g1219 ( .A1(n_15), .A2(n_100), .B1(n_412), .B2(n_783), .C(n_1071), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_16), .A2(n_76), .B1(n_1476), .B2(n_1478), .Y(n_1494) );
AOI22xp33_ASAP7_75t_L g1591 ( .A1(n_17), .A2(n_316), .B1(n_1468), .B2(n_1473), .Y(n_1591) );
OAI221xp5_ASAP7_75t_L g544 ( .A1(n_18), .A2(n_321), .B1(n_545), .B2(n_547), .C(n_549), .Y(n_544) );
OAI21xp33_ASAP7_75t_SL g616 ( .A1(n_18), .A2(n_617), .B(n_618), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g1398 ( .A1(n_19), .A2(n_59), .B1(n_1041), .B2(n_1276), .Y(n_1398) );
AOI221xp5_ASAP7_75t_L g1413 ( .A1(n_19), .A2(n_294), .B1(n_688), .B2(n_915), .C(n_1414), .Y(n_1413) );
AOI221xp5_ASAP7_75t_L g979 ( .A1(n_20), .A2(n_78), .B1(n_646), .B2(n_980), .C(n_982), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g1022 ( .A1(n_20), .A2(n_177), .B1(n_515), .B2(n_516), .Y(n_1022) );
INVx2_ASAP7_75t_L g459 ( .A(n_21), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_22), .A2(n_149), .B1(n_604), .B2(n_676), .Y(n_1169) );
AOI22xp5_ASAP7_75t_L g1192 ( .A1(n_22), .A2(n_292), .B1(n_701), .B2(n_709), .Y(n_1192) );
CKINVDCx5p33_ASAP7_75t_R g1308 ( .A(n_23), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_24), .A2(n_159), .B1(n_1038), .B2(n_1044), .Y(n_1043) );
INVxp67_ASAP7_75t_SL g1083 ( .A(n_24), .Y(n_1083) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_25), .A2(n_271), .B1(n_575), .B2(n_578), .Y(n_574) );
INVx1_ASAP7_75t_L g614 ( .A(n_25), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_26), .Y(n_1388) );
AOI22xp5_ASAP7_75t_L g1499 ( .A1(n_27), .A2(n_194), .B1(n_1468), .B2(n_1473), .Y(n_1499) );
INVx1_ASAP7_75t_L g1252 ( .A(n_28), .Y(n_1252) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_28), .A2(n_126), .B1(n_1274), .B2(n_1276), .C(n_1277), .Y(n_1273) );
INVx1_ASAP7_75t_L g1713 ( .A(n_29), .Y(n_1713) );
AOI221x1_ASAP7_75t_SL g1718 ( .A1(n_29), .A2(n_174), .B1(n_413), .B2(n_604), .C(n_1719), .Y(n_1718) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_30), .Y(n_338) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_30), .B(n_336), .Y(n_1469) );
AOI22xp33_ASAP7_75t_L g1589 ( .A1(n_31), .A2(n_165), .B1(n_1476), .B2(n_1590), .Y(n_1589) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_32), .A2(n_210), .B1(n_1020), .B2(n_1047), .Y(n_1113) );
AOI22xp5_ASAP7_75t_L g1139 ( .A1(n_32), .A2(n_277), .B1(n_678), .B2(n_820), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1508 ( .A1(n_33), .A2(n_176), .B1(n_1476), .B2(n_1478), .Y(n_1508) );
INVx1_ASAP7_75t_L g1708 ( .A(n_34), .Y(n_1708) );
AOI22xp33_ASAP7_75t_L g1725 ( .A1(n_34), .A2(n_160), .B1(n_370), .B2(n_422), .Y(n_1725) );
INVx1_ASAP7_75t_L g1335 ( .A(n_35), .Y(n_1335) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_35), .A2(n_54), .B1(n_1259), .B2(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1263 ( .A(n_36), .Y(n_1263) );
OAI22xp33_ASAP7_75t_L g1271 ( .A1(n_36), .A2(n_45), .B1(n_545), .B2(n_547), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_37), .A2(n_230), .B1(n_520), .B2(n_942), .Y(n_1206) );
AOI221xp5_ASAP7_75t_L g1216 ( .A1(n_37), .A2(n_260), .B1(n_645), .B2(n_647), .C(n_795), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_38), .A2(n_805), .B1(n_806), .B2(n_807), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_38), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g1706 ( .A(n_39), .Y(n_1706) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_40), .A2(n_256), .B1(n_1012), .B2(n_1038), .Y(n_1037) );
INVxp67_ASAP7_75t_SL g1073 ( .A(n_40), .Y(n_1073) );
INVxp67_ASAP7_75t_SL g1162 ( .A(n_41), .Y(n_1162) );
AOI22xp33_ASAP7_75t_SL g1193 ( .A1(n_41), .A2(n_74), .B1(n_515), .B2(n_1040), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g1295 ( .A1(n_42), .A2(n_557), .B1(n_1296), .B2(n_1299), .Y(n_1295) );
INVx1_ASAP7_75t_L g1314 ( .A(n_42), .Y(n_1314) );
CKINVDCx5p33_ASAP7_75t_R g1199 ( .A(n_43), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_44), .A2(n_171), .B1(n_604), .B2(n_677), .Y(n_833) );
INVx1_ASAP7_75t_L g865 ( .A(n_44), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g1256 ( .A1(n_45), .A2(n_286), .B1(n_618), .B2(n_1257), .C(n_1259), .Y(n_1256) );
AOI22xp5_ASAP7_75t_L g1484 ( .A1(n_46), .A2(n_145), .B1(n_1476), .B2(n_1478), .Y(n_1484) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_47), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g1353 ( .A1(n_48), .A2(n_308), .B1(n_703), .B2(n_707), .C(n_1354), .Y(n_1353) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_48), .A2(n_155), .B1(n_688), .B2(n_980), .Y(n_1360) );
INVx1_ASAP7_75t_L g1210 ( .A(n_49), .Y(n_1210) );
INVx1_ASAP7_75t_L g890 ( .A(n_50), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_50), .A2(n_166), .B1(n_624), .B2(n_674), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g1332 ( .A1(n_51), .A2(n_175), .B1(n_553), .B2(n_557), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g1365 ( .A(n_51), .Y(n_1365) );
CKINVDCx5p33_ASAP7_75t_R g1246 ( .A(n_52), .Y(n_1246) );
INVx1_ASAP7_75t_L g1302 ( .A(n_53), .Y(n_1302) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_53), .A2(n_56), .B1(n_408), .B2(n_677), .Y(n_1323) );
INVx1_ASAP7_75t_L g1357 ( .A(n_54), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_55), .A2(n_201), .B1(n_676), .B2(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g859 ( .A(n_55), .Y(n_859) );
AOI221xp5_ASAP7_75t_L g1290 ( .A1(n_56), .A2(n_315), .B1(n_701), .B2(n_1048), .C(n_1291), .Y(n_1290) );
OAI222xp33_ASAP7_75t_L g363 ( .A1(n_57), .A2(n_68), .B1(n_364), .B2(n_372), .C1(n_386), .C2(n_399), .Y(n_363) );
INVx1_ASAP7_75t_L g488 ( .A(n_57), .Y(n_488) );
INVxp67_ASAP7_75t_SL g1261 ( .A(n_58), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g1278 ( .A1(n_58), .A2(n_557), .B1(n_1279), .B2(n_1280), .Y(n_1278) );
AOI22xp33_ASAP7_75t_SL g1411 ( .A1(n_59), .A2(n_131), .B1(n_427), .B2(n_921), .Y(n_1411) );
AOI21xp33_ASAP7_75t_L g580 ( .A1(n_60), .A2(n_581), .B(n_584), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_60), .A2(n_91), .B1(n_644), .B2(n_646), .C(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g1094 ( .A(n_61), .Y(n_1094) );
INVx1_ASAP7_75t_L g1336 ( .A(n_62), .Y(n_1336) );
OAI21xp33_ASAP7_75t_L g1379 ( .A1(n_62), .A2(n_617), .B(n_618), .Y(n_1379) );
CKINVDCx5p33_ASAP7_75t_R g1103 ( .A(n_63), .Y(n_1103) );
INVx1_ASAP7_75t_L g1265 ( .A(n_64), .Y(n_1265) );
OAI222xp33_ASAP7_75t_L g1268 ( .A1(n_64), .A2(n_275), .B1(n_286), .B2(n_556), .C1(n_1269), .C2(n_1270), .Y(n_1268) );
XOR2x2_ASAP7_75t_L g538 ( .A(n_65), .B(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_66), .A2(n_298), .B1(n_763), .B2(n_764), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_66), .A2(n_312), .B1(n_624), .B2(n_781), .C(n_783), .Y(n_780) );
INVx1_ASAP7_75t_L g668 ( .A(n_67), .Y(n_668) );
INVx1_ASAP7_75t_L g497 ( .A(n_68), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g810 ( .A1(n_69), .A2(n_108), .B1(n_791), .B2(n_811), .C(n_814), .Y(n_810) );
INVx1_ASAP7_75t_L g841 ( .A(n_69), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g1341 ( .A(n_70), .Y(n_1341) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_71), .A2(n_326), .B1(n_515), .B2(n_938), .Y(n_945) );
AOI221xp5_ASAP7_75t_L g952 ( .A1(n_71), .A2(n_182), .B1(n_413), .B2(n_832), .C(n_953), .Y(n_952) );
CKINVDCx5p33_ASAP7_75t_R g1178 ( .A(n_72), .Y(n_1178) );
XOR2xp5_ASAP7_75t_L g1195 ( .A(n_73), .B(n_1196), .Y(n_1195) );
AOI221xp5_ASAP7_75t_L g1167 ( .A1(n_74), .A2(n_102), .B1(n_419), .B2(n_624), .C(n_1168), .Y(n_1167) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_75), .A2(n_183), .B1(n_441), .B2(n_507), .Y(n_1003) );
INVx1_ASAP7_75t_L g816 ( .A(n_77), .Y(n_816) );
OAI221xp5_ASAP7_75t_SL g848 ( .A1(n_77), .A2(n_104), .B1(n_491), .B2(n_500), .C(n_754), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_78), .A2(n_258), .B1(n_516), .B2(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g986 ( .A(n_79), .Y(n_986) );
AOI221xp5_ASAP7_75t_L g1436 ( .A1(n_80), .A2(n_302), .B1(n_1276), .B2(n_1346), .C(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1459 ( .A(n_80), .Y(n_1459) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_81), .A2(n_191), .B1(n_553), .B2(n_557), .Y(n_552) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_81), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g1467 ( .A1(n_82), .A2(n_193), .B1(n_1468), .B2(n_1473), .Y(n_1467) );
INVx1_ASAP7_75t_L g1224 ( .A(n_83), .Y(n_1224) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_84), .A2(n_98), .B1(n_703), .B2(n_707), .C(n_1047), .Y(n_1046) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_84), .A2(n_256), .B1(n_677), .B2(n_678), .Y(n_1084) );
AOI222xp33_ASAP7_75t_L g585 ( .A1(n_85), .A2(n_136), .B1(n_311), .B2(n_471), .C1(n_524), .C2(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g650 ( .A(n_85), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g1248 ( .A(n_86), .Y(n_1248) );
OAI22xp33_ASAP7_75t_L g1309 ( .A1(n_87), .A2(n_133), .B1(n_545), .B2(n_547), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_87), .A2(n_273), .B1(n_1257), .B2(n_1259), .Y(n_1324) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_88), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_88), .A2(n_263), .B1(n_515), .B2(n_516), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g1253 ( .A(n_89), .Y(n_1253) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_90), .A2(n_217), .B1(n_535), .B2(n_734), .C(n_736), .Y(n_733) );
OAI211xp5_ASAP7_75t_L g774 ( .A1(n_90), .A2(n_775), .B(n_776), .C(n_784), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g560 ( .A1(n_91), .A2(n_208), .B1(n_561), .B2(n_564), .C(n_567), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_92), .A2(n_262), .B1(n_1018), .B2(n_1020), .Y(n_1017) );
INVx1_ASAP7_75t_L g336 ( .A(n_93), .Y(n_336) );
INVx1_ASAP7_75t_L g1298 ( .A(n_94), .Y(n_1298) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_94), .A2(n_315), .B1(n_604), .B2(n_677), .Y(n_1319) );
INVx1_ASAP7_75t_L g1262 ( .A(n_95), .Y(n_1262) );
INVx1_ASAP7_75t_L g543 ( .A(n_96), .Y(n_543) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_96), .A2(n_600), .B(n_606), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_97), .A2(n_137), .B1(n_413), .B2(n_419), .C(n_832), .Y(n_834) );
INVx1_ASAP7_75t_L g853 ( .A(n_97), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g1070 ( .A1(n_98), .A2(n_143), .B1(n_832), .B2(n_1071), .C(n_1072), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_99), .A2(n_247), .B1(n_441), .B2(n_507), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g1202 ( .A1(n_100), .A2(n_235), .B1(n_1203), .B2(n_1204), .Y(n_1202) );
INVx1_ASAP7_75t_L g900 ( .A(n_101), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_101), .A2(n_146), .B1(n_604), .B2(n_677), .Y(n_916) );
XOR2x2_ASAP7_75t_L g1420 ( .A(n_103), .B(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g827 ( .A(n_104), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_105), .Y(n_887) );
INVx1_ASAP7_75t_L g436 ( .A(n_106), .Y(n_436) );
INVx1_ASAP7_75t_L g1689 ( .A(n_107), .Y(n_1689) );
OAI22xp5_ASAP7_75t_L g1726 ( .A1(n_107), .A2(n_234), .B1(n_1257), .B2(n_1259), .Y(n_1726) );
INVx1_ASAP7_75t_L g839 ( .A(n_108), .Y(n_839) );
INVx1_ASAP7_75t_L g1434 ( .A(n_109), .Y(n_1434) );
INVx1_ASAP7_75t_L g1439 ( .A(n_110), .Y(n_1439) );
XOR2x2_ASAP7_75t_L g924 ( .A(n_111), .B(n_925), .Y(n_924) );
OAI221xp5_ASAP7_75t_L g880 ( .A1(n_112), .A2(n_270), .B1(n_553), .B2(n_557), .C(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g922 ( .A(n_112), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g1090 ( .A1(n_113), .A2(n_1091), .B1(n_1092), .B2(n_1146), .Y(n_1090) );
INVx1_ASAP7_75t_L g1146 ( .A(n_113), .Y(n_1146) );
AOI22xp5_ASAP7_75t_L g1488 ( .A1(n_113), .A2(n_295), .B1(n_1468), .B2(n_1473), .Y(n_1488) );
INVx1_ASAP7_75t_L g1438 ( .A(n_114), .Y(n_1438) );
INVx1_ASAP7_75t_L g822 ( .A(n_115), .Y(n_822) );
OAI21xp33_ASAP7_75t_L g846 ( .A1(n_115), .A2(n_477), .B(n_847), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_116), .Y(n_1389) );
CKINVDCx5p33_ASAP7_75t_R g1293 ( .A(n_117), .Y(n_1293) );
OAI22xp5_ASAP7_75t_L g1435 ( .A1(n_118), .A2(n_179), .B1(n_575), .B2(n_578), .Y(n_1435) );
OAI22xp5_ASAP7_75t_L g1448 ( .A1(n_118), .A2(n_266), .B1(n_442), .B2(n_609), .Y(n_1448) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_119), .A2(n_239), .B1(n_676), .B2(n_678), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_119), .A2(n_310), .B1(n_515), .B2(n_703), .C(n_707), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g1498 ( .A1(n_120), .A2(n_197), .B1(n_1476), .B2(n_1478), .Y(n_1498) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_121), .Y(n_927) );
OAI211xp5_ASAP7_75t_SL g1165 ( .A1(n_122), .A2(n_406), .B(n_1166), .C(n_1170), .Y(n_1165) );
INVx1_ASAP7_75t_L g1187 ( .A(n_122), .Y(n_1187) );
AOI22xp33_ASAP7_75t_SL g1395 ( .A1(n_123), .A2(n_281), .B1(n_534), .B2(n_1396), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g1415 ( .A1(n_123), .A2(n_272), .B1(n_427), .B2(n_921), .Y(n_1415) );
OAI22xp5_ASAP7_75t_L g1426 ( .A1(n_124), .A2(n_203), .B1(n_553), .B2(n_557), .Y(n_1426) );
INVxp67_ASAP7_75t_SL g1446 ( .A(n_124), .Y(n_1446) );
OAI222xp33_ASAP7_75t_L g1153 ( .A1(n_125), .A2(n_252), .B1(n_962), .B2(n_1154), .C1(n_1155), .C2(n_1159), .Y(n_1153) );
INVx1_ASAP7_75t_L g1181 ( .A(n_125), .Y(n_1181) );
INVx1_ASAP7_75t_L g1236 ( .A(n_126), .Y(n_1236) );
INVx1_ASAP7_75t_L g752 ( .A(n_127), .Y(n_752) );
INVx1_ASAP7_75t_L g382 ( .A(n_128), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_128), .A2(n_186), .B1(n_520), .B2(n_523), .Y(n_519) );
XNOR2x1_ASAP7_75t_L g1149 ( .A(n_129), .B(n_1150), .Y(n_1149) );
AOI22xp5_ASAP7_75t_L g1503 ( .A1(n_129), .A2(n_209), .B1(n_1468), .B2(n_1473), .Y(n_1503) );
INVx1_ASAP7_75t_L g934 ( .A(n_130), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_131), .A2(n_294), .B1(n_471), .B2(n_523), .Y(n_1399) );
INVx1_ASAP7_75t_L g1061 ( .A(n_132), .Y(n_1061) );
INVx1_ASAP7_75t_L g1315 ( .A(n_133), .Y(n_1315) );
AOI221xp5_ASAP7_75t_SL g831 ( .A1(n_134), .A2(n_291), .B1(n_413), .B2(n_795), .C(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g862 ( .A(n_134), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_135), .Y(n_829) );
INVx1_ASAP7_75t_L g628 ( .A(n_136), .Y(n_628) );
INVx1_ASAP7_75t_L g866 ( .A(n_137), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_138), .A2(n_284), .B1(n_520), .B2(n_940), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_138), .A2(n_248), .B1(n_955), .B2(n_956), .Y(n_954) );
INVx1_ASAP7_75t_L g1343 ( .A(n_139), .Y(n_1343) );
AOI22xp33_ASAP7_75t_SL g1361 ( .A1(n_139), .A2(n_150), .B1(n_1362), .B2(n_1363), .Y(n_1361) );
INVxp67_ASAP7_75t_SL g739 ( .A(n_140), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g794 ( .A1(n_140), .A2(n_238), .B1(n_647), .B2(n_781), .C(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g883 ( .A(n_141), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_141), .A2(n_305), .B1(n_442), .B2(n_609), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g1700 ( .A(n_142), .Y(n_1700) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_143), .A2(n_167), .B1(n_704), .B2(n_1040), .C(n_1041), .Y(n_1039) );
INVxp67_ASAP7_75t_SL g1098 ( .A(n_144), .Y(n_1098) );
OAI221xp5_ASAP7_75t_L g1114 ( .A1(n_144), .A2(n_549), .B1(n_553), .B2(n_1115), .C(n_1122), .Y(n_1114) );
INVx1_ASAP7_75t_L g893 ( .A(n_146), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g1112 ( .A1(n_147), .A2(n_704), .B(n_1018), .Y(n_1112) );
INVx1_ASAP7_75t_L g1132 ( .A(n_147), .Y(n_1132) );
INVx1_ASAP7_75t_L g1121 ( .A(n_148), .Y(n_1121) );
AOI22xp33_ASAP7_75t_SL g1134 ( .A1(n_148), .A2(n_210), .B1(n_836), .B2(n_955), .Y(n_1134) );
INVx1_ASAP7_75t_L g1352 ( .A(n_150), .Y(n_1352) );
INVx1_ASAP7_75t_L g1198 ( .A(n_151), .Y(n_1198) );
OAI221xp5_ASAP7_75t_L g1425 ( .A1(n_152), .A2(n_266), .B1(n_545), .B2(n_547), .C(n_549), .Y(n_1425) );
INVxp67_ASAP7_75t_SL g1444 ( .A(n_152), .Y(n_1444) );
INVx1_ASAP7_75t_L g771 ( .A(n_153), .Y(n_771) );
INVx1_ASAP7_75t_L g1304 ( .A(n_154), .Y(n_1304) );
AOI221xp5_ASAP7_75t_L g1344 ( .A1(n_155), .A2(n_283), .B1(n_704), .B2(n_1345), .C(n_1346), .Y(n_1344) );
OAI221xp5_ASAP7_75t_L g1055 ( .A1(n_156), .A2(n_158), .B1(n_760), .B2(n_1056), .C(n_1058), .Y(n_1055) );
INVx1_ASAP7_75t_L g1171 ( .A(n_157), .Y(n_1171) );
INVxp67_ASAP7_75t_SL g1067 ( .A(n_158), .Y(n_1067) );
INVxp33_ASAP7_75t_SL g1074 ( .A(n_159), .Y(n_1074) );
INVx1_ASAP7_75t_L g1702 ( .A(n_160), .Y(n_1702) );
INVx2_ASAP7_75t_L g1471 ( .A(n_161), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_161), .B(n_1472), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_161), .B(n_278), .Y(n_1479) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_162), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_162), .A2(n_296), .B1(n_533), .B2(n_534), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g1483 ( .A1(n_163), .A2(n_257), .B1(n_1468), .B2(n_1473), .Y(n_1483) );
INVx1_ASAP7_75t_L g1211 ( .A(n_164), .Y(n_1211) );
INVx1_ASAP7_75t_L g898 ( .A(n_166), .Y(n_898) );
INVx1_ASAP7_75t_L g1081 ( .A(n_167), .Y(n_1081) );
INVx1_ASAP7_75t_L g923 ( .A(n_168), .Y(n_923) );
OAI21xp33_ASAP7_75t_L g663 ( .A1(n_169), .A2(n_664), .B(n_666), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_169), .A2(n_268), .B1(n_715), .B2(n_716), .C(n_718), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g1489 ( .A1(n_170), .A2(n_288), .B1(n_1476), .B2(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g852 ( .A(n_171), .Y(n_852) );
OAI21xp5_ASAP7_75t_SL g1330 ( .A1(n_172), .A2(n_878), .B(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1356 ( .A(n_172), .Y(n_1356) );
CKINVDCx5p33_ASAP7_75t_R g1697 ( .A(n_173), .Y(n_1697) );
INVx1_ASAP7_75t_L g1704 ( .A(n_174), .Y(n_1704) );
INVx1_ASAP7_75t_L g1373 ( .A(n_175), .Y(n_1373) );
INVxp67_ASAP7_75t_SL g997 ( .A(n_177), .Y(n_997) );
CKINVDCx5p33_ASAP7_75t_R g1393 ( .A(n_178), .Y(n_1393) );
OAI211xp5_ASAP7_75t_L g1441 ( .A1(n_179), .A2(n_878), .B(n_1442), .C(n_1445), .Y(n_1441) );
INVx1_ASAP7_75t_L g1060 ( .A(n_181), .Y(n_1060) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_181), .A2(n_223), .B1(n_442), .B2(n_609), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_182), .A2(n_192), .B1(n_515), .B2(n_938), .Y(n_937) );
OAI211xp5_ASAP7_75t_L g977 ( .A1(n_183), .A2(n_406), .B(n_978), .C(n_985), .Y(n_977) );
CKINVDCx5p33_ASAP7_75t_R g1124 ( .A(n_184), .Y(n_1124) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_185), .A2(n_300), .B1(n_415), .B2(n_674), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_185), .A2(n_218), .B1(n_520), .B2(n_703), .C(n_704), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_186), .A2(n_327), .B1(n_422), .B2(n_426), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_187), .A2(n_235), .B1(n_676), .B2(n_678), .Y(n_1217) );
AOI22xp33_ASAP7_75t_SL g1400 ( .A1(n_188), .A2(n_272), .B1(n_462), .B2(n_534), .Y(n_1400) );
AOI221xp5_ASAP7_75t_L g1407 ( .A1(n_188), .A2(n_281), .B1(n_646), .B2(n_783), .C(n_1408), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_189), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g496 ( .A(n_189), .Y(n_496) );
INVx1_ASAP7_75t_L g531 ( .A(n_189), .Y(n_531) );
OAI211xp5_ASAP7_75t_L g1333 ( .A1(n_190), .A2(n_549), .B(n_720), .C(n_1334), .Y(n_1333) );
CKINVDCx5p33_ASAP7_75t_R g1378 ( .A(n_190), .Y(n_1378) );
INVxp67_ASAP7_75t_SL g591 ( .A(n_191), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_192), .A2(n_326), .B1(n_676), .B2(n_956), .Y(n_968) );
XOR2xp5_ASAP7_75t_L g1681 ( .A(n_193), .B(n_1682), .Y(n_1681) );
AOI22xp5_ASAP7_75t_L g1734 ( .A1(n_193), .A2(n_1735), .B1(n_1740), .B2(n_1745), .Y(n_1734) );
INVx1_ASAP7_75t_L g1229 ( .A(n_195), .Y(n_1229) );
OAI221xp5_ASAP7_75t_SL g991 ( .A1(n_196), .A2(n_279), .B1(n_364), .B2(n_961), .C(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g1007 ( .A(n_196), .Y(n_1007) );
INVx1_ASAP7_75t_L g903 ( .A(n_198), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_198), .A2(n_301), .B1(n_427), .B2(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g1493 ( .A1(n_199), .A2(n_289), .B1(n_1468), .B2(n_1473), .Y(n_1493) );
OAI22xp33_ASAP7_75t_L g1690 ( .A1(n_200), .A2(n_290), .B1(n_751), .B2(n_1042), .Y(n_1690) );
INVx1_ASAP7_75t_L g1730 ( .A(n_200), .Y(n_1730) );
INVx1_ASAP7_75t_L g863 ( .A(n_201), .Y(n_863) );
CKINVDCx5p33_ASAP7_75t_R g1404 ( .A(n_202), .Y(n_1404) );
INVxp67_ASAP7_75t_SL g1443 ( .A(n_203), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_204), .A2(n_309), .B1(n_676), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_204), .A2(n_239), .B1(n_515), .B2(n_701), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_205), .A2(n_282), .B1(n_929), .B2(n_930), .Y(n_928) );
OAI211xp5_ASAP7_75t_L g949 ( .A1(n_205), .A2(n_950), .B(n_951), .C(n_957), .Y(n_949) );
INVx1_ASAP7_75t_L g377 ( .A(n_206), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g525 ( .A1(n_206), .A2(n_327), .B1(n_523), .B2(n_526), .Y(n_525) );
BUFx3_ASAP7_75t_L g455 ( .A(n_207), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_208), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g569 ( .A(n_211), .Y(n_569) );
OAI21xp5_ASAP7_75t_SL g1418 ( .A1(n_212), .A2(n_441), .B(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g667 ( .A(n_213), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g1305 ( .A1(n_214), .A2(n_273), .B1(n_1110), .B2(n_1306), .C(n_1307), .Y(n_1305) );
OAI211xp5_ASAP7_75t_L g1312 ( .A1(n_214), .A2(n_722), .B(n_1313), .C(n_1316), .Y(n_1312) );
OAI21xp5_ASAP7_75t_SL g440 ( .A1(n_215), .A2(n_441), .B(n_460), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g1292 ( .A(n_216), .Y(n_1292) );
OAI221xp5_ASAP7_75t_SL g785 ( .A1(n_217), .A2(n_304), .B1(n_399), .B2(n_786), .C(n_788), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_218), .A2(n_310), .B1(n_688), .B2(n_689), .Y(n_687) );
OAI21xp5_ASAP7_75t_L g1173 ( .A1(n_219), .A2(n_929), .B(n_1174), .Y(n_1173) );
XOR2xp5_ASAP7_75t_L g974 ( .A(n_220), .B(n_975), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_221), .A2(n_262), .B1(n_685), .B2(n_984), .Y(n_983) );
OAI22xp33_ASAP7_75t_L g946 ( .A1(n_222), .A2(n_322), .B1(n_766), .B2(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g958 ( .A(n_222), .Y(n_958) );
INVx1_ASAP7_75t_L g1050 ( .A(n_223), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_224), .Y(n_1002) );
CKINVDCx5p33_ASAP7_75t_R g1097 ( .A(n_225), .Y(n_1097) );
INVx1_ASAP7_75t_L g1432 ( .A(n_226), .Y(n_1432) );
AOI22xp5_ASAP7_75t_L g1475 ( .A1(n_227), .A2(n_246), .B1(n_1476), .B2(n_1478), .Y(n_1475) );
CKINVDCx5p33_ASAP7_75t_R g1242 ( .A(n_228), .Y(n_1242) );
INVx1_ASAP7_75t_L g432 ( .A(n_229), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_231), .A2(n_248), .B1(n_520), .B2(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g964 ( .A(n_231), .Y(n_964) );
OAI211xp5_ASAP7_75t_L g884 ( .A1(n_232), .A2(n_508), .B(n_549), .C(n_885), .Y(n_884) );
INVxp33_ASAP7_75t_SL g911 ( .A(n_232), .Y(n_911) );
INVx1_ASAP7_75t_L g1424 ( .A(n_233), .Y(n_1424) );
OAI221xp5_ASAP7_75t_L g1693 ( .A1(n_234), .A2(n_251), .B1(n_491), .B2(n_500), .C(n_854), .Y(n_1693) );
BUFx3_ASAP7_75t_L g353 ( .A(n_236), .Y(n_353) );
INVx1_ASAP7_75t_L g369 ( .A(n_236), .Y(n_369) );
OAI211xp5_ASAP7_75t_L g405 ( .A1(n_237), .A2(n_406), .B(n_410), .C(n_429), .Y(n_405) );
INVx1_ASAP7_75t_L g505 ( .A(n_237), .Y(n_505) );
INVx1_ASAP7_75t_L g757 ( .A(n_238), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g1142 ( .A(n_240), .B(n_1143), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g1710 ( .A(n_241), .Y(n_1710) );
OAI322xp33_ASAP7_75t_SL g737 ( .A1(n_242), .A2(n_738), .A3(n_745), .B1(n_748), .B2(n_756), .C1(n_765), .C2(n_766), .Y(n_737) );
OAI22xp33_ASAP7_75t_SL g796 ( .A1(n_242), .A2(n_247), .B1(n_406), .B2(n_797), .Y(n_796) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_243), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_244), .Y(n_815) );
INVx1_ASAP7_75t_L g1105 ( .A(n_245), .Y(n_1105) );
CKINVDCx5p33_ASAP7_75t_R g1300 ( .A(n_249), .Y(n_1300) );
INVx1_ASAP7_75t_L g761 ( .A(n_250), .Y(n_761) );
OA222x2_ASAP7_75t_L g1727 ( .A1(n_251), .A2(n_265), .B1(n_313), .B2(n_600), .C1(n_617), .C2(n_664), .Y(n_1727) );
INVx1_ASAP7_75t_L g1184 ( .A(n_252), .Y(n_1184) );
OAI21xp5_ASAP7_75t_L g1225 ( .A1(n_253), .A2(n_441), .B(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g572 ( .A(n_254), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g1118 ( .A(n_255), .Y(n_1118) );
XOR2x2_ASAP7_75t_L g360 ( .A(n_257), .B(n_361), .Y(n_360) );
INVxp67_ASAP7_75t_SL g995 ( .A(n_258), .Y(n_995) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_259), .A2(n_727), .B1(n_728), .B2(n_801), .Y(n_726) );
INVx1_ASAP7_75t_L g801 ( .A(n_259), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_259), .A2(n_727), .B1(n_728), .B2(n_801), .Y(n_868) );
AOI211xp5_ASAP7_75t_L g1428 ( .A1(n_261), .A2(n_703), .B(n_1429), .C(n_1431), .Y(n_1428) );
INVx1_ASAP7_75t_L g1456 ( .A(n_261), .Y(n_1456) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_263), .A2(n_296), .B1(n_412), .B2(n_413), .C(n_419), .Y(n_411) );
INVx1_ASAP7_75t_L g453 ( .A(n_264), .Y(n_453) );
INVx1_ASAP7_75t_L g468 ( .A(n_264), .Y(n_468) );
INVx1_ASAP7_75t_L g1692 ( .A(n_265), .Y(n_1692) );
INVx1_ASAP7_75t_L g682 ( .A(n_267), .Y(n_682) );
INVxp67_ASAP7_75t_SL g723 ( .A(n_268), .Y(n_723) );
CKINVDCx5p33_ASAP7_75t_R g1240 ( .A(n_269), .Y(n_1240) );
INVxp67_ASAP7_75t_SL g909 ( .A(n_270), .Y(n_909) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_271), .Y(n_597) );
INVx1_ASAP7_75t_L g1059 ( .A(n_274), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g1062 ( .A(n_274), .B(n_878), .Y(n_1062) );
INVx1_ASAP7_75t_L g1283 ( .A(n_275), .Y(n_1283) );
CKINVDCx5p33_ASAP7_75t_R g1405 ( .A(n_276), .Y(n_1405) );
INVx1_ASAP7_75t_L g1125 ( .A(n_277), .Y(n_1125) );
INVx1_ASAP7_75t_L g1472 ( .A(n_278), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_278), .B(n_1471), .Y(n_1477) );
INVx1_ASAP7_75t_L g1008 ( .A(n_279), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_280), .Y(n_485) );
AOI221xp5_ASAP7_75t_SL g1366 ( .A1(n_283), .A2(n_285), .B1(n_980), .B2(n_1367), .C(n_1368), .Y(n_1366) );
AOI21xp33_ASAP7_75t_L g967 ( .A1(n_284), .A2(n_413), .B(n_795), .Y(n_967) );
INVx1_ASAP7_75t_L g1351 ( .A(n_285), .Y(n_1351) );
OAI22xp5_ASAP7_75t_L g1327 ( .A1(n_287), .A2(n_1328), .B1(n_1329), .B2(n_1382), .Y(n_1327) );
INVx1_ASAP7_75t_L g1382 ( .A(n_287), .Y(n_1382) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_287), .A2(n_319), .B1(n_1468), .B2(n_1473), .Y(n_1509) );
INVx1_ASAP7_75t_L g1729 ( .A(n_290), .Y(n_1729) );
INVx1_ASAP7_75t_L g856 ( .A(n_291), .Y(n_856) );
INVx1_ASAP7_75t_L g1157 ( .A(n_292), .Y(n_1157) );
INVx1_ASAP7_75t_L g1430 ( .A(n_293), .Y(n_1430) );
INVx1_ASAP7_75t_L g1223 ( .A(n_297), .Y(n_1223) );
INVxp67_ASAP7_75t_SL g793 ( .A(n_298), .Y(n_793) );
INVx1_ASAP7_75t_L g1106 ( .A(n_299), .Y(n_1106) );
OAI221xp5_ASAP7_75t_L g1135 ( .A1(n_299), .A2(n_617), .B1(n_1136), .B2(n_1140), .C(n_1141), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_300), .A2(n_309), .B1(n_701), .B2(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g895 ( .A(n_301), .Y(n_895) );
INVx1_ASAP7_75t_L g1452 ( .A(n_302), .Y(n_1452) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_304), .Y(n_730) );
INVx1_ASAP7_75t_L g886 ( .A(n_305), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g1392 ( .A(n_306), .Y(n_1392) );
CKINVDCx5p33_ASAP7_75t_R g1297 ( .A(n_307), .Y(n_1297) );
INVx1_ASAP7_75t_L g1369 ( .A(n_308), .Y(n_1369) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_311), .A2(n_412), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g755 ( .A(n_312), .Y(n_755) );
INVx1_ASAP7_75t_L g1687 ( .A(n_313), .Y(n_1687) );
CKINVDCx5p33_ASAP7_75t_R g1237 ( .A(n_314), .Y(n_1237) );
INVx1_ASAP7_75t_L g1088 ( .A(n_317), .Y(n_1088) );
XOR2xp5_ASAP7_75t_L g1385 ( .A(n_318), .B(n_1386), .Y(n_1385) );
INVx2_ASAP7_75t_L g439 ( .A(n_320), .Y(n_439) );
INVx1_ASAP7_75t_L g448 ( .A(n_320), .Y(n_448) );
INVx1_ASAP7_75t_L g483 ( .A(n_320), .Y(n_483) );
INVx1_ASAP7_75t_L g607 ( .A(n_321), .Y(n_607) );
INVx1_ASAP7_75t_L g959 ( .A(n_322), .Y(n_959) );
INVx1_ASAP7_75t_L g1286 ( .A(n_323), .Y(n_1286) );
CKINVDCx5p33_ASAP7_75t_R g1108 ( .A(n_324), .Y(n_1108) );
OAI21xp33_ASAP7_75t_SL g877 ( .A1(n_325), .A2(n_878), .B(n_879), .Y(n_877) );
INVx1_ASAP7_75t_L g882 ( .A(n_325), .Y(n_882) );
INVx1_ASAP7_75t_L g742 ( .A(n_328), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_354), .B(n_1461), .Y(n_329) );
BUFx4f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_339), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g1733 ( .A(n_333), .B(n_342), .Y(n_1733) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g1739 ( .A(n_335), .B(n_338), .Y(n_1739) );
INVx1_ASAP7_75t_L g1749 ( .A(n_335), .Y(n_1749) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g1751 ( .A(n_338), .B(n_1749), .Y(n_1751) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g385 ( .A(n_343), .B(n_352), .Y(n_385) );
AND2x4_ASAP7_75t_L g420 ( .A(n_343), .B(n_353), .Y(n_420) );
AND2x4_ASAP7_75t_SL g1732 ( .A(n_344), .B(n_1733), .Y(n_1732) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_346), .B(n_351), .Y(n_345) );
BUFx4f_ASAP7_75t_L g627 ( .A(n_346), .Y(n_627) );
INVxp67_ASAP7_75t_L g1251 ( .A(n_346), .Y(n_1251) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx3_ASAP7_75t_L g390 ( .A(n_347), .Y(n_390) );
BUFx4f_ASAP7_75t_L g792 ( .A(n_347), .Y(n_792) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x2_ASAP7_75t_L g371 ( .A(n_349), .B(n_350), .Y(n_371) );
NAND2x1_ASAP7_75t_L g376 ( .A(n_349), .B(n_350), .Y(n_376) );
INVx2_ASAP7_75t_L g381 ( .A(n_349), .Y(n_381) );
INVx2_ASAP7_75t_L g397 ( .A(n_349), .Y(n_397) );
AND2x2_ASAP7_75t_L g417 ( .A(n_349), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g445 ( .A(n_349), .Y(n_445) );
OR2x2_ASAP7_75t_L g380 ( .A(n_350), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_350), .B(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_L g402 ( .A(n_350), .Y(n_402) );
AND2x2_ASAP7_75t_L g409 ( .A(n_350), .B(n_397), .Y(n_409) );
INVx2_ASAP7_75t_L g418 ( .A(n_350), .Y(n_418) );
INVx1_ASAP7_75t_L g425 ( .A(n_350), .Y(n_425) );
INVxp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
XOR2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_1027), .Y(n_354) );
XNOR2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_870), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B1(n_653), .B2(n_869), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_537), .B2(n_652), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND3x1_ASAP7_75t_L g361 ( .A(n_362), .B(n_474), .C(n_486), .Y(n_361) );
O2A1O1Ixp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_405), .B(n_437), .C(n_440), .Y(n_362) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g775 ( .A(n_365), .Y(n_775) );
INVx2_ASAP7_75t_L g1154 ( .A(n_365), .Y(n_1154) );
INVx4_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g1215 ( .A(n_367), .Y(n_1215) );
AND2x4_ASAP7_75t_SL g367 ( .A(n_368), .B(n_370), .Y(n_367) );
AND2x4_ASAP7_75t_L g407 ( .A(n_368), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g431 ( .A(n_368), .B(n_424), .Y(n_431) );
AND2x4_ASAP7_75t_L g434 ( .A(n_368), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g594 ( .A(n_368), .B(n_435), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_368), .B(n_483), .Y(n_603) );
BUFx2_ASAP7_75t_L g817 ( .A(n_368), .Y(n_817) );
BUFx3_ASAP7_75t_L g412 ( .A(n_370), .Y(n_412) );
AND2x6_ASAP7_75t_L g428 ( .A(n_370), .B(n_404), .Y(n_428) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_370), .Y(n_645) );
BUFx3_ASAP7_75t_L g674 ( .A(n_370), .Y(n_674) );
INVx1_ASAP7_75t_L g782 ( .A(n_370), .Y(n_782) );
BUFx3_ASAP7_75t_L g832 ( .A(n_370), .Y(n_832) );
BUFx3_ASAP7_75t_L g915 ( .A(n_370), .Y(n_915) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g691 ( .A(n_371), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_377), .B1(n_378), .B2(n_382), .C(n_383), .Y(n_372) );
INVx5_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g617 ( .A(n_375), .B(n_603), .Y(n_617) );
OR2x2_ASAP7_75t_L g670 ( .A(n_375), .B(n_603), .Y(n_670) );
BUFx3_ASAP7_75t_L g1247 ( .A(n_375), .Y(n_1247) );
BUFx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_376), .Y(n_619) );
OAI221xp5_ASAP7_75t_L g1321 ( .A1(n_378), .A2(n_1292), .B1(n_1297), .B2(n_1322), .C(n_1323), .Y(n_1321) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g1131 ( .A(n_379), .Y(n_1131) );
BUFx2_ASAP7_75t_L g1245 ( .A(n_379), .Y(n_1245) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g813 ( .A(n_380), .Y(n_813) );
BUFx3_ASAP7_75t_L g1080 ( .A(n_380), .Y(n_1080) );
INVx1_ASAP7_75t_L g1724 ( .A(n_380), .Y(n_1724) );
AND2x2_ASAP7_75t_L g424 ( .A(n_381), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g795 ( .A(n_385), .Y(n_795) );
INVx2_ASAP7_75t_L g999 ( .A(n_385), .Y(n_999) );
OAI221xp5_ASAP7_75t_L g1155 ( .A1(n_385), .A2(n_1078), .B1(n_1156), .B2(n_1157), .C(n_1158), .Y(n_1155) );
INVx1_ASAP7_75t_L g1414 ( .A(n_385), .Y(n_1414) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_391), .B2(n_398), .Y(n_386) );
OAI221xp5_ASAP7_75t_L g776 ( .A1(n_388), .A2(n_742), .B1(n_761), .B2(n_777), .C(n_780), .Y(n_776) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g649 ( .A(n_390), .Y(n_649) );
BUFx3_ASAP7_75t_L g1720 ( .A(n_390), .Y(n_1720) );
BUFx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_394), .Y(n_630) );
INVx2_ASAP7_75t_L g651 ( .A(n_394), .Y(n_651) );
INVx4_ASAP7_75t_L g779 ( .A(n_394), .Y(n_779) );
INVx1_ASAP7_75t_L g996 ( .A(n_394), .Y(n_996) );
INVx1_ASAP7_75t_L g1164 ( .A(n_394), .Y(n_1164) );
INVx2_ASAP7_75t_SL g1238 ( .A(n_394), .Y(n_1238) );
INVx8_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g962 ( .A(n_400), .Y(n_962) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g613 ( .A(n_402), .Y(n_613) );
BUFx2_ASAP7_75t_L g826 ( .A(n_402), .Y(n_826) );
INVx1_ASAP7_75t_L g823 ( .A(n_403), .Y(n_823) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_404), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_404), .B(n_424), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_404), .B(n_439), .Y(n_611) );
AND2x2_ASAP7_75t_L g825 ( .A(n_404), .B(n_826), .Y(n_825) );
INVx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_SL g950 ( .A(n_407), .Y(n_950) );
AOI221xp5_ASAP7_75t_L g1218 ( .A1(n_407), .A2(n_428), .B1(n_1198), .B2(n_1219), .C(n_1220), .Y(n_1218) );
AOI221xp5_ASAP7_75t_L g1406 ( .A1(n_407), .A2(n_428), .B1(n_1388), .B2(n_1407), .C(n_1411), .Y(n_1406) );
INVx1_ASAP7_75t_L g686 ( .A(n_408), .Y(n_686) );
BUFx2_ASAP7_75t_L g836 ( .A(n_408), .Y(n_836) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_408), .Y(n_956) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx3_ASAP7_75t_L g427 ( .A(n_409), .Y(n_427) );
INVx2_ASAP7_75t_L g605 ( .A(n_409), .Y(n_605) );
BUFx3_ASAP7_75t_L g678 ( .A(n_409), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_421), .B(n_428), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_412), .A2(n_427), .B1(n_815), .B2(n_816), .Y(n_814) );
A2O1A1Ixp33_ASAP7_75t_L g819 ( .A1(n_412), .A2(n_820), .B(n_822), .C(n_823), .Y(n_819) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g688 ( .A(n_414), .Y(n_688) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
HB1xp67_ASAP7_75t_L g1367 ( .A(n_415), .Y(n_1367) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g1071 ( .A(n_416), .Y(n_1071) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_417), .Y(n_435) );
BUFx3_ASAP7_75t_L g647 ( .A(n_417), .Y(n_647) );
INVx4_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g640 ( .A(n_420), .B(n_641), .Y(n_640) );
INVx4_ASAP7_75t_L g783 ( .A(n_420), .Y(n_783) );
INVx1_ASAP7_75t_SL g953 ( .A(n_420), .Y(n_953) );
AND2x2_ASAP7_75t_SL g1255 ( .A(n_420), .B(n_457), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1320 ( .A(n_420), .B(n_641), .Y(n_1320) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_SL g921 ( .A(n_423), .Y(n_921) );
INVx2_ASAP7_75t_L g955 ( .A(n_423), .Y(n_955) );
INVx1_ASAP7_75t_L g1362 ( .A(n_423), .Y(n_1362) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_424), .Y(n_677) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g1364 ( .A(n_427), .Y(n_1364) );
INVx1_ASAP7_75t_L g784 ( .A(n_428), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g951 ( .A1(n_428), .A2(n_952), .B(n_954), .Y(n_951) );
AOI21xp5_ASAP7_75t_L g978 ( .A1(n_428), .A2(n_979), .B(n_983), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g1166 ( .A1(n_428), .A2(n_1167), .B(n_1169), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B1(n_433), .B2(n_436), .Y(n_429) );
INVx1_ASAP7_75t_L g797 ( .A(n_430), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_430), .A2(n_434), .B1(n_958), .B2(n_959), .Y(n_957) );
HB1xp67_ASAP7_75t_L g987 ( .A(n_430), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_430), .A2(n_434), .B1(n_1171), .B2(n_1172), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_430), .A2(n_434), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1403 ( .A1(n_430), .A2(n_433), .B1(n_1404), .B2(n_1405), .Y(n_1403) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g598 ( .A(n_431), .B(n_593), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_432), .A2(n_436), .B1(n_461), .B2(n_470), .Y(n_460) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_434), .Y(n_787) );
INVx1_ASAP7_75t_L g990 ( .A(n_434), .Y(n_990) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_435), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_437), .A2(n_541), .B(n_559), .C(n_590), .Y(n_540) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
AND3x4_ASAP7_75t_L g512 ( .A(n_438), .B(n_496), .C(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_438), .A2(n_693), .B1(n_721), .B2(n_723), .Y(n_692) );
OAI31xp33_ASAP7_75t_SL g879 ( .A1(n_438), .A2(n_880), .A3(n_884), .B(n_888), .Y(n_879) );
INVx1_ASAP7_75t_L g972 ( .A(n_438), .Y(n_972) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g634 ( .A(n_439), .Y(n_634) );
AND2x4_ASAP7_75t_L g441 ( .A(n_442), .B(n_449), .Y(n_441) );
INVx2_ASAP7_75t_SL g615 ( .A(n_442), .Y(n_615) );
AND2x4_ASAP7_75t_L g929 ( .A(n_442), .B(n_449), .Y(n_929) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g828 ( .A(n_443), .Y(n_828) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_443), .B(n_446), .Y(n_1259) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_L g509 ( .A(n_446), .Y(n_509) );
INVx1_ASAP7_75t_L g593 ( .A(n_446), .Y(n_593) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g457 ( .A(n_447), .Y(n_457) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g844 ( .A(n_449), .Y(n_844) );
OR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_456), .Y(n_449) );
INVx4_ASAP7_75t_L g566 ( .A(n_450), .Y(n_566) );
BUFx6f_ASAP7_75t_L g854 ( .A(n_450), .Y(n_854) );
INVx3_ASAP7_75t_L g1111 ( .A(n_450), .Y(n_1111) );
OAI221xp5_ASAP7_75t_L g1291 ( .A1(n_450), .A2(n_573), .B1(n_1292), .B2(n_1293), .C(n_1294), .Y(n_1291) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g550 ( .A(n_451), .Y(n_550) );
BUFx3_ASAP7_75t_L g754 ( .A(n_451), .Y(n_754) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_453), .B(n_455), .Y(n_480) );
INVx2_ASAP7_75t_L g503 ( .A(n_453), .Y(n_503) );
INVx2_ASAP7_75t_L g491 ( .A(n_454), .Y(n_491) );
AND2x4_ASAP7_75t_L g524 ( .A(n_454), .B(n_502), .Y(n_524) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g465 ( .A(n_455), .Y(n_465) );
AND2x4_ASAP7_75t_L g518 ( .A(n_455), .B(n_503), .Y(n_518) );
OR2x2_ASAP7_75t_L g587 ( .A(n_455), .B(n_467), .Y(n_587) );
INVx1_ASAP7_75t_L g469 ( .A(n_456), .Y(n_469) );
OR2x2_ASAP7_75t_L g477 ( .A(n_456), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g769 ( .A(n_456), .Y(n_769) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g642 ( .A(n_457), .Y(n_642) );
OR2x2_ASAP7_75t_L g747 ( .A(n_457), .B(n_705), .Y(n_747) );
INVx1_ASAP7_75t_L g555 ( .A(n_458), .Y(n_555) );
INVx1_ASAP7_75t_L g577 ( .A(n_458), .Y(n_577) );
INVx3_ASAP7_75t_L g494 ( .A(n_459), .Y(n_494) );
BUFx3_ASAP7_75t_L g513 ( .A(n_459), .Y(n_513) );
NAND2xp33_ASAP7_75t_SL g705 ( .A(n_459), .B(n_496), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_461), .B(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_461), .A2(n_470), .B1(n_1404), .B2(n_1405), .Y(n_1419) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_469), .Y(n_461) );
AND2x4_ASAP7_75t_L g1175 ( .A(n_462), .B(n_469), .Y(n_1175) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx8_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
INVx3_ASAP7_75t_L g533 ( .A(n_463), .Y(n_533) );
INVx2_ASAP7_75t_L g763 ( .A(n_463), .Y(n_763) );
INVx8_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2x1p5_ASAP7_75t_L g508 ( .A(n_464), .B(n_493), .Y(n_508) );
BUFx3_ASAP7_75t_L g571 ( .A(n_464), .Y(n_571) );
AND2x2_ASAP7_75t_L g576 ( .A(n_464), .B(n_577), .Y(n_576) );
BUFx3_ASAP7_75t_L g1048 ( .A(n_464), .Y(n_1048) );
HB1xp67_ASAP7_75t_L g1203 ( .A(n_464), .Y(n_1203) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
AND2x4_ASAP7_75t_L g472 ( .A(n_465), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVxp67_ASAP7_75t_L g473 ( .A(n_468), .Y(n_473) );
AND2x4_ASAP7_75t_L g470 ( .A(n_469), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g732 ( .A(n_470), .Y(n_732) );
INVx2_ASAP7_75t_L g947 ( .A(n_470), .Y(n_947) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_471), .Y(n_526) );
INVx3_ASAP7_75t_L g710 ( .A(n_471), .Y(n_710) );
INVx3_ASAP7_75t_L g1019 ( .A(n_471), .Y(n_1019) );
INVx2_ASAP7_75t_SL g1123 ( .A(n_471), .Y(n_1123) );
BUFx8_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_472), .Y(n_522) );
INVx2_ASAP7_75t_L g556 ( .A(n_472), .Y(n_556) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_472), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_485), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_475), .A2(n_771), .B(n_772), .Y(n_770) );
AOI21xp33_ASAP7_75t_L g926 ( .A1(n_475), .A2(n_927), .B(n_928), .Y(n_926) );
AOI21xp5_ASAP7_75t_L g1001 ( .A1(n_475), .A2(n_1002), .B(n_1003), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_475), .B(n_1178), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1197 ( .A1(n_475), .A2(n_1188), .B1(n_1198), .B2(n_1199), .C(n_1200), .Y(n_1197) );
AOI221xp5_ASAP7_75t_L g1387 ( .A1(n_475), .A2(n_1188), .B1(n_1388), .B2(n_1389), .C(n_1390), .Y(n_1387) );
INVx8_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g905 ( .A(n_478), .Y(n_905) );
BUFx3_ASAP7_75t_L g1342 ( .A(n_478), .Y(n_1342) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_479), .Y(n_717) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g744 ( .A(n_480), .Y(n_744) );
INVx1_ASAP7_75t_L g665 ( .A(n_481), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_481), .B(n_1145), .Y(n_1144) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
AND2x4_ASAP7_75t_L g492 ( .A(n_482), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g638 ( .A(n_482), .Y(n_638) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g530 ( .A(n_483), .Y(n_530) );
INVx1_ASAP7_75t_L g639 ( .A(n_484), .Y(n_639) );
AND4x1_ASAP7_75t_SL g486 ( .A(n_487), .B(n_504), .C(n_510), .D(n_535), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B1(n_497), .B2(n_498), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_489), .A2(n_498), .B1(n_1007), .B2(n_1008), .Y(n_1006) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
AND2x6_ASAP7_75t_L g546 ( .A(n_490), .B(n_493), .Y(n_546) );
AND2x2_ASAP7_75t_L g735 ( .A(n_490), .B(n_492), .Y(n_735) );
NAND2x1_ASAP7_75t_L g1183 ( .A(n_490), .B(n_492), .Y(n_1183) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x4_ASAP7_75t_L g498 ( .A(n_492), .B(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g536 ( .A(n_492), .B(n_517), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g847 ( .A1(n_492), .A2(n_515), .B(n_815), .C(n_848), .Y(n_847) );
AND2x4_ASAP7_75t_SL g1185 ( .A(n_492), .B(n_499), .Y(n_1185) );
AND2x2_ASAP7_75t_L g548 ( .A(n_493), .B(n_501), .Y(n_548) );
INVx1_ASAP7_75t_L g551 ( .A(n_493), .Y(n_551) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
NAND3x1_ASAP7_75t_L g529 ( .A(n_494), .B(n_530), .C(n_531), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g589 ( .A(n_494), .B(n_531), .Y(n_589) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g573 ( .A(n_496), .B(n_513), .Y(n_573) );
INVx1_ASAP7_75t_L g736 ( .A(n_498), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_498), .A2(n_735), .B1(n_934), .B2(n_935), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_498), .A2(n_735), .B1(n_1210), .B2(n_1211), .Y(n_1209) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_498), .A2(n_1182), .B1(n_1392), .B2(n_1393), .Y(n_1391) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx5_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g1188 ( .A(n_507), .Y(n_1188) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g542 ( .A(n_508), .Y(n_542) );
OR2x2_ASAP7_75t_L g930 ( .A(n_508), .B(n_509), .Y(n_930) );
AOI33xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_514), .A3(n_519), .B1(n_525), .B2(n_527), .B3(n_532), .Y(n_510) );
AOI33xp33_ASAP7_75t_L g1009 ( .A1(n_511), .A2(n_1010), .A3(n_1013), .B1(n_1017), .B2(n_1021), .B3(n_1022), .Y(n_1009) );
AOI33xp33_ASAP7_75t_L g1394 ( .A1(n_511), .A2(n_527), .A3(n_1395), .B1(n_1398), .B2(n_1399), .B3(n_1400), .Y(n_1394) );
BUFx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI33xp33_ASAP7_75t_L g936 ( .A1(n_512), .A2(n_937), .A3(n_939), .B1(n_941), .B2(n_943), .B3(n_945), .Y(n_936) );
AOI33xp33_ASAP7_75t_L g1189 ( .A1(n_512), .A2(n_1190), .A3(n_1191), .B1(n_1192), .B2(n_1193), .B3(n_1194), .Y(n_1189) );
AOI33xp33_ASAP7_75t_L g1201 ( .A1(n_512), .A2(n_943), .A3(n_1202), .B1(n_1206), .B2(n_1207), .B3(n_1208), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_515), .A2(n_1040), .B1(n_1097), .B2(n_1103), .Y(n_1102) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_517), .A2(n_533), .B1(n_661), .B2(n_682), .Y(n_718) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g534 ( .A(n_518), .Y(n_534) );
AND2x2_ASAP7_75t_L g579 ( .A(n_518), .B(n_577), .Y(n_579) );
BUFx3_ASAP7_75t_L g703 ( .A(n_518), .Y(n_703) );
BUFx2_ASAP7_75t_L g764 ( .A(n_518), .Y(n_764) );
BUFx2_ASAP7_75t_L g938 ( .A(n_518), .Y(n_938) );
BUFx2_ASAP7_75t_L g1040 ( .A(n_518), .Y(n_1040) );
INVx2_ASAP7_75t_L g1205 ( .A(n_518), .Y(n_1205) );
INVx8_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_521), .A2(n_856), .B1(n_857), .B2(n_859), .Y(n_855) );
INVx5_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx3_ASAP7_75t_L g760 ( .A(n_522), .Y(n_760) );
INVx2_ASAP7_75t_SL g1042 ( .A(n_522), .Y(n_1042) );
INVx2_ASAP7_75t_SL g1045 ( .A(n_522), .Y(n_1045) );
HB1xp67_ASAP7_75t_L g1699 ( .A(n_522), .Y(n_1699) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g558 ( .A(n_524), .B(n_555), .Y(n_558) );
INVx5_ASAP7_75t_L g568 ( .A(n_524), .Y(n_568) );
BUFx12f_ASAP7_75t_L g701 ( .A(n_524), .Y(n_701) );
BUFx2_ASAP7_75t_L g1038 ( .A(n_524), .Y(n_1038) );
BUFx3_ASAP7_75t_L g1276 ( .A(n_524), .Y(n_1276) );
INVx1_ASAP7_75t_L g765 ( .A(n_527), .Y(n_765) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g1194 ( .A(n_528), .Y(n_1194) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_L g1021 ( .A(n_529), .Y(n_1021) );
A2O1A1Ixp33_ASAP7_75t_L g1691 ( .A1(n_533), .A2(n_1692), .B(n_1693), .C(n_1694), .Y(n_1691) );
AND4x1_ASAP7_75t_L g1179 ( .A(n_535), .B(n_1180), .C(n_1186), .D(n_1189), .Y(n_1179) );
NAND3xp33_ASAP7_75t_L g1200 ( .A(n_535), .B(n_1201), .C(n_1209), .Y(n_1200) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NOR3xp33_ASAP7_75t_L g931 ( .A(n_536), .B(n_932), .C(n_946), .Y(n_931) );
INVx3_ASAP7_75t_L g1026 ( .A(n_536), .Y(n_1026) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_538), .Y(n_652) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_595), .Y(n_539) );
AOI211xp5_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_543), .B(n_544), .C(n_552), .Y(n_541) );
INVx2_ASAP7_75t_L g720 ( .A(n_542), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_542), .A2(n_1053), .B1(n_1055), .B2(n_1061), .Y(n_1052) );
AOI221xp5_ASAP7_75t_L g1267 ( .A1(n_542), .A2(n_712), .B1(n_1262), .B2(n_1268), .C(n_1271), .Y(n_1267) );
AOI221xp5_ASAP7_75t_L g1303 ( .A1(n_542), .A2(n_712), .B1(n_1304), .B2(n_1305), .C(n_1309), .Y(n_1303) );
AOI211xp5_ASAP7_75t_L g1423 ( .A1(n_542), .A2(n_1424), .B(n_1425), .C(n_1426), .Y(n_1423) );
INVx4_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_546), .A2(n_548), .B1(n_886), .B2(n_887), .Y(n_885) );
AOI221xp5_ASAP7_75t_L g1049 ( .A1(n_546), .A2(n_548), .B1(n_698), .B2(n_1050), .C(n_1051), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_546), .A2(n_548), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_546), .A2(n_548), .B1(n_1335), .B2(n_1336), .Y(n_1334) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_548), .Y(n_697) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_549), .Y(n_698) );
OR2x6_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g583 ( .A(n_550), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g1296 ( .A1(n_550), .A2(n_588), .B1(n_851), .B2(n_1297), .C(n_1298), .Y(n_1296) );
INVx1_ASAP7_75t_L g1694 ( .A(n_551), .Y(n_1694) );
OR2x6_ASAP7_75t_SL g553 ( .A(n_554), .B(n_556), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_555), .Y(n_713) );
INVx1_ASAP7_75t_L g741 ( .A(n_556), .Y(n_741) );
INVx3_ASAP7_75t_L g843 ( .A(n_556), .Y(n_843) );
BUFx2_ASAP7_75t_L g1015 ( .A(n_556), .Y(n_1015) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_558), .B(n_800), .Y(n_1145) );
NOR3xp33_ASAP7_75t_SL g559 ( .A(n_560), .B(n_574), .C(n_580), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g715 ( .A(n_563), .Y(n_715) );
INVx2_ASAP7_75t_L g1294 ( .A(n_563), .Y(n_1294) );
INVx2_ASAP7_75t_L g1347 ( .A(n_563), .Y(n_1347) );
BUFx6f_ASAP7_75t_L g1350 ( .A(n_563), .Y(n_1350) );
BUFx6f_ASAP7_75t_L g1712 ( .A(n_563), .Y(n_1712) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g899 ( .A(n_566), .Y(n_899) );
INVx1_ASAP7_75t_L g1703 ( .A(n_566), .Y(n_1703) );
OAI221xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_570), .B2(n_572), .C(n_573), .Y(n_567) );
INVx2_ASAP7_75t_L g940 ( .A(n_568), .Y(n_940) );
INVx2_ASAP7_75t_R g942 ( .A(n_568), .Y(n_942) );
INVx1_ASAP7_75t_L g1020 ( .A(n_568), .Y(n_1020) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_569), .A2(n_649), .B1(n_650), .B2(n_651), .Y(n_648) );
INVx2_ASAP7_75t_L g1012 ( .A(n_570), .Y(n_1012) );
INVx2_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_571), .B(n_1308), .Y(n_1307) );
BUFx3_ASAP7_75t_L g1354 ( .A(n_571), .Y(n_1354) );
INVx1_ASAP7_75t_L g1397 ( .A(n_571), .Y(n_1397) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_572), .A2(n_627), .B1(n_628), .B2(n_629), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g889 ( .A1(n_573), .A2(n_710), .B1(n_854), .B2(n_890), .C(n_891), .Y(n_889) );
OAI221xp5_ASAP7_75t_L g1277 ( .A1(n_573), .A2(n_754), .B1(n_861), .B2(n_1242), .C(n_1246), .Y(n_1277) );
OAI21xp33_ASAP7_75t_L g1429 ( .A1(n_573), .A2(n_710), .B(n_1430), .Y(n_1429) );
OAI221xp5_ASAP7_75t_L g1709 ( .A1(n_573), .A2(n_899), .B1(n_1710), .B2(n_1711), .C(n_1713), .Y(n_1709) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_576), .A2(n_579), .B1(n_882), .B2(n_883), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_576), .A2(n_579), .B1(n_1356), .B2(n_1357), .Y(n_1355) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx2_ASAP7_75t_SL g767 ( .A(n_586), .Y(n_767) );
INVx3_ASAP7_75t_L g894 ( .A(n_586), .Y(n_894) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx3_ASAP7_75t_L g751 ( .A(n_587), .Y(n_751) );
BUFx4f_ASAP7_75t_L g851 ( .A(n_587), .Y(n_851) );
BUFx3_ASAP7_75t_L g1269 ( .A(n_587), .Y(n_1269) );
INVx3_ASAP7_75t_L g707 ( .A(n_588), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g897 ( .A1(n_588), .A2(n_751), .B1(n_898), .B2(n_899), .C(n_900), .Y(n_897) );
OAI221xp5_ASAP7_75t_L g1115 ( .A1(n_588), .A2(n_1116), .B1(n_1118), .B2(n_1119), .C(n_1121), .Y(n_1115) );
OAI221xp5_ASAP7_75t_L g1279 ( .A1(n_588), .A2(n_751), .B1(n_754), .B2(n_1237), .C(n_1248), .Y(n_1279) );
OAI221xp5_ASAP7_75t_L g1437 ( .A1(n_588), .A2(n_751), .B1(n_754), .B2(n_1438), .C(n_1439), .Y(n_1437) );
OAI221xp5_ASAP7_75t_L g1701 ( .A1(n_588), .A2(n_1269), .B1(n_1702), .B2(n_1703), .C(n_1704), .Y(n_1701) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g867 ( .A(n_589), .B(n_634), .Y(n_867) );
OR2x6_ASAP7_75t_L g944 ( .A(n_589), .B(n_634), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g722 ( .A(n_592), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_592), .B(n_909), .Y(n_908) );
HB1xp67_ASAP7_75t_L g1068 ( .A(n_592), .Y(n_1068) );
AOI222xp33_ASAP7_75t_L g1093 ( .A1(n_592), .A2(n_598), .B1(n_1094), .B2(n_1095), .C1(n_1097), .C2(n_1098), .Y(n_1093) );
NAND2xp33_ASAP7_75t_SL g1282 ( .A(n_592), .B(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1375 ( .A(n_592), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_592), .B(n_1446), .Y(n_1445) );
AOI22xp33_ASAP7_75t_SL g1728 ( .A1(n_592), .A2(n_598), .B1(n_1729), .B2(n_1730), .Y(n_1728) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_621), .Y(n_595) );
AOI211xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_599), .C(n_616), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_598), .B(n_661), .Y(n_660) );
INVx3_ASAP7_75t_L g878 ( .A(n_598), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_598), .B(n_1265), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_598), .B(n_1308), .Y(n_1311) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_601), .A2(n_667), .B1(n_668), .B2(n_669), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g910 ( .A1(n_601), .A2(n_911), .B(n_912), .Y(n_910) );
INVxp67_ASAP7_75t_L g1065 ( .A(n_601), .Y(n_1065) );
INVx1_ASAP7_75t_L g1096 ( .A(n_601), .Y(n_1096) );
AOI222xp33_ASAP7_75t_L g1260 ( .A1(n_601), .A2(n_637), .B1(n_669), .B2(n_1261), .C1(n_1262), .C2(n_1263), .Y(n_1260) );
AOI211xp5_ASAP7_75t_L g1377 ( .A1(n_601), .A2(n_1378), .B(n_1379), .C(n_1380), .Y(n_1377) );
AOI222xp33_ASAP7_75t_L g1442 ( .A1(n_601), .A2(n_637), .B1(n_669), .B2(n_1424), .C1(n_1443), .C2(n_1444), .Y(n_1442) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
AOI332xp33_ASAP7_75t_L g1313 ( .A1(n_602), .A2(n_604), .A3(n_638), .B1(n_639), .B2(n_669), .B3(n_1304), .C1(n_1314), .C2(n_1315), .Y(n_1313) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_614), .B2(n_615), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_608), .A2(n_615), .B1(n_681), .B2(n_682), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_608), .A2(n_615), .B1(n_1103), .B2(n_1105), .Y(n_1141) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_SL g1258 ( .A(n_609), .Y(n_1258) );
HB1xp67_ASAP7_75t_L g1381 ( .A(n_609), .Y(n_1381) );
NAND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g620 ( .A(n_610), .Y(n_620) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_618), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g1076 ( .A1(n_618), .A2(n_1077), .B(n_1085), .Y(n_1076) );
OAI21xp5_ASAP7_75t_SL g1127 ( .A1(n_618), .A2(n_1128), .B(n_1130), .Y(n_1127) );
OAI21xp5_ASAP7_75t_L g1721 ( .A1(n_618), .A2(n_1140), .B(n_1722), .Y(n_1721) );
OR2x6_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx4_ASAP7_75t_L g966 ( .A(n_619), .Y(n_966) );
BUFx4f_ASAP7_75t_L g1133 ( .A(n_619), .Y(n_1133) );
BUFx4f_ASAP7_75t_L g1138 ( .A(n_619), .Y(n_1138) );
BUFx4f_ASAP7_75t_L g1156 ( .A(n_619), .Y(n_1156) );
BUFx6f_ASAP7_75t_L g1322 ( .A(n_619), .Y(n_1322) );
BUFx4f_ASAP7_75t_L g1451 ( .A(n_619), .Y(n_1451) );
AOI322xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_625), .A3(n_631), .B1(n_636), .B2(n_637), .C1(n_640), .C2(n_643), .Y(n_621) );
BUFx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_627), .A2(n_1236), .B1(n_1237), .B2(n_1238), .Y(n_1235) );
INVx5_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx6_ASAP7_75t_L g1075 ( .A(n_630), .Y(n_1075) );
OAI33xp33_ASAP7_75t_L g1449 ( .A1(n_632), .A2(n_1254), .A3(n_1450), .B1(n_1453), .B2(n_1455), .B3(n_1458), .Y(n_1449) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI31xp33_ASAP7_75t_L g672 ( .A1(n_633), .A2(n_673), .A3(n_675), .B(n_679), .Y(n_672) );
INVx4_ASAP7_75t_L g918 ( .A(n_633), .Y(n_918) );
INVx2_ASAP7_75t_L g1086 ( .A(n_633), .Y(n_1086) );
INVx2_ASAP7_75t_L g1234 ( .A(n_633), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g1717 ( .A(n_633), .Y(n_1717) );
AND2x4_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g800 ( .A(n_634), .Y(n_800) );
AOI332xp33_ASAP7_75t_L g913 ( .A1(n_637), .A2(n_640), .A3(n_914), .B1(n_916), .B2(n_917), .B3(n_919), .C1(n_920), .C2(n_922), .Y(n_913) );
AOI322xp5_ASAP7_75t_L g1359 ( .A1(n_637), .A2(n_640), .A3(n_1360), .B1(n_1361), .B2(n_1365), .C1(n_1366), .C2(n_1371), .Y(n_1359) );
AND2x4_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_640), .B(n_684), .C(n_687), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g1069 ( .A1(n_640), .A2(n_1070), .B(n_1076), .C(n_1087), .Y(n_1069) );
CKINVDCx5p33_ASAP7_75t_R g1140 ( .A(n_640), .Y(n_1140) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g981 ( .A(n_645), .Y(n_981) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g1458 ( .A1(n_649), .A2(n_1238), .B1(n_1434), .B2(n_1459), .Y(n_1458) );
OAI22xp5_ASAP7_75t_L g1453 ( .A1(n_651), .A2(n_1432), .B1(n_1439), .B2(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g869 ( .A(n_653), .Y(n_869) );
XNOR2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_725), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI21x1_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_658), .B(n_724), .Y(n_656) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_657), .B(n_660), .C(n_662), .D(n_692), .Y(n_724) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .C(n_692), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_671), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_667), .A2(n_712), .B1(n_714), .B2(n_719), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g907 ( .A1(n_669), .A2(n_679), .B(n_887), .Y(n_907) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND3xp33_ASAP7_75t_SL g671 ( .A(n_672), .B(n_680), .C(n_683), .Y(n_671) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_676), .Y(n_984) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx3_ASAP7_75t_L g821 ( .A(n_677), .Y(n_821) );
NOR3xp33_ASAP7_75t_L g1316 ( .A(n_679), .B(n_1317), .C(n_1324), .Y(n_1316) );
OR3x1_ASAP7_75t_L g1447 ( .A(n_679), .B(n_1448), .C(n_1449), .Y(n_1447) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
BUFx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g1410 ( .A(n_691), .Y(n_1410) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_699), .C(n_711), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g1272 ( .A(n_698), .B(n_1273), .C(n_1278), .Y(n_1272) );
NOR3xp33_ASAP7_75t_L g1289 ( .A(n_698), .B(n_1290), .C(n_1295), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B1(n_706), .B2(n_708), .Y(n_699) );
BUFx2_ASAP7_75t_L g1016 ( .A(n_701), .Y(n_1016) );
BUFx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_710), .A2(n_902), .B1(n_903), .B2(n_904), .Y(n_901) );
INVx1_ASAP7_75t_L g1685 ( .A(n_712), .Y(n_1685) );
BUFx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g1054 ( .A(n_713), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_716), .A2(n_1123), .B1(n_1124), .B2(n_1125), .Y(n_1122) );
CKINVDCx8_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
INVx3_ASAP7_75t_L g896 ( .A(n_717), .Y(n_896) );
INVx3_ASAP7_75t_L g1301 ( .A(n_717), .Y(n_1301) );
INVx1_ASAP7_75t_L g1433 ( .A(n_717), .Y(n_1433) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_802), .B1(n_803), .B2(n_868), .Y(n_725) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND3x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_770), .C(n_773), .Y(n_728) );
AOI211xp5_ASAP7_75t_SL g729 ( .A1(n_730), .A2(n_731), .B(n_733), .C(n_737), .Y(n_729) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B1(n_742), .B2(n_743), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI221xp5_ASAP7_75t_L g756 ( .A1(n_743), .A2(n_757), .B1(n_758), .B2(n_761), .C(n_762), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g1696 ( .A1(n_743), .A2(n_1697), .B1(n_1698), .B2(n_1700), .Y(n_1696) );
BUFx3_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g858 ( .A(n_744), .Y(n_858) );
BUFx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI33xp33_ASAP7_75t_L g849 ( .A1(n_746), .A2(n_850), .A3(n_855), .B1(n_860), .B2(n_864), .B3(n_867), .Y(n_849) );
BUFx4f_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B1(n_753), .B2(n_755), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI221xp5_ASAP7_75t_L g788 ( .A1(n_752), .A2(n_777), .B1(n_789), .B2(n_793), .C(n_794), .Y(n_788) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_754), .A2(n_851), .B1(n_865), .B2(n_866), .Y(n_864) );
INVx2_ASAP7_75t_L g1117 ( .A(n_754), .Y(n_1117) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_760), .A2(n_1300), .B1(n_1301), .B2(n_1302), .Y(n_1299) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_763), .A2(n_938), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
OR2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
OR2x6_ASAP7_75t_L g1024 ( .A(n_767), .B(n_768), .Y(n_1024) );
INVx2_ASAP7_75t_SL g1340 ( .A(n_767), .Y(n_1340) );
INVxp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_L g842 ( .A(n_769), .B(n_843), .Y(n_842) );
OAI31xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_785), .A3(n_796), .B(n_798), .Y(n_773) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g1168 ( .A(n_782), .Y(n_1168) );
HB1xp67_ASAP7_75t_SL g982 ( .A(n_783), .Y(n_982) );
INVxp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
OAI22xp33_ASAP7_75t_L g1072 ( .A1(n_791), .A2(n_1073), .B1(n_1074), .B2(n_1075), .Y(n_1072) );
INVx3_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx6f_ASAP7_75t_L g994 ( .A(n_792), .Y(n_994) );
O2A1O1Ixp33_ASAP7_75t_SL g1152 ( .A1(n_798), .A2(n_1153), .B(n_1165), .C(n_1173), .Y(n_1152) );
AOI21xp5_ASAP7_75t_SL g1401 ( .A1(n_798), .A2(n_1402), .B(n_1418), .Y(n_1401) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g1034 ( .A1(n_799), .A2(n_1035), .B(n_1062), .Y(n_1034) );
INVx2_ASAP7_75t_L g1281 ( .A(n_799), .Y(n_1281) );
OAI31xp33_ASAP7_75t_SL g1331 ( .A1(n_799), .A2(n_1332), .A3(n_1333), .B(n_1337), .Y(n_1331) );
BUFx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
AOI21xp5_ASAP7_75t_SL g808 ( .A1(n_800), .A2(n_809), .B(n_830), .Y(n_808) );
INVx1_ASAP7_75t_L g1715 ( .A(n_800), .Y(n_1715) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_837), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_817), .B(n_818), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g1450 ( .A1(n_811), .A2(n_1430), .B1(n_1451), .B2(n_1452), .Y(n_1450) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g1137 ( .A(n_812), .Y(n_1137) );
INVx4_ASAP7_75t_L g1241 ( .A(n_812), .Y(n_1241) );
INVx4_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_824), .Y(n_818) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g1221 ( .A(n_821), .Y(n_1221) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_825), .A2(n_827), .B1(n_828), .B2(n_829), .Y(n_824) );
AOI222xp33_ASAP7_75t_L g1214 ( .A1(n_825), .A2(n_1210), .B1(n_1211), .B2(n_1215), .C1(n_1216), .C2(n_1217), .Y(n_1214) );
INVx1_ASAP7_75t_L g1417 ( .A(n_825), .Y(n_1417) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_829), .A2(n_841), .B1(n_842), .B2(n_844), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_830) );
NAND3xp33_ASAP7_75t_SL g837 ( .A(n_838), .B(n_840), .C(n_845), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_842), .A2(n_1171), .B1(n_1172), .B2(n_1175), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_842), .A2(n_1175), .B1(n_1223), .B2(n_1224), .Y(n_1226) );
INVx2_ASAP7_75t_L g861 ( .A(n_843), .Y(n_861) );
INVx2_ASAP7_75t_L g1306 ( .A(n_843), .Y(n_1306) );
NOR2xp33_ASAP7_75t_SL g845 ( .A(n_846), .B(n_849), .Y(n_845) );
OAI22xp33_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B1(n_853), .B2(n_854), .Y(n_850) );
INVx1_ASAP7_75t_L g1120 ( .A(n_851), .Y(n_1120) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_857), .A2(n_861), .B1(n_862), .B2(n_863), .Y(n_860) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
BUFx2_ASAP7_75t_L g1057 ( .A(n_858), .Y(n_1057) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
XNOR2xp5_ASAP7_75t_L g872 ( .A(n_873), .B(n_973), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
XNOR2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_924), .Y(n_874) );
XOR2x2_ASAP7_75t_L g875 ( .A(n_876), .B(n_923), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_877), .B(n_906), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_892), .B1(n_897), .B2(n_901), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_894), .B1(n_895), .B2(n_896), .Y(n_892) );
BUFx4f_ASAP7_75t_SL g1707 ( .A(n_894), .Y(n_1707) );
OAI22xp5_ASAP7_75t_L g1280 ( .A1(n_896), .A2(n_1019), .B1(n_1240), .B2(n_1253), .Y(n_1280) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
NAND4xp25_ASAP7_75t_SL g906 ( .A(n_907), .B(n_908), .C(n_910), .D(n_913), .Y(n_906) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_917), .Y(n_1129) );
INVx2_ASAP7_75t_SL g917 ( .A(n_918), .Y(n_917) );
NAND3xp33_ASAP7_75t_SL g925 ( .A(n_926), .B(n_931), .C(n_948), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_930), .B(n_1096), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_933), .B(n_936), .Y(n_932) );
HB1xp67_ASAP7_75t_L g1345 ( .A(n_938), .Y(n_1345) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
OAI21xp5_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_960), .B(n_969), .Y(n_948) );
BUFx2_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
OAI211xp5_ASAP7_75t_SL g963 ( .A1(n_964), .A2(n_965), .B(n_967), .C(n_968), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g1239 ( .A1(n_965), .A2(n_1240), .B1(n_1241), .B2(n_1242), .Y(n_1239) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx2_ASAP7_75t_L g1082 ( .A(n_966), .Y(n_1082) );
INVx1_ASAP7_75t_L g1457 ( .A(n_966), .Y(n_1457) );
AOI21xp5_ASAP7_75t_L g1212 ( .A1(n_969), .A2(n_1213), .B(n_1225), .Y(n_1212) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
OAI21xp33_ASAP7_75t_L g1099 ( .A1(n_970), .A2(n_1100), .B(n_1114), .Y(n_1099) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
BUFx2_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_972), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1310 ( .A(n_972), .Y(n_1310) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
NAND3xp33_ASAP7_75t_SL g975 ( .A(n_976), .B(n_1001), .C(n_1004), .Y(n_975) );
OAI21xp33_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_991), .B(n_1000), .Y(n_976) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_987), .B1(n_988), .B2(n_989), .Y(n_985) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
OAI221xp5_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_995), .B1(n_996), .B2(n_997), .C(n_998), .Y(n_992) );
OAI22xp5_ASAP7_75t_SL g1368 ( .A1(n_993), .A2(n_1341), .B1(n_1369), .B2(n_1370), .Y(n_1368) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx2_ASAP7_75t_L g1161 ( .A(n_994), .Y(n_1161) );
INVx3_ASAP7_75t_L g1454 ( .A(n_994), .Y(n_1454) );
NOR3xp33_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1023), .C(n_1025), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1009), .Y(n_1005) );
BUFx2_ASAP7_75t_SL g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx2_ASAP7_75t_SL g1025 ( .A(n_1026), .Y(n_1025) );
NAND3xp33_ASAP7_75t_SL g1390 ( .A(n_1026), .B(n_1391), .C(n_1394), .Y(n_1390) );
AOI22xp5_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1029), .B1(n_1325), .B2(n_1326), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
XNOR2x1_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1147), .Y(n_1030) );
XNOR2x2_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1090), .Y(n_1031) );
AOI21xp5_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1088), .B(n_1089), .Y(n_1032) );
AND3x1_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1063), .C(n_1069), .Y(n_1033) );
AOI31xp33_ASAP7_75t_L g1089 ( .A1(n_1034), .A2(n_1063), .A3(n_1069), .B(n_1088), .Y(n_1089) );
NAND3xp33_ASAP7_75t_SL g1035 ( .A(n_1036), .B(n_1049), .C(n_1052), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1039), .B1(n_1043), .B2(n_1046), .Y(n_1036) );
INVx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
BUFx2_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1048), .Y(n_1275) );
INVxp67_ASAP7_75t_L g1101 ( .A(n_1053), .Y(n_1101) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1705 ( .A1(n_1056), .A2(n_1706), .B1(n_1707), .B2(n_1708), .Y(n_1705) );
INVx3_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1066), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1068), .Y(n_1066) );
OAI221xp5_ASAP7_75t_L g1722 ( .A1(n_1075), .A2(n_1700), .B1(n_1710), .B2(n_1723), .C(n_1725), .Y(n_1722) );
OAI221xp5_ASAP7_75t_L g1077 ( .A1(n_1078), .A2(n_1081), .B1(n_1082), .B2(n_1083), .C(n_1084), .Y(n_1077) );
INVx3_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx2_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
OAI221xp5_ASAP7_75t_L g1318 ( .A1(n_1080), .A2(n_1133), .B1(n_1293), .B2(n_1300), .C(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1085), .Y(n_1371) );
BUFx6f_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
NAND3xp33_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1099), .C(n_1126), .Y(n_1092) );
OAI211xp5_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1102), .B(n_1104), .C(n_1107), .Y(n_1100) );
OAI211xp5_ASAP7_75t_L g1107 ( .A1(n_1108), .A2(n_1109), .B(n_1112), .C(n_1113), .Y(n_1107) );
OAI221xp5_ASAP7_75t_L g1136 ( .A1(n_1108), .A2(n_1118), .B1(n_1137), .B2(n_1138), .C(n_1139), .Y(n_1136) );
HB1xp67_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx2_ASAP7_75t_L g1270 ( .A(n_1111), .Y(n_1270) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
OAI221xp5_ASAP7_75t_L g1130 ( .A1(n_1124), .A2(n_1131), .B1(n_1132), .B2(n_1133), .C(n_1134), .Y(n_1130) );
NOR3xp33_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1135), .C(n_1142), .Y(n_1126) );
INVxp67_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
XNOR2xp5_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1227), .Y(n_1147) );
XNOR2xp5_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1195), .Y(n_1148) );
NOR2x1p5_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1176), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g1159 ( .A1(n_1160), .A2(n_1161), .B1(n_1162), .B2(n_1163), .Y(n_1159) );
BUFx3_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1179), .Y(n_1176) );
AOI22xp5_ASAP7_75t_L g1180 ( .A1(n_1181), .A2(n_1182), .B1(n_1184), .B2(n_1185), .Y(n_1180) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1188), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1212), .Y(n_1196) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1205), .Y(n_1688) );
NAND3xp33_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1218), .C(n_1222), .Y(n_1213) );
AOI222xp33_ASAP7_75t_L g1412 ( .A1(n_1215), .A2(n_1392), .B1(n_1393), .B2(n_1413), .C1(n_1415), .C2(n_1416), .Y(n_1412) );
XNOR2x1_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1284), .Y(n_1227) );
XNOR2x1_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1230), .Y(n_1228) );
NOR2x1_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1266), .Y(n_1230) );
NAND3xp33_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1260), .C(n_1264), .Y(n_1231) );
NOR2xp33_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1256), .Y(n_1232) );
OAI33xp33_ASAP7_75t_L g1233 ( .A1(n_1234), .A2(n_1235), .A3(n_1239), .B1(n_1243), .B2(n_1249), .B3(n_1254), .Y(n_1233) );
OAI22xp5_ASAP7_75t_SL g1317 ( .A1(n_1234), .A2(n_1318), .B1(n_1320), .B2(n_1321), .Y(n_1317) );
OAI22xp5_ASAP7_75t_L g1249 ( .A1(n_1238), .A2(n_1250), .B1(n_1252), .B2(n_1253), .Y(n_1249) );
HB1xp67_ASAP7_75t_L g1370 ( .A(n_1238), .Y(n_1370) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_1244), .A2(n_1246), .B1(n_1247), .B2(n_1248), .Y(n_1243) );
OAI22xp5_ASAP7_75t_L g1455 ( .A1(n_1244), .A2(n_1438), .B1(n_1456), .B2(n_1457), .Y(n_1455) );
INVx4_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g1719 ( .A1(n_1247), .A2(n_1697), .B1(n_1706), .B2(n_1720), .Y(n_1719) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVx2_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
A2O1A1Ixp33_ASAP7_75t_L g1266 ( .A1(n_1267), .A2(n_1272), .B(n_1281), .C(n_1282), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g1431 ( .A1(n_1269), .A2(n_1432), .B1(n_1433), .B2(n_1434), .Y(n_1431) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
AOI221xp5_ASAP7_75t_SL g1686 ( .A1(n_1276), .A2(n_1687), .B1(n_1688), .B2(n_1689), .C(n_1690), .Y(n_1686) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1281), .Y(n_1440) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
XNOR2x1_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1287), .Y(n_1285) );
OR2x2_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1312), .Y(n_1287) );
A2O1A1Ixp33_ASAP7_75t_L g1288 ( .A1(n_1289), .A2(n_1303), .B(n_1310), .C(n_1311), .Y(n_1288) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
OA22x2_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1383), .B1(n_1384), .B2(n_1460), .Y(n_1326) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1327), .Y(n_1460) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
NOR2x1_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1358), .Y(n_1329) );
NAND3xp33_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1348), .C(n_1355), .Y(n_1337) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_1339), .A2(n_1341), .B1(n_1342), .B2(n_1343), .C(n_1344), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
OAI221xp5_ASAP7_75t_L g1348 ( .A1(n_1342), .A2(n_1349), .B1(n_1351), .B2(n_1352), .C(n_1353), .Y(n_1348) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1372), .Y(n_1358) );
INVx1_ASAP7_75t_SL g1363 ( .A(n_1364), .Y(n_1363) );
AOI21xp5_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1374), .B(n_1376), .Y(n_1372) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
XNOR2xp5_ASAP7_75t_L g1384 ( .A(n_1385), .B(n_1420), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1387), .B(n_1401), .Y(n_1386) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
NAND3xp33_ASAP7_75t_SL g1402 ( .A(n_1403), .B(n_1406), .C(n_1412), .Y(n_1402) );
INVx2_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
AOI211x1_ASAP7_75t_L g1421 ( .A1(n_1422), .A2(n_1440), .B(n_1441), .C(n_1447), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1427), .Y(n_1422) );
NOR3xp33_ASAP7_75t_L g1427 ( .A(n_1428), .B(n_1435), .C(n_1436), .Y(n_1427) );
OAI221xp5_ASAP7_75t_L g1461 ( .A1(n_1462), .A2(n_1676), .B1(n_1679), .B2(n_1731), .C(n_1734), .Y(n_1461) );
AOI211xp5_ASAP7_75t_L g1462 ( .A1(n_1463), .A2(n_1588), .B(n_1592), .C(n_1651), .Y(n_1462) );
NAND5xp2_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1523), .C(n_1539), .D(n_1558), .E(n_1580), .Y(n_1463) );
AOI211xp5_ASAP7_75t_L g1464 ( .A1(n_1465), .A2(n_1495), .B(n_1504), .C(n_1516), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1466), .B(n_1480), .Y(n_1465) );
INVx2_ASAP7_75t_L g1514 ( .A(n_1466), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1466), .B(n_1482), .Y(n_1533) );
AOI311xp33_ASAP7_75t_L g1558 ( .A1(n_1466), .A2(n_1559), .A3(n_1564), .B(n_1568), .C(n_1576), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1584 ( .A(n_1466), .B(n_1517), .Y(n_1584) );
OR2x2_ASAP7_75t_L g1610 ( .A(n_1466), .B(n_1611), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1466), .B(n_1491), .Y(n_1630) );
NAND2xp5_ASAP7_75t_L g1649 ( .A(n_1466), .B(n_1487), .Y(n_1649) );
OR2x2_ASAP7_75t_L g1666 ( .A(n_1466), .B(n_1487), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1467), .B(n_1475), .Y(n_1466) );
AND2x4_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1470), .Y(n_1468) );
AND2x6_ASAP7_75t_L g1473 ( .A(n_1469), .B(n_1474), .Y(n_1473) );
AND2x6_ASAP7_75t_L g1476 ( .A(n_1469), .B(n_1477), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1478 ( .A(n_1469), .B(n_1479), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1469), .B(n_1479), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1469), .B(n_1479), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1472), .Y(n_1470) );
INVx2_ASAP7_75t_L g1678 ( .A(n_1473), .Y(n_1678) );
HB1xp67_ASAP7_75t_L g1748 ( .A(n_1474), .Y(n_1748) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1485), .Y(n_1480) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1481), .Y(n_1512) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1481), .B(n_1566), .Y(n_1565) );
OR2x2_ASAP7_75t_L g1577 ( .A(n_1481), .B(n_1521), .Y(n_1577) );
OAI21xp33_ASAP7_75t_L g1598 ( .A1(n_1481), .A2(n_1599), .B(n_1600), .Y(n_1598) );
OAI332xp33_ASAP7_75t_L g1643 ( .A1(n_1481), .A2(n_1584), .A3(n_1644), .B1(n_1646), .B2(n_1647), .B3(n_1648), .C1(n_1649), .C2(n_1650), .Y(n_1643) );
OR2x2_ASAP7_75t_L g1644 ( .A(n_1481), .B(n_1645), .Y(n_1644) );
CKINVDCx5p33_ASAP7_75t_R g1481 ( .A(n_1482), .Y(n_1481) );
NOR2xp33_ASAP7_75t_L g1542 ( .A(n_1482), .B(n_1543), .Y(n_1542) );
INVx3_ASAP7_75t_L g1547 ( .A(n_1482), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1482), .B(n_1575), .Y(n_1581) );
NOR2xp33_ASAP7_75t_L g1607 ( .A(n_1482), .B(n_1550), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1611 ( .A(n_1482), .B(n_1485), .Y(n_1611) );
OR2x2_ASAP7_75t_L g1665 ( .A(n_1482), .B(n_1666), .Y(n_1665) );
AND2x4_ASAP7_75t_SL g1482 ( .A(n_1483), .B(n_1484), .Y(n_1482) );
NAND2xp5_ASAP7_75t_L g1663 ( .A(n_1485), .B(n_1533), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1486), .B(n_1491), .Y(n_1485) );
OR2x2_ASAP7_75t_L g1517 ( .A(n_1486), .B(n_1492), .Y(n_1517) );
AOI322xp5_ASAP7_75t_L g1580 ( .A1(n_1486), .A2(n_1566), .A3(n_1581), .B1(n_1582), .B2(n_1583), .C1(n_1585), .C2(n_1587), .Y(n_1580) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1487), .B(n_1492), .Y(n_1515) );
NOR2xp33_ASAP7_75t_L g1531 ( .A(n_1487), .B(n_1532), .Y(n_1531) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_1487), .B(n_1551), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1487), .B(n_1514), .Y(n_1602) );
NOR3xp33_ASAP7_75t_SL g1636 ( .A(n_1487), .B(n_1512), .C(n_1588), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1489), .Y(n_1487) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1492), .Y(n_1545) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1492), .Y(n_1551) );
NAND2xp5_ASAP7_75t_L g1645 ( .A(n_1492), .B(n_1514), .Y(n_1645) );
NAND2x1_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1494), .Y(n_1492) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1495), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1500), .Y(n_1495) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1497), .Y(n_1519) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1497), .Y(n_1530) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1497), .B(n_1500), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_1497), .B(n_1501), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1499), .Y(n_1497) );
OR2x2_ASAP7_75t_L g1554 ( .A(n_1500), .B(n_1506), .Y(n_1554) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1500), .B(n_1507), .Y(n_1567) );
HB1xp67_ASAP7_75t_SL g1616 ( .A(n_1500), .Y(n_1616) );
NAND2xp5_ASAP7_75t_L g1648 ( .A(n_1500), .B(n_1605), .Y(n_1648) );
CKINVDCx5p33_ASAP7_75t_R g1500 ( .A(n_1501), .Y(n_1500) );
NAND2xp5_ASAP7_75t_L g1521 ( .A(n_1501), .B(n_1522), .Y(n_1521) );
OR2x2_ASAP7_75t_L g1526 ( .A(n_1501), .B(n_1507), .Y(n_1526) );
HB1xp67_ASAP7_75t_SL g1552 ( .A(n_1501), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1501), .B(n_1519), .Y(n_1587) );
AND2x4_ASAP7_75t_L g1501 ( .A(n_1502), .B(n_1503), .Y(n_1501) );
NOR2xp33_ASAP7_75t_L g1504 ( .A(n_1505), .B(n_1510), .Y(n_1504) );
OAI32xp33_ASAP7_75t_L g1640 ( .A1(n_1505), .A2(n_1506), .A3(n_1570), .B1(n_1600), .B2(n_1641), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1650 ( .A(n_1505), .B(n_1536), .Y(n_1650) );
INVx2_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_1506), .B(n_1586), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1656 ( .A(n_1506), .B(n_1623), .Y(n_1656) );
INVx2_ASAP7_75t_SL g1506 ( .A(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1507), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1507), .B(n_1547), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1508), .B(n_1509), .Y(n_1507) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
O2A1O1Ixp33_ASAP7_75t_L g1606 ( .A1(n_1511), .A2(n_1607), .B(n_1608), .C(n_1609), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1511 ( .A(n_1512), .B(n_1513), .Y(n_1511) );
OR2x2_ASAP7_75t_L g1537 ( .A(n_1512), .B(n_1538), .Y(n_1537) );
AOI221xp5_ASAP7_75t_L g1523 ( .A1(n_1513), .A2(n_1524), .B1(n_1527), .B2(n_1531), .C(n_1534), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1514), .B(n_1515), .Y(n_1513) );
OR2x2_ASAP7_75t_L g1538 ( .A(n_1514), .B(n_1517), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1544 ( .A(n_1514), .B(n_1545), .Y(n_1544) );
OR2x2_ASAP7_75t_L g1549 ( .A(n_1514), .B(n_1550), .Y(n_1549) );
NAND2xp5_ASAP7_75t_L g1557 ( .A(n_1514), .B(n_1547), .Y(n_1557) );
OR2x2_ASAP7_75t_L g1595 ( .A(n_1514), .B(n_1596), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1514), .B(n_1563), .Y(n_1600) );
OR2x2_ASAP7_75t_L g1659 ( .A(n_1514), .B(n_1556), .Y(n_1659) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1515), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1515), .B(n_1533), .Y(n_1586) );
NAND2xp5_ASAP7_75t_L g1596 ( .A(n_1515), .B(n_1547), .Y(n_1596) );
NOR2xp33_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1518), .Y(n_1516) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1517), .Y(n_1562) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1518), .Y(n_1608) );
NAND2xp5_ASAP7_75t_L g1518 ( .A(n_1519), .B(n_1520), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1519), .B(n_1525), .Y(n_1524) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1519), .Y(n_1575) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1519), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1519), .B(n_1574), .Y(n_1672) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1521), .Y(n_1599) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1521), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_1522), .B(n_1541), .Y(n_1540) );
INVx2_ASAP7_75t_L g1574 ( .A(n_1522), .Y(n_1574) );
NAND2xp5_ASAP7_75t_L g1528 ( .A(n_1525), .B(n_1529), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1525), .B(n_1547), .Y(n_1639) );
INVx2_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
NOR2xp33_ASAP7_75t_L g1674 ( .A(n_1526), .B(n_1547), .Y(n_1674) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
OAI332xp33_ASAP7_75t_L g1625 ( .A1(n_1530), .A2(n_1565), .A3(n_1611), .B1(n_1626), .B2(n_1627), .B3(n_1628), .C1(n_1629), .C2(n_1632), .Y(n_1625) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1533), .B(n_1563), .Y(n_1570) );
NOR2xp33_ASAP7_75t_L g1534 ( .A(n_1535), .B(n_1537), .Y(n_1534) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
AOI21xp33_ASAP7_75t_L g1576 ( .A1(n_1538), .A2(n_1577), .B(n_1578), .Y(n_1576) );
INVx2_ASAP7_75t_L g1621 ( .A(n_1538), .Y(n_1621) );
AOI221xp5_ASAP7_75t_L g1539 ( .A1(n_1540), .A2(n_1542), .B1(n_1546), .B2(n_1552), .C(n_1553), .Y(n_1539) );
OAI31xp33_ASAP7_75t_L g1652 ( .A1(n_1541), .A2(n_1594), .A3(n_1653), .B(n_1655), .Y(n_1652) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
A2O1A1Ixp33_ASAP7_75t_L g1673 ( .A1(n_1545), .A2(n_1633), .B(n_1674), .C(n_1675), .Y(n_1673) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1548), .Y(n_1546) );
NOR2xp33_ASAP7_75t_L g1603 ( .A(n_1547), .B(n_1554), .Y(n_1603) );
CKINVDCx14_ASAP7_75t_R g1620 ( .A(n_1547), .Y(n_1620) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1548), .B(n_1574), .Y(n_1654) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1550), .Y(n_1563) );
A2O1A1Ixp33_ASAP7_75t_L g1593 ( .A1(n_1552), .A2(n_1594), .B(n_1597), .C(n_1605), .Y(n_1593) );
NOR2xp33_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1555), .Y(n_1553) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1554), .Y(n_1582) );
OAI22xp33_ASAP7_75t_L g1662 ( .A1(n_1554), .A2(n_1571), .B1(n_1578), .B2(n_1663), .Y(n_1662) );
OR2x2_ASAP7_75t_L g1555 ( .A(n_1556), .B(n_1557), .Y(n_1555) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1557), .Y(n_1572) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
NOR2xp33_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1563), .Y(n_1561) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_1562), .B(n_1572), .Y(n_1571) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1566), .Y(n_1624) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
OR2x2_ASAP7_75t_L g1613 ( .A(n_1567), .B(n_1614), .Y(n_1613) );
AOI21xp5_ASAP7_75t_L g1568 ( .A1(n_1569), .A2(n_1571), .B(n_1573), .Y(n_1568) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
OAI22xp5_ASAP7_75t_L g1609 ( .A1(n_1573), .A2(n_1610), .B1(n_1612), .B2(n_1613), .Y(n_1609) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1573), .Y(n_1660) );
OR2x2_ASAP7_75t_L g1573 ( .A(n_1574), .B(n_1575), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1574), .B(n_1575), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_1574), .B(n_1586), .Y(n_1585) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1574), .Y(n_1647) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1604 ( .A(n_1582), .B(n_1583), .Y(n_1604) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
NOR2xp33_ASAP7_75t_SL g1632 ( .A(n_1587), .B(n_1633), .Y(n_1632) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1587), .Y(n_1667) );
INVx3_ASAP7_75t_L g1605 ( .A(n_1588), .Y(n_1605) );
NOR2xp33_ASAP7_75t_L g1633 ( .A(n_1588), .B(n_1614), .Y(n_1633) );
NOR3xp33_ASAP7_75t_L g1664 ( .A(n_1588), .B(n_1665), .C(n_1667), .Y(n_1664) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1589), .B(n_1591), .Y(n_1588) );
NAND4xp25_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1606), .C(n_1615), .D(n_1634), .Y(n_1592) );
AOI22xp5_ASAP7_75t_L g1668 ( .A1(n_1594), .A2(n_1623), .B1(n_1669), .B2(n_1672), .Y(n_1668) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1596), .Y(n_1641) );
NAND3xp33_ASAP7_75t_SL g1597 ( .A(n_1598), .B(n_1601), .C(n_1604), .Y(n_1597) );
INVx2_ASAP7_75t_L g1612 ( .A(n_1600), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1623 ( .A(n_1600), .B(n_1620), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1602), .B(n_1603), .Y(n_1601) );
CKINVDCx14_ASAP7_75t_R g1626 ( .A(n_1602), .Y(n_1626) );
CKINVDCx14_ASAP7_75t_R g1627 ( .A(n_1605), .Y(n_1627) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1605), .B(n_1614), .Y(n_1642) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1613), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1613), .B(n_1670), .Y(n_1669) );
AOI211xp5_ASAP7_75t_L g1615 ( .A1(n_1616), .A2(n_1617), .B(n_1618), .C(n_1625), .Y(n_1615) );
AOI21xp33_ASAP7_75t_L g1618 ( .A1(n_1619), .A2(n_1622), .B(n_1624), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1620), .B(n_1621), .Y(n_1619) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1623), .Y(n_1622) );
CKINVDCx14_ASAP7_75t_R g1661 ( .A(n_1627), .Y(n_1661) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1631), .Y(n_1629) );
OAI21xp5_ASAP7_75t_L g1637 ( .A1(n_1630), .A2(n_1638), .B(n_1640), .Y(n_1637) );
INVxp67_ASAP7_75t_SL g1646 ( .A(n_1633), .Y(n_1646) );
AOI221xp5_ASAP7_75t_L g1634 ( .A1(n_1635), .A2(n_1636), .B1(n_1637), .B2(n_1642), .C(n_1643), .Y(n_1634) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
NAND4xp25_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1657), .C(n_1668), .D(n_1673), .Y(n_1651) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
AOI311xp33_ASAP7_75t_L g1657 ( .A1(n_1658), .A2(n_1660), .A3(n_1661), .B(n_1662), .C(n_1664), .Y(n_1657) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1663), .Y(n_1675) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
CKINVDCx20_ASAP7_75t_R g1676 ( .A(n_1677), .Y(n_1676) );
CKINVDCx20_ASAP7_75t_R g1677 ( .A(n_1678), .Y(n_1677) );
INVx2_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
HB1xp67_ASAP7_75t_L g1743 ( .A(n_1682), .Y(n_1743) );
NAND4xp75_ASAP7_75t_L g1682 ( .A(n_1683), .B(n_1716), .C(n_1727), .D(n_1728), .Y(n_1682) );
OAI21x1_ASAP7_75t_L g1683 ( .A1(n_1684), .A2(n_1695), .B(n_1714), .Y(n_1683) );
OAI21xp5_ASAP7_75t_L g1684 ( .A1(n_1685), .A2(n_1686), .B(n_1691), .Y(n_1684) );
OAI22xp5_ASAP7_75t_L g1695 ( .A1(n_1696), .A2(n_1701), .B1(n_1705), .B2(n_1709), .Y(n_1695) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
INVx2_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
AOI211x1_ASAP7_75t_L g1716 ( .A1(n_1717), .A2(n_1718), .B(n_1721), .C(n_1726), .Y(n_1716) );
INVx2_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
INVx2_ASAP7_75t_L g1731 ( .A(n_1732), .Y(n_1731) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
HB1xp67_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
BUFx3_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
INVxp67_ASAP7_75t_SL g1740 ( .A(n_1741), .Y(n_1740) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
INVx2_ASAP7_75t_SL g1745 ( .A(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
OAI21xp5_ASAP7_75t_L g1747 ( .A1(n_1748), .A2(n_1749), .B(n_1750), .Y(n_1747) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
endmodule