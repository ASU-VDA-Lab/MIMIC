module fake_jpeg_5374_n_251 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_5),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_31),
.B(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_20),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_26),
.B(n_18),
.C(n_22),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_57),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_28),
.B1(n_17),
.B2(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_49),
.B1(n_36),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_21),
.B1(n_22),
.B2(n_27),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_36),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_60),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_23),
.B1(n_16),
.B2(n_56),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_69),
.Y(n_84)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_68),
.Y(n_83)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_73),
.Y(n_88)
);

AO21x1_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_59),
.B(n_41),
.Y(n_71)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_39),
.B(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_43),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_16),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_41),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_104),
.Y(n_126)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_91),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_63),
.B(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_74),
.B1(n_78),
.B2(n_67),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_94),
.B1(n_77),
.B2(n_70),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2x1p5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_34),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_95),
.B(n_79),
.Y(n_119)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_97),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_56),
.B1(n_44),
.B2(n_58),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_39),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_65),
.B1(n_75),
.B2(n_60),
.Y(n_108)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_20),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_69),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_106),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_110),
.B(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_109),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_71),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_73),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_65),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_87),
.B1(n_110),
.B2(n_109),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_66),
.B(n_39),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_122),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_66),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_137),
.B1(n_101),
.B2(n_126),
.Y(n_164)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_116),
.B1(n_124),
.B2(n_119),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_99),
.B1(n_82),
.B2(n_104),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_115),
.B1(n_82),
.B2(n_113),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_142),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_123),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_120),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_126),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_150),
.B(n_163),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_106),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_152),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_125),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_138),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_35),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_121),
.C(n_95),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_129),
.C(n_143),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_117),
.B(n_132),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_159),
.A2(n_161),
.B(n_129),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_145),
.A2(n_117),
.B(n_90),
.C(n_88),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_159),
.B1(n_153),
.B2(n_152),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_101),
.B1(n_118),
.B2(n_97),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_15),
.B1(n_29),
.B2(n_24),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_128),
.B(n_83),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_86),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_174),
.B1(n_175),
.B2(n_181),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_172),
.A2(n_182),
.B(n_35),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_179),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_134),
.B1(n_142),
.B2(n_128),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_134),
.B1(n_147),
.B2(n_139),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_155),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_148),
.C(n_135),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_76),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_64),
.B1(n_86),
.B2(n_91),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_35),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_91),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_186),
.B1(n_177),
.B2(n_166),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_29),
.B1(n_24),
.B2(n_25),
.Y(n_186)
);

AOI21x1_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_161),
.B(n_169),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_193),
.B(n_197),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_191),
.B1(n_202),
.B2(n_177),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_178),
.A2(n_158),
.B1(n_157),
.B2(n_155),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_195),
.B(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_155),
.Y(n_198)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_0),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_2),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_200),
.A2(n_2),
.B(n_3),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_171),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_185),
.A2(n_29),
.B1(n_24),
.B2(n_76),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_171),
.C(n_184),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_213),
.C(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_207),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_189),
.B(n_182),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_196),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_191),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_209),
.A2(n_210),
.B(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_199),
.B(n_182),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_214),
.B(n_201),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_35),
.C(n_68),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_2),
.B(n_3),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_216),
.B(n_15),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_221),
.Y(n_228)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_211),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_222),
.B(n_223),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_3),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_194),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_194),
.B(n_192),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_206),
.C(n_207),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_224),
.A2(n_33),
.B(n_30),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_225),
.A2(n_68),
.B1(n_4),
.B2(n_6),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_231),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_226),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_35),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_229),
.B(n_224),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_33),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_229),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_237),
.B(n_15),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_218),
.Y(n_237)
);

OAI21x1_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_33),
.B(n_30),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_SL g241 ( 
.A1(n_239),
.A2(n_236),
.B(n_238),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_12),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_29),
.A3(n_24),
.B1(n_20),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_10),
.C2(n_11),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_6),
.B(n_10),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_247),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_246),
.A2(n_12),
.B(n_25),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_12),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_249),
.Y(n_251)
);


endmodule