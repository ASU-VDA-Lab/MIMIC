module real_jpeg_15525_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_1),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_1),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_1),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_1),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_1),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_1),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_1),
.B(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_1),
.A2(n_4),
.B1(n_304),
.B2(n_306),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_1),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_2),
.Y(n_181)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_2),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_3),
.A2(n_20),
.B(n_22),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_4),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_4),
.B(n_244),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_4),
.B(n_372),
.Y(n_371)
);

AOI31xp33_ASAP7_75t_SL g404 ( 
.A1(n_4),
.A2(n_303),
.A3(n_405),
.B(n_407),
.Y(n_404)
);

NAND2x1_ASAP7_75t_SL g446 ( 
.A(n_4),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_4),
.B(n_112),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_4),
.B(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_4),
.B(n_519),
.Y(n_518)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_5),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_5),
.Y(n_209)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_5),
.Y(n_425)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_6),
.Y(n_112)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_6),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_6),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_6),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_7),
.Y(n_183)
);

NAND2x1_ASAP7_75t_SL g185 ( 
.A(n_7),
.B(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_7),
.B(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g270 ( 
.A(n_7),
.B(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g322 ( 
.A(n_7),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_7),
.B(n_112),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_7),
.B(n_412),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_7),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_8),
.B(n_69),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_8),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_8),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_8),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_8),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_8),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_8),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g369 ( 
.A(n_8),
.B(n_260),
.Y(n_369)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_9),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_9),
.Y(n_228)
);

BUFx4f_ASAP7_75t_L g414 ( 
.A(n_9),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_9),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_10),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_10),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_10),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_10),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_10),
.B(n_510),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_10),
.B(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_10),
.B(n_530),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_11),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_11),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_11),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_11),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_11),
.B(n_568),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_12),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_12),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_13),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_13),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_13),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_13),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_13),
.B(n_226),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_13),
.B(n_260),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_14),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_14),
.Y(n_148)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_14),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_14),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_15),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_15),
.B(n_71),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_15),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_15),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_15),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_15),
.B(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_15),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_15),
.B(n_327),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_16),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_16),
.B(n_97),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_16),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_16),
.B(n_88),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_16),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_16),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_16),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_16),
.B(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g186 ( 
.A(n_18),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_563),
.B(n_571),
.C(n_573),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_120),
.B(n_562),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2x1_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_76),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_27),
.B(n_76),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_58),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_44),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_29),
.B(n_44),
.C(n_58),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_36),
.C(n_39),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_30),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_30),
.A2(n_36),
.B1(n_51),
.B2(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_SL g565 ( 
.A(n_30),
.B(n_46),
.C(n_53),
.Y(n_565)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_34),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_35),
.Y(n_165)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_35),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_68),
.C(n_73),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_36),
.A2(n_62),
.B1(n_73),
.B2(n_74),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_38),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_53),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_46),
.A2(n_52),
.B1(n_567),
.B2(n_571),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_49),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_111),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_50),
.B(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_67),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_60),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_119),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_66),
.Y(n_224)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_66),
.Y(n_325)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

XOR2x1_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_72),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_73),
.A2(n_74),
.B1(n_110),
.B2(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_74),
.B(n_107),
.C(n_110),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_115),
.C(n_116),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_106),
.C(n_113),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_78),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_95),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_96),
.C(n_100),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.C(n_91),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_175)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_83),
.Y(n_338)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_84),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_85),
.Y(n_308)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_91),
.B(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_106),
.B(n_113),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_107),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_110),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_110),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_110),
.B(n_160),
.C(n_168),
.Y(n_192)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21x1_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_293),
.B(n_557),
.Y(n_120)
);

NOR3x1_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_197),
.C(n_287),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_122),
.A2(n_558),
.B(n_561),
.Y(n_557)
);

NOR2xp67_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_123),
.B(n_125),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_189),
.C(n_194),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_126),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_174),
.C(n_176),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_128),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_142),
.C(n_159),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_129),
.B(n_142),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_130),
.B(n_132),
.C(n_137),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_137),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_141),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_149),
.C(n_154),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_143),
.B(n_154),
.Y(n_220)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_147),
.Y(n_448)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_149),
.B(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_153),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_158),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_164),
.Y(n_271)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_168),
.A2(n_169),
.B1(n_179),
.B2(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_179),
.C(n_182),
.Y(n_178)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_172),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_174),
.B(n_176),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_185),
.C(n_187),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_178),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_222),
.C(n_225),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_179),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_179),
.A2(n_225),
.B1(n_233),
.B2(n_241),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_181),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_182),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_182),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_182),
.A2(n_230),
.B1(n_315),
.B2(n_364),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_187),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_185),
.B(n_259),
.C(n_263),
.Y(n_258)
);

XNOR2x2_ASAP7_75t_SL g300 ( 
.A(n_185),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_187),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_187),
.A2(n_216),
.B1(n_217),
.B2(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_189),
.A2(n_194),
.B1(n_195),
.B2(n_291),
.Y(n_290)
);

INVxp33_ASAP7_75t_SL g291 ( 
.A(n_189),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_193),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_190),
.B(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_192),
.B(n_193),
.Y(n_282)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_276),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_198),
.B(n_276),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_234),
.C(n_237),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_199),
.B(n_234),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_218),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_204),
.B(n_278),
.C(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_216),
.C(n_217),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_205),
.B(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.C(n_215),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_206),
.B(n_215),
.Y(n_256)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_216),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.C(n_229),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_219),
.B(n_221),
.Y(n_347)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_228),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_229),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_230),
.B(n_310),
.C(n_315),
.Y(n_309)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_237),
.B(n_387),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_257),
.C(n_272),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_238),
.B(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.C(n_255),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_239),
.B(n_242),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.C(n_250),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_243),
.A2(n_250),
.B1(n_251),
.B2(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_243),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_247),
.B(n_383),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_249),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_250),
.B(n_442),
.C(n_446),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_250),
.A2(n_251),
.B1(n_442),
.B2(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g356 ( 
.A(n_255),
.B(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_257),
.B(n_273),
.Y(n_344)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.C(n_269),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g340 ( 
.A(n_258),
.B(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_263),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_262),
.Y(n_418)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_266),
.B(n_270),
.Y(n_341)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_267),
.Y(n_525)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_269),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_269),
.A2(n_270),
.B1(n_420),
.B2(n_421),
.Y(n_541)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_281),
.C(n_286),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_280)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_288),
.A2(n_559),
.B(n_560),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_292),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_289),
.B(n_292),
.Y(n_560)
);

AO21x2_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_391),
.B(n_554),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_385),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_350),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_296),
.B(n_350),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_342),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_297),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_319),
.C(n_339),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_299),
.B(n_354),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.C(n_309),
.Y(n_299)
);

XNOR2x1_ASAP7_75t_L g426 ( 
.A(n_300),
.B(n_427),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_302),
.A2(n_303),
.B1(n_309),
.B2(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_305),
.B(n_408),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_309),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_314),
.Y(n_466)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_315),
.Y(n_364)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_320),
.A2(n_339),
.B1(n_340),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_330),
.C(n_337),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_321),
.B(n_380),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.C(n_326),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_322),
.B(n_326),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_322),
.B(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_322),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_324),
.B(n_403),
.Y(n_402)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_330),
.A2(n_331),
.B1(n_337),
.B2(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_337),
.Y(n_381)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_345),
.B1(n_348),
.B2(n_349),
.Y(n_342)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_343),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_345),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_389),
.C(n_390),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_356),
.C(n_358),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_352),
.A2(n_353),
.B1(n_356),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_379),
.C(n_382),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_360),
.B(n_400),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_365),
.C(n_370),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XNOR2x1_ASAP7_75t_SL g451 ( 
.A(n_362),
.B(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_365),
.B(n_370),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_369),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_366),
.B(n_369),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_368),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_375),
.C(n_376),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_371),
.A2(n_375),
.B1(n_438),
.B2(n_439),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_371),
.Y(n_438)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_375),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_375),
.B(n_506),
.C(n_508),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_375),
.A2(n_439),
.B1(n_508),
.B2(n_509),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_376),
.B(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_378),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_382),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_385),
.A2(n_555),
.B(n_556),
.Y(n_554)
);

AND2x2_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_386),
.B(n_388),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_453),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_397),
.C(n_429),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_394),
.B(n_398),
.Y(n_455)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_401),
.C(n_426),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_426),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.C(n_409),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_404),
.Y(n_434)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_434),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_419),
.C(n_420),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g540 ( 
.A(n_410),
.B(n_541),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_415),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_411),
.B(n_415),
.Y(n_492)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_411),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_411),
.A2(n_517),
.B1(n_518),
.B2(n_527),
.Y(n_526)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_418),
.Y(n_476)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NOR2x1_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_432),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.C(n_451),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_433),
.B(n_552),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_435),
.B(n_451),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_440),
.C(n_449),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_436),
.B(n_546),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_441),
.B(n_450),
.Y(n_546)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_442),
.Y(n_499)
);

INVx8_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XOR2x2_ASAP7_75t_L g497 ( 
.A(n_446),
.B(n_498),
.Y(n_497)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_455),
.C(n_456),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_457),
.A2(n_549),
.B(n_553),
.Y(n_456)
);

AOI21x1_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_535),
.B(n_548),
.Y(n_457)
);

OAI21x1_ASAP7_75t_SL g458 ( 
.A1(n_459),
.A2(n_500),
.B(n_534),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_488),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_460),
.B(n_488),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_468),
.C(n_477),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_461),
.B(n_503),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_467),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_467),
.C(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_468),
.A2(n_469),
.B1(n_477),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_474),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_470),
.B(n_474),
.Y(n_507)
);

INVx5_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_473),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_477),
.Y(n_504)
);

AO22x1_ASAP7_75t_SL g477 ( 
.A1(n_478),
.A2(n_483),
.B1(n_486),
.B2(n_487),
.Y(n_477)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_478),
.Y(n_486)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_483),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_483),
.B(n_486),
.Y(n_490)
);

INVx6_ASAP7_75t_L g520 ( 
.A(n_484),
.Y(n_520)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_487),
.B(n_529),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_494),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_489),
.B(n_495),
.C(n_497),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

MAJx2_ASAP7_75t_L g543 ( 
.A(n_490),
.B(n_492),
.C(n_493),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_497),
.Y(n_494)
);

AOI21x1_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_511),
.B(n_533),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_505),
.Y(n_501)
);

NOR2x1_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_505),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_506),
.A2(n_507),
.B1(n_514),
.B2(n_515),
.Y(n_513)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_512),
.A2(n_521),
.B(n_532),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_SL g512 ( 
.A(n_513),
.B(n_516),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_513),
.B(n_516),
.Y(n_532)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_518),
.Y(n_527)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_528),
.B(n_531),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_526),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_523),
.B(n_526),
.Y(n_531)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_536),
.B(n_547),
.Y(n_535)
);

NOR2x1p5_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_547),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_538),
.B1(n_544),
.B2(n_545),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_538),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_539),
.A2(n_540),
.B1(n_542),
.B2(n_543),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_539),
.B(n_543),
.C(n_544),
.Y(n_550)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NOR2xp67_ASAP7_75t_SL g549 ( 
.A(n_550),
.B(n_551),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_550),
.B(n_551),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_572),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_564),
.B(n_572),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_566),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_567),
.Y(n_571)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_574),
.Y(n_573)
);


endmodule