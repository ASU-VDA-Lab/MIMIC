module real_jpeg_4580_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_0),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_0),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_0),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_0),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_0),
.B(n_52),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_0),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_0),
.Y(n_151)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_2),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_2),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_2),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_2),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_2),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_2),
.B(n_115),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_2),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_3),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_3),
.B(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_3),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_3),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_3),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_3),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_3),
.B(n_164),
.Y(n_403)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_4),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_4),
.Y(n_255)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_6),
.B(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_6),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_6),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_6),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_6),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_6),
.B(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_6),
.B(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_7),
.Y(n_149)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_7),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_7),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_7),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_7),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_8),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_8),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g377 ( 
.A(n_8),
.Y(n_377)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_11),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_11),
.B(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_11),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_11),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_11),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_11),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_11),
.B(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_11),
.A2(n_372),
.B(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_12),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_12),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_13),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_13),
.B(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_13),
.B(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_13),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_13),
.B(n_226),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_13),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_13),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_13),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_14),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_14),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_14),
.B(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_14),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_14),
.B(n_115),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_15),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_15),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_15),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_15),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_15),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_15),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_15),
.B(n_286),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_15),
.B(n_52),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_452),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_200),
.B(n_450),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_168),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_20),
.B(n_168),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_97),
.C(n_125),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_21),
.B(n_97),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_68),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_22),
.B(n_69),
.C(n_85),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_44),
.C(n_54),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_23),
.B(n_44),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_24),
.B(n_33),
.C(n_38),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_24),
.A2(n_25),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_24),
.B(n_120),
.C(n_124),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_24),
.A2(n_25),
.B1(n_144),
.B2(n_145),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_25),
.B(n_145),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_29),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_29),
.Y(n_356)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_38),
.B2(n_43),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_37),
.Y(n_159)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_37),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_37),
.Y(n_334)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_38),
.A2(n_43),
.B1(n_463),
.B2(n_464),
.Y(n_462)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_42),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.C(n_51),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_45),
.B(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g317 ( 
.A(n_47),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_48),
.B(n_51),
.Y(n_141)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_50),
.Y(n_217)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_54),
.B(n_421),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_60),
.C(n_63),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_55),
.A2(n_66),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_55),
.B(n_381),
.C(n_384),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_57),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_58),
.Y(n_242)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_62),
.A2(n_63),
.B1(n_74),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_62),
.A2(n_63),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_71),
.C(n_74),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_63),
.B(n_235),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_85),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_77),
.C(n_81),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_70),
.B(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_71),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_71),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_71),
.A2(n_128),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_73),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_74),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_74),
.A2(n_131),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_74),
.B(n_337),
.Y(n_365)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_77),
.A2(n_81),
.B1(n_93),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_87),
.B1(n_88),
.B2(n_93),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_84),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_88),
.B(n_93),
.C(n_96),
.Y(n_189)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_92),
.Y(n_361)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_117),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_99),
.B(n_100),
.C(n_117),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_113),
.B2(n_114),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_107),
.B1(n_111),
.B2(n_112),
.Y(n_102)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_105),
.Y(n_220)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_106),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_107),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_111),
.C(n_114),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_107),
.B(n_134),
.Y(n_396)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_133),
.C(n_135),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_124),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_120),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_122),
.A2(n_124),
.B1(n_181),
.B2(n_184),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_122),
.A2(n_124),
.B1(n_325),
.B2(n_329),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_122),
.B(n_325),
.C(n_330),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_124),
.B(n_176),
.C(n_181),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_125),
.B(n_427),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_142),
.C(n_165),
.Y(n_125)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_126),
.B(n_423),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_140),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_127),
.B(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_128),
.B(n_192),
.C(n_196),
.Y(n_461)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_132),
.B(n_140),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_135),
.B(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_L g423 ( 
.A(n_142),
.B(n_165),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_156),
.C(n_160),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_143),
.B(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_150),
.C(n_154),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_144),
.A2(n_145),
.B1(n_154),
.B2(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_149),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_150),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_150),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_150),
.A2(n_175),
.B1(n_176),
.B2(n_412),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_152),
.Y(n_328)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_154),
.Y(n_415)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_155),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_156),
.A2(n_160),
.B1(n_161),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_156),
.Y(n_406)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_159),
.Y(n_294)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_169),
.B(n_171),
.C(n_185),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_185),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_171),
.B(n_459),
.Y(n_458)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.CI(n_174),
.CON(n_171),
.SN(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_175),
.A2(n_176),
.B1(n_358),
.B2(n_362),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_175),
.B(n_351),
.C(n_362),
.Y(n_397)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_181),
.Y(n_184)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_186),
.B(n_188),
.C(n_191),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_194),
.B(n_239),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_196),
.Y(n_199)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_198),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI221xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_389),
.B1(n_443),
.B2(n_448),
.C(n_449),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_344),
.B(n_388),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_305),
.B(n_343),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_280),
.B(n_304),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_247),
.B(n_279),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_236),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_207),
.B(n_236),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_221),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_208),
.B(n_222),
.C(n_233),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_209),
.B(n_214),
.C(n_218),
.Y(n_290)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_233),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_228),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_224),
.B(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.C(n_243),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_238),
.A2(n_243),
.B1(n_244),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_238),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_273),
.B(n_278),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_263),
.B(n_272),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_260),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_260),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_256),
.Y(n_274)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_282),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_289),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_283),
.B(n_290),
.C(n_291),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_288),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_296),
.C(n_303),
.Y(n_339)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_299),
.B2(n_303),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_299),
.Y(n_303)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_342),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_342),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_322),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_311),
.C(n_322),
.Y(n_345)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_311)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_316),
.B2(n_318),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_313),
.B(n_318),
.C(n_319),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_335),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_339),
.C(n_341),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_330),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_325),
.Y(n_329)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_335)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_336),
.Y(n_341)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_345),
.B(n_346),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_368),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_348),
.B(n_349),
.C(n_368),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_363),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_350),
.B(n_364),
.C(n_367),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_357),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_358),
.Y(n_362)
);

INVx6_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_365),
.B1(n_366),
.B2(n_367),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_387),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_378),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_370),
.B(n_378),
.C(n_387),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_372),
.B(n_376),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_402),
.C(n_403),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_417),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_384),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

NOR3xp33_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_425),
.C(n_429),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_390),
.A2(n_444),
.B(n_447),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_418),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_391),
.B(n_418),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_407),
.C(n_409),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_392),
.B(n_407),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_400),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_401),
.C(n_404),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_397),
.C(n_398),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_399),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_403),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.C(n_416),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_416),
.Y(n_433)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_424),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_422),
.C(n_424),
.Y(n_428)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_425),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_428),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_439),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_430),
.A2(n_445),
.B(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_437),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_437),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_434),
.C(n_435),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_434),
.B(n_435),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_440),
.B(n_441),
.Y(n_445)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_472),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_455),
.B(n_456),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_465),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_468),
.A2(n_469),
.B1(n_470),
.B2(n_471),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_468),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_469),
.Y(n_471)
);


endmodule