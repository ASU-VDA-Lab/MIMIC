module fake_jpeg_483_n_652 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_652);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_652;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_67),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_27),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_66),
.B(n_70),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_23),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_68),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_0),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_71),
.B(n_86),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_73),
.Y(n_208)
);

INVx2_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_74),
.B(n_5),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_27),
.B(n_18),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_75),
.B(n_81),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_51),
.Y(n_77)
);

CKINVDCx6p67_ASAP7_75t_R g228 ( 
.A(n_77),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_82),
.B(n_85),
.Y(n_177)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_84),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_18),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_100),
.Y(n_160)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_90),
.B(n_93),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_91),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_32),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_94),
.B(n_35),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_95),
.Y(n_224)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_97),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_0),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_98),
.B(n_101),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_1),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_56),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_103),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_32),
.B(n_2),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_105),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_56),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_106),
.B(n_119),
.Y(n_197)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_21),
.Y(n_112)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_46),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_113),
.B(n_116),
.Y(n_218)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_41),
.B(n_3),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_42),
.B(n_4),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_54),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_122),
.B(n_123),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_42),
.B(n_4),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_54),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_125),
.B(n_63),
.Y(n_221)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_47),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_47),
.Y(n_130)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_70),
.A2(n_22),
.B1(n_26),
.B2(n_30),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_165),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_53),
.B1(n_29),
.B2(n_34),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_77),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_138),
.B(n_144),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_81),
.A2(n_22),
.B1(n_26),
.B2(n_30),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_99),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g155 ( 
.A(n_74),
.B(n_53),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_155),
.B(n_171),
.Y(n_295)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_58),
.A2(n_53),
.B1(n_29),
.B2(n_54),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_159),
.A2(n_204),
.B1(n_215),
.B2(n_222),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_163),
.B(n_91),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_98),
.A2(n_25),
.B1(n_36),
.B2(n_50),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_113),
.A2(n_31),
.B1(n_36),
.B2(n_50),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_166),
.A2(n_174),
.B1(n_202),
.B2(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_97),
.A2(n_35),
.B1(n_114),
.B2(n_104),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_80),
.A2(n_25),
.B1(n_31),
.B2(n_29),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_124),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_180),
.B(n_188),
.Y(n_309)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_96),
.Y(n_184)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_59),
.A2(n_45),
.B1(n_34),
.B2(n_54),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_185),
.A2(n_84),
.B1(n_127),
.B2(n_117),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_126),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_189),
.Y(n_266)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_190),
.Y(n_288)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_192),
.Y(n_291)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_194),
.Y(n_300)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_94),
.A2(n_4),
.B(n_5),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_198),
.A2(n_203),
.B(n_222),
.Y(n_276)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_201),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_60),
.A2(n_62),
.B1(n_72),
.B2(n_115),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_118),
.A2(n_54),
.B(n_45),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_111),
.A2(n_45),
.B1(n_34),
.B2(n_54),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_129),
.A2(n_57),
.B1(n_38),
.B2(n_20),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_73),
.A2(n_57),
.B1(n_38),
.B2(n_20),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_211),
.A2(n_219),
.B1(n_9),
.B2(n_10),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_212),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_64),
.B(n_57),
.C(n_20),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_212),
.C(n_217),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_109),
.A2(n_20),
.B1(n_7),
.B2(n_8),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_76),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_61),
.B(n_6),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_220),
.B(n_225),
.Y(n_232)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_128),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_92),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_61),
.B(n_91),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_228),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_229),
.B(n_230),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_228),
.Y(n_230)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_149),
.Y(n_233)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_233),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_95),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_235),
.B(n_238),
.Y(n_316)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_236),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_87),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_239),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_160),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_241),
.B(n_245),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_242),
.A2(n_275),
.B1(n_296),
.B2(n_305),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_169),
.B(n_79),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_243),
.B(n_249),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_134),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_248),
.B(n_147),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_173),
.B(n_130),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_L g323 ( 
.A(n_251),
.B(n_276),
.C(n_310),
.Y(n_323)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_154),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_253),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_198),
.B(n_9),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_255),
.B(n_260),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_132),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_274),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_143),
.A2(n_110),
.B1(n_78),
.B2(n_69),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_258),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_259),
.A2(n_262),
.B1(n_267),
.B2(n_193),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_11),
.Y(n_260)
);

OA22x2_ASAP7_75t_L g261 ( 
.A1(n_137),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_261)
);

OA22x2_ASAP7_75t_L g360 ( 
.A1(n_261),
.A2(n_233),
.B1(n_239),
.B2(n_301),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_211),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_262)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_263),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_135),
.Y(n_264)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_264),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_145),
.A2(n_15),
.B1(n_16),
.B2(n_156),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_265),
.A2(n_270),
.B1(n_289),
.B2(n_312),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_204),
.A2(n_172),
.B1(n_164),
.B2(n_170),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_161),
.Y(n_268)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_268),
.Y(n_319)
);

INVx4_ASAP7_75t_SL g269 ( 
.A(n_196),
.Y(n_269)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_179),
.A2(n_170),
.B1(n_151),
.B2(n_185),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_159),
.B(n_15),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_271),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_210),
.B(n_148),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_272),
.B(n_290),
.Y(n_335)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_152),
.Y(n_273)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_227),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_177),
.A2(n_191),
.B1(n_168),
.B2(n_183),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_168),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_277),
.B(n_278),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_183),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_131),
.Y(n_279)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_178),
.Y(n_281)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_153),
.A2(n_217),
.B(n_179),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_282),
.A2(n_306),
.B(n_286),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_142),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_283),
.B(n_284),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_151),
.Y(n_284)
);

AND2x4_ASAP7_75t_L g285 ( 
.A(n_159),
.B(n_157),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_285),
.A2(n_286),
.B(n_306),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_200),
.B(n_226),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_286),
.B(n_287),
.C(n_306),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_133),
.B(n_162),
.Y(n_287)
);

INVx11_ASAP7_75t_L g289 ( 
.A(n_193),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_176),
.B(n_182),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_131),
.Y(n_292)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_154),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_302),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_208),
.A2(n_135),
.B1(n_187),
.B2(n_158),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_196),
.B(n_207),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_308),
.Y(n_344)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_186),
.Y(n_298)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_178),
.Y(n_299)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_299),
.Y(n_339)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_207),
.Y(n_301)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_301),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g302 ( 
.A(n_154),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_152),
.Y(n_303)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_303),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_146),
.Y(n_304)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_146),
.A2(n_187),
.B1(n_158),
.B2(n_224),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_205),
.B(n_206),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_208),
.Y(n_307)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_307),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_153),
.B(n_206),
.Y(n_308)
);

AND2x4_ASAP7_75t_SL g310 ( 
.A(n_205),
.B(n_139),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_224),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_269),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_147),
.A2(n_139),
.B1(n_141),
.B2(n_175),
.Y(n_312)
);

AO22x2_ASAP7_75t_SL g313 ( 
.A1(n_271),
.A2(n_215),
.B1(n_150),
.B2(n_175),
.Y(n_313)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_295),
.A2(n_214),
.B1(n_141),
.B2(n_150),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_314),
.A2(n_325),
.B1(n_352),
.B2(n_365),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_320),
.B(n_324),
.C(n_334),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_235),
.B(n_214),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_331),
.A2(n_368),
.B(n_291),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_243),
.B(n_249),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_346),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_293),
.B(n_272),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_351),
.Y(n_377)
);

OAI32xp33_ASAP7_75t_L g349 ( 
.A1(n_285),
.A2(n_238),
.A3(n_271),
.B1(n_255),
.B2(n_246),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_349),
.B(n_360),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_240),
.B(n_232),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_295),
.A2(n_285),
.B1(n_276),
.B2(n_254),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_285),
.A2(n_252),
.B1(n_267),
.B2(n_262),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_353),
.A2(n_372),
.B1(n_325),
.B2(n_364),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_248),
.B(n_251),
.C(n_234),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_247),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g357 ( 
.A(n_231),
.B(n_251),
.CI(n_260),
.CON(n_357),
.SN(n_357)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_357),
.B(n_288),
.Y(n_390)
);

O2A1O1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_254),
.A2(n_310),
.B(n_261),
.C(n_308),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_361),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_309),
.B(n_290),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_297),
.B(n_287),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_373),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_254),
.A2(n_261),
.B1(n_282),
.B2(n_307),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_287),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_371),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_261),
.A2(n_237),
.B1(n_244),
.B2(n_254),
.Y(n_369)
);

OAI22x1_ASAP7_75t_L g383 ( 
.A1(n_369),
.A2(n_303),
.B1(n_273),
.B2(n_292),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_236),
.B(n_250),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_310),
.A2(n_298),
.B1(n_266),
.B2(n_268),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_266),
.B(n_300),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_315),
.Y(n_374)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_374),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_358),
.A2(n_289),
.B1(n_263),
.B2(n_299),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_376),
.A2(n_409),
.B1(n_370),
.B2(n_338),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_379),
.A2(n_381),
.B1(n_383),
.B2(n_384),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_236),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_380),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_353),
.A2(n_304),
.B1(n_264),
.B2(n_281),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_382),
.B(n_354),
.C(n_347),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_317),
.A2(n_280),
.B1(n_257),
.B2(n_300),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_317),
.B(n_288),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_395),
.Y(n_426)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_319),
.Y(n_388)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_388),
.Y(n_425)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_319),
.Y(n_389)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_389),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_390),
.B(n_417),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_345),
.A2(n_291),
.B1(n_250),
.B2(n_279),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_392),
.A2(n_405),
.B1(n_406),
.B2(n_383),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_344),
.B(n_334),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_396),
.Y(n_438)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_397),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_318),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_401),
.Y(n_433)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_399),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_400),
.A2(n_402),
.B(n_415),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_343),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_368),
.A2(n_349),
.B(n_352),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_403),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_316),
.B(n_344),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_407),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_324),
.A2(n_253),
.B1(n_302),
.B2(n_335),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_359),
.A2(n_302),
.B1(n_335),
.B2(n_316),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_361),
.B(n_330),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_330),
.B(n_320),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_413),
.Y(n_435)
);

CKINVDCx6p67_ASAP7_75t_R g409 ( 
.A(n_329),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_363),
.A2(n_323),
.B1(n_331),
.B2(n_355),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_412),
.A2(n_420),
.B1(n_333),
.B2(n_356),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_350),
.B(n_342),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_322),
.B(n_341),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_414),
.B(n_418),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_350),
.A2(n_358),
.B(n_313),
.Y(n_415)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_357),
.B(n_372),
.C(n_360),
.Y(n_416)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_339),
.C(n_333),
.Y(n_430)
);

AOI21xp33_ASAP7_75t_L g417 ( 
.A1(n_357),
.A2(n_337),
.B(n_360),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_326),
.B(n_370),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_321),
.A2(n_313),
.B(n_360),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_419),
.A2(n_327),
.B(n_385),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_313),
.A2(n_367),
.B1(n_362),
.B2(n_315),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_354),
.Y(n_421)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_424),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_428),
.B(n_456),
.C(n_458),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_430),
.B(n_393),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_409),
.Y(n_431)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_431),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_409),
.Y(n_432)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_432),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_402),
.A2(n_419),
.B(n_415),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_434),
.A2(n_440),
.B(n_420),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_394),
.A2(n_347),
.B(n_332),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_409),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_441),
.B(n_444),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_378),
.Y(n_443)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_443),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_384),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_392),
.B(n_339),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_461),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_450),
.A2(n_459),
.B1(n_397),
.B2(n_444),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_451),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_387),
.B(n_362),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_453),
.B(n_391),
.Y(n_479)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_454),
.Y(n_490)
);

AOI21x1_ASAP7_75t_L g455 ( 
.A1(n_400),
.A2(n_328),
.B(n_338),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_455),
.A2(n_460),
.B(n_416),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_393),
.B(n_328),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_386),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_457),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_382),
.B(n_332),
.C(n_367),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_385),
.A2(n_327),
.B1(n_411),
.B2(n_394),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_379),
.A2(n_411),
.B1(n_381),
.B2(n_394),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_462),
.A2(n_391),
.B1(n_395),
.B2(n_407),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_453),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_465),
.A2(n_475),
.B1(n_482),
.B2(n_438),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_467),
.A2(n_470),
.B(n_476),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_434),
.A2(n_375),
.B(n_406),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_471),
.B(n_487),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_398),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_473),
.B(n_492),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_433),
.Y(n_474)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_474),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_433),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_442),
.A2(n_375),
.B(n_412),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_447),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_477),
.B(n_486),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_479),
.B(n_483),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_428),
.C(n_413),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_480),
.B(n_497),
.C(n_423),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_460),
.A2(n_405),
.B(n_404),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_481),
.A2(n_484),
.B(n_491),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_447),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_442),
.A2(n_455),
.B(n_436),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_435),
.B(n_408),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_422),
.Y(n_488)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_440),
.A2(n_401),
.B(n_410),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_439),
.B(n_410),
.Y(n_492)
);

MAJx2_ASAP7_75t_L g493 ( 
.A(n_435),
.B(n_390),
.C(n_377),
.Y(n_493)
);

MAJx2_ASAP7_75t_L g529 ( 
.A(n_493),
.B(n_437),
.C(n_452),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_450),
.A2(n_388),
.B1(n_389),
.B2(n_396),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_494),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_461),
.A2(n_421),
.B(n_399),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_499),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_496),
.A2(n_429),
.B1(n_448),
.B2(n_438),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_458),
.B(n_427),
.C(n_426),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_425),
.Y(n_498)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_498),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_462),
.A2(n_430),
.B(n_457),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_430),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_500),
.B(n_437),
.Y(n_533)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_490),
.Y(n_501)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_501),
.Y(n_541)
);

NOR2x1_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_476),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_505),
.B(n_509),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_479),
.B(n_423),
.Y(n_506)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_506),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_507),
.B(n_533),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_469),
.B(n_426),
.Y(n_508)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_508),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_463),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_466),
.B(n_480),
.C(n_471),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_510),
.B(n_520),
.C(n_524),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_427),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_512),
.B(n_516),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_465),
.B(n_459),
.Y(n_514)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_514),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_466),
.B(n_454),
.Y(n_516)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_518),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_519),
.A2(n_526),
.B1(n_472),
.B2(n_467),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_425),
.C(n_449),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_463),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_521),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_494),
.Y(n_523)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_523),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_449),
.C(n_446),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_481),
.Y(n_525)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_525),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_496),
.A2(n_429),
.B1(n_448),
.B2(n_446),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_490),
.Y(n_528)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_528),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_529),
.B(n_486),
.Y(n_538)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_498),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_495),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_470),
.B(n_452),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_491),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_475),
.B(n_422),
.C(n_445),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_534),
.C(n_507),
.Y(n_547)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_537),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_538),
.B(n_547),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_508),
.B(n_482),
.Y(n_542)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_542),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_544),
.A2(n_560),
.B1(n_517),
.B2(n_511),
.Y(n_575)
);

OA21x2_ASAP7_75t_L g545 ( 
.A1(n_527),
.A2(n_472),
.B(n_499),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_545),
.A2(n_552),
.B(n_515),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_548),
.B(n_555),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_506),
.B(n_489),
.Y(n_549)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_549),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_527),
.A2(n_484),
.B(n_472),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_535),
.B(n_489),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_510),
.B(n_464),
.C(n_485),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_556),
.B(n_564),
.C(n_522),
.Y(n_565)
);

BUFx24_ASAP7_75t_SL g558 ( 
.A(n_503),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_558),
.B(n_441),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_519),
.A2(n_478),
.B1(n_485),
.B2(n_464),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_531),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_561),
.B(n_562),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_514),
.B(n_488),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_516),
.B(n_468),
.C(n_445),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_565),
.B(n_574),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_552),
.A2(n_515),
.B(n_513),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_567),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_546),
.B(n_522),
.C(n_512),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_569),
.B(n_573),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_571),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_546),
.B(n_520),
.C(n_524),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_547),
.B(n_529),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_575),
.A2(n_557),
.B1(n_568),
.B2(n_537),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_556),
.B(n_505),
.C(n_502),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_576),
.B(n_579),
.C(n_587),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_555),
.Y(n_577)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_577),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_553),
.B(n_502),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_578),
.B(n_584),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_553),
.B(n_526),
.C(n_468),
.Y(n_579)
);

INVxp33_ASAP7_75t_L g581 ( 
.A(n_542),
.Y(n_581)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_581),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_583),
.B(n_541),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_540),
.B(n_532),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_536),
.B(n_564),
.Y(n_585)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_585),
.Y(n_595)
);

A2O1A1O1Ixp25_ASAP7_75t_L g586 ( 
.A1(n_538),
.A2(n_501),
.B(n_528),
.C(n_530),
.D(n_432),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_586),
.A2(n_563),
.B(n_545),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_540),
.B(n_431),
.C(n_488),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_591),
.B(n_593),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_576),
.A2(n_545),
.B(n_551),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_565),
.B(n_551),
.C(n_548),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_598),
.B(n_602),
.C(n_603),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_599),
.B(n_543),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_601),
.A2(n_539),
.B1(n_586),
.B2(n_554),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_573),
.B(n_559),
.C(n_560),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_569),
.B(n_544),
.C(n_550),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_584),
.Y(n_604)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_604),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_579),
.B(n_550),
.C(n_562),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_605),
.B(n_587),
.C(n_594),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_582),
.Y(n_606)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_606),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_598),
.B(n_578),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_607),
.B(n_608),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_595),
.A2(n_570),
.B1(n_581),
.B2(n_580),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_610),
.B(n_614),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_589),
.B(n_577),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_611),
.B(n_588),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_597),
.B(n_572),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_612),
.B(n_621),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_589),
.A2(n_575),
.B1(n_543),
.B2(n_554),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_613),
.A2(n_616),
.B(n_592),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_574),
.C(n_566),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_615),
.B(n_619),
.C(n_600),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_600),
.A2(n_571),
.B(n_567),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_603),
.B(n_566),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_617),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_590),
.B(n_539),
.C(n_549),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_609),
.B(n_605),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_623),
.B(n_627),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_622),
.A2(n_616),
.B(n_609),
.Y(n_628)
);

AOI21xp33_ASAP7_75t_L g639 ( 
.A1(n_628),
.A2(n_629),
.B(n_632),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_620),
.B(n_602),
.Y(n_631)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_631),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_610),
.B(n_596),
.C(n_604),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_633),
.B(n_607),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_625),
.B(n_619),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_634),
.B(n_641),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_630),
.A2(n_622),
.B(n_618),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_635),
.A2(n_637),
.B(n_626),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_625),
.A2(n_601),
.B(n_615),
.C(n_478),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g643 ( 
.A(n_640),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_627),
.B(n_617),
.C(n_612),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_636),
.B(n_633),
.C(n_624),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_642),
.B(n_645),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_638),
.B(n_626),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_641),
.C(n_637),
.Y(n_647)
);

A2O1A1O1Ixp25_ASAP7_75t_L g649 ( 
.A1(n_647),
.A2(n_643),
.B(n_644),
.C(n_639),
.D(n_504),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_649),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_650),
.B(n_648),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_651),
.B(n_504),
.Y(n_652)
);


endmodule