module fake_netlist_6_3987_n_612 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_612);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_612;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_167;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_599;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_420;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_311;
wire n_403;
wire n_253;
wire n_583;
wire n_596;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_32),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_10),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_6),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_17),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_27),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_74),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_42),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_29),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_106),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_2),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_40),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_49),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_104),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_54),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_48),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_18),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_60),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_82),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_38),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_51),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_13),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_0),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_14),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_0),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_35),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_53),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_15),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_92),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_63),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_45),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_66),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_98),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_120),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_80),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_30),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_9),
.Y(n_178)
);

BUFx8_ASAP7_75t_SL g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_37),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_1),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_69),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_3),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_26),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_28),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_93),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_109),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_2),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_47),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_65),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_58),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_56),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_19),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_133),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_176),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_169),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_145),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_150),
.B(n_3),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_151),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_164),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_179),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_181),
.Y(n_221)
);

BUFx2_ASAP7_75t_SL g222 ( 
.A(n_153),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g223 ( 
.A(n_159),
.B(n_4),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_134),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_135),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_139),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_136),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_163),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_L g234 ( 
.A(n_159),
.B(n_4),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_189),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_140),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_141),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_142),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_SL g243 ( 
.A(n_197),
.B(n_194),
.Y(n_243)
);

XNOR2x1_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_5),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_198),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_191),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_143),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_199),
.B(n_144),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_227),
.B(n_147),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_R g268 ( 
.A(n_201),
.B(n_5),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_224),
.B(n_149),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_152),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_222),
.B(n_155),
.Y(n_281)
);

NAND2x1_ASAP7_75t_L g282 ( 
.A(n_209),
.B(n_156),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_233),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_233),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_204),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

AND2x6_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_11),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_275),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_242),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

NAND3xp33_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_173),
.C(n_193),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_250),
.B(n_219),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_261),
.B(n_219),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_190),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_258),
.B(n_157),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_258),
.B(n_158),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_272),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_246),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_165),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

AND2x6_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_12),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_268),
.A2(n_188),
.B1(n_186),
.B2(n_185),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_167),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_249),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_268),
.A2(n_175),
.B1(n_174),
.B2(n_172),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_269),
.B(n_168),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_261),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_255),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_254),
.Y(n_321)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

OR2x2_ASAP7_75t_SL g323 ( 
.A(n_287),
.B(n_271),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_264),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_281),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_271),
.B(n_171),
.Y(n_326)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_288),
.B(n_6),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_255),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_263),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_16),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_269),
.B(n_7),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_256),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_273),
.B(n_20),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_245),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_273),
.B(n_21),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_245),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_247),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_247),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_257),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_283),
.B(n_285),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_262),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_265),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_267),
.B(n_22),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_260),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_270),
.Y(n_346)
);

NAND3xp33_ASAP7_75t_L g347 ( 
.A(n_277),
.B(n_8),
.C(n_9),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_243),
.B(n_23),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_243),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_286),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_291),
.Y(n_352)
);

AO22x2_ASAP7_75t_L g353 ( 
.A1(n_347),
.A2(n_244),
.B1(n_286),
.B2(n_284),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_309),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_341),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_283),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_312),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_302),
.B(n_24),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_299),
.B(n_25),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_319),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

AO22x2_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_8),
.B1(n_10),
.B2(n_285),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_292),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_297),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_340),
.Y(n_367)
);

BUFx8_ASAP7_75t_L g368 ( 
.A(n_298),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_320),
.B(n_31),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_304),
.Y(n_370)
);

AO22x2_ASAP7_75t_L g371 ( 
.A1(n_348),
.A2(n_285),
.B1(n_283),
.B2(n_274),
.Y(n_371)
);

NAND2x1p5_ASAP7_75t_L g372 ( 
.A(n_305),
.B(n_283),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_325),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_317),
.B(n_285),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_345),
.Y(n_375)
);

OA22x2_ASAP7_75t_L g376 ( 
.A1(n_313),
.A2(n_316),
.B1(n_346),
.B2(n_348),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_251),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_337),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_320),
.B(n_33),
.Y(n_380)
);

AO22x2_ASAP7_75t_L g381 ( 
.A1(n_300),
.A2(n_34),
.B1(n_36),
.B2(n_39),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_349),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_310),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_296),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_301),
.Y(n_386)
);

OR2x6_ASAP7_75t_L g387 ( 
.A(n_308),
.B(n_41),
.Y(n_387)
);

OA22x2_ASAP7_75t_L g388 ( 
.A1(n_313),
.A2(n_131),
.B1(n_44),
.B2(n_46),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_328),
.B(n_43),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_50),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_305),
.B(n_52),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_301),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_329),
.Y(n_398)
);

BUFx8_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_329),
.B(n_55),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_336),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_L g402 ( 
.A(n_330),
.B(n_289),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_336),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_338),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_339),
.B(n_57),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_322),
.B(n_307),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_350),
.B(n_322),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_386),
.B(n_322),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_397),
.B(n_332),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_373),
.B(n_332),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_360),
.B(n_374),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_407),
.B(n_332),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_407),
.B(n_339),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_354),
.B(n_306),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_351),
.B(n_321),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_SL g417 ( 
.A(n_355),
.B(n_314),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_382),
.B(n_321),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_392),
.B(n_316),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_SL g420 ( 
.A(n_375),
.B(n_331),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_356),
.B(n_295),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_372),
.B(n_327),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_376),
.B(n_344),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_SL g424 ( 
.A(n_377),
.B(n_333),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_357),
.B(n_296),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_361),
.B(n_303),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_363),
.B(n_335),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_366),
.B(n_303),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_358),
.B(n_294),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_294),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g431 ( 
.A(n_359),
.B(n_323),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_400),
.B(n_293),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_400),
.B(n_293),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_367),
.B(n_330),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_379),
.B(n_330),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_389),
.B(n_311),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_394),
.B(n_311),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_387),
.B(n_311),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_390),
.B(n_311),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_395),
.B(n_289),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_387),
.B(n_289),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_385),
.B(n_289),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_385),
.B(n_59),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_383),
.B(n_61),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_370),
.B(n_62),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_384),
.B(n_64),
.Y(n_446)
);

NAND2xp33_ASAP7_75t_SL g447 ( 
.A(n_365),
.B(n_393),
.Y(n_447)
);

AOI31xp67_ASAP7_75t_L g448 ( 
.A1(n_423),
.A2(n_406),
.A3(n_380),
.B(n_369),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_416),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_437),
.A2(n_402),
.B(n_391),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_396),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_435),
.A2(n_430),
.B(n_440),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_419),
.A2(n_388),
.B(n_352),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_436),
.A2(n_352),
.B(n_364),
.Y(n_454)
);

OAI21xp33_ASAP7_75t_L g455 ( 
.A1(n_412),
.A2(n_353),
.B(n_362),
.Y(n_455)
);

AOI31xp67_ASAP7_75t_L g456 ( 
.A1(n_429),
.A2(n_427),
.A3(n_434),
.B(n_439),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_431),
.A2(n_405),
.B(n_404),
.C(n_403),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_438),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_422),
.B(n_401),
.Y(n_459)
);

A2O1A1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_424),
.A2(n_398),
.B(n_378),
.C(n_364),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

AOI21x1_ASAP7_75t_SL g462 ( 
.A1(n_445),
.A2(n_381),
.B(n_362),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_421),
.B(n_353),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_411),
.B(n_410),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_442),
.A2(n_381),
.B(n_371),
.Y(n_465)
);

A2O1A1Ixp33_ASAP7_75t_L g466 ( 
.A1(n_420),
.A2(n_371),
.B(n_368),
.C(n_399),
.Y(n_466)
);

O2A1O1Ixp5_ASAP7_75t_L g467 ( 
.A1(n_408),
.A2(n_368),
.B(n_68),
.C(n_70),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_428),
.A2(n_67),
.B(n_71),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_445),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_432),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_413),
.B(n_399),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_409),
.B(n_128),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_72),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_447),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_458),
.Y(n_476)
);

OR2x6_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_441),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_458),
.Y(n_478)
);

INVx3_ASAP7_75t_SL g479 ( 
.A(n_475),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_418),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_463),
.A2(n_417),
.B1(n_441),
.B2(n_443),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_450),
.A2(n_452),
.B(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_470),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_458),
.Y(n_484)
);

AO21x2_ASAP7_75t_L g485 ( 
.A1(n_460),
.A2(n_457),
.B(n_453),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_474),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_459),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_455),
.A2(n_446),
.B1(n_444),
.B2(n_425),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_473),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_451),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_454),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_469),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_461),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_468),
.A2(n_414),
.B(n_75),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_464),
.B(n_73),
.Y(n_495)
);

AO32x2_ASAP7_75t_L g496 ( 
.A1(n_462),
.A2(n_77),
.A3(n_78),
.B1(n_81),
.B2(n_83),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_465),
.A2(n_474),
.B(n_467),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_472),
.A2(n_456),
.B(n_448),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_466),
.Y(n_499)
);

OAI22xp33_ASAP7_75t_L g500 ( 
.A1(n_475),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_498),
.A2(n_87),
.B(n_88),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_493),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_89),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_476),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_491),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_496),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_476),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_477),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_483),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_496),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_482),
.A2(n_90),
.B(n_94),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_496),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_487),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_487),
.A2(n_96),
.B(n_97),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_479),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_489),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_495),
.A2(n_99),
.B(n_101),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_482),
.A2(n_102),
.B(n_103),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_486),
.B(n_105),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_477),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_492),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_485),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_485),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_497),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_495),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_494),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_486),
.B(n_107),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_476),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_513),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_502),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_R g531 ( 
.A(n_515),
.B(n_499),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_R g532 ( 
.A(n_515),
.B(n_478),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_508),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_R g534 ( 
.A(n_528),
.B(n_484),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_520),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_R g536 ( 
.A(n_528),
.B(n_504),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_502),
.B(n_477),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_519),
.B(n_480),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_R g539 ( 
.A(n_519),
.B(n_108),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_525),
.B(n_481),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_521),
.B(n_481),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_R g542 ( 
.A(n_519),
.B(n_112),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_R g543 ( 
.A(n_528),
.B(n_488),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_504),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_R g545 ( 
.A(n_519),
.B(n_113),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_514),
.B(n_500),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_509),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_114),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_526),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_R g550 ( 
.A(n_527),
.B(n_525),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_509),
.B(n_117),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_529),
.B(n_523),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_547),
.B(n_516),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_540),
.B(n_516),
.Y(n_554)
);

AOI222xp33_ASAP7_75t_L g555 ( 
.A1(n_548),
.A2(n_517),
.B1(n_512),
.B2(n_506),
.C1(n_510),
.C2(n_521),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_530),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_537),
.B(n_505),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_541),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_535),
.B(n_505),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_543),
.B(n_522),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_549),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_544),
.B(n_507),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_549),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_546),
.A2(n_510),
.B1(n_512),
.B2(n_506),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_538),
.B(n_518),
.Y(n_565)
);

NAND2x1_ASAP7_75t_SL g566 ( 
.A(n_550),
.B(n_523),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_553),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_558),
.B(n_565),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_556),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_559),
.B(n_538),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_557),
.B(n_522),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_561),
.B(n_549),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_563),
.B(n_532),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_553),
.B(n_562),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_568),
.B(n_564),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_572),
.B(n_567),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_569),
.B(n_564),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_574),
.B(n_552),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_567),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_569),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_570),
.B(n_560),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_578),
.B(n_571),
.Y(n_582)
);

AO221x2_ASAP7_75t_L g583 ( 
.A1(n_577),
.A2(n_566),
.B1(n_573),
.B2(n_554),
.C(n_542),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_581),
.A2(n_545),
.B1(n_539),
.B2(n_546),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_580),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_577),
.B(n_555),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_585),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_586),
.B(n_575),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_582),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_583),
.B(n_576),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_584),
.B(n_579),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_590),
.B(n_576),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_587),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_589),
.B(n_579),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_592),
.A2(n_588),
.B1(n_591),
.B2(n_531),
.Y(n_595)
);

INVxp67_ASAP7_75t_SL g596 ( 
.A(n_592),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_596),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_597),
.B(n_595),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_597),
.B1(n_593),
.B2(n_594),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_599),
.A2(n_507),
.B1(n_551),
.B2(n_524),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_600),
.B(n_555),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_601),
.B(n_534),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_602),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_603),
.Y(n_604)
);

AOI31xp33_ASAP7_75t_L g605 ( 
.A1(n_604),
.A2(n_536),
.A3(n_119),
.B(n_121),
.Y(n_605)
);

OAI322xp33_ASAP7_75t_L g606 ( 
.A1(n_605),
.A2(n_524),
.A3(n_518),
.B1(n_526),
.B2(n_124),
.C1(n_125),
.C2(n_126),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_606),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_606),
.A2(n_518),
.B1(n_511),
.B2(n_501),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_607),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_608),
.Y(n_610)
);

AOI221xp5_ASAP7_75t_L g611 ( 
.A1(n_609),
.A2(n_526),
.B1(n_122),
.B2(n_123),
.C(n_118),
.Y(n_611)
);

AOI211xp5_ASAP7_75t_L g612 ( 
.A1(n_611),
.A2(n_610),
.B(n_511),
.C(n_501),
.Y(n_612)
);


endmodule