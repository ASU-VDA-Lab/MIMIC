module fake_jpeg_30894_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_10),
.B(n_15),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_44),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

CKINVDCx10_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_47),
.Y(n_108)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_20),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_52),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_28),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_34),
.B1(n_38),
.B2(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_2),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_60),
.Y(n_92)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_19),
.B(n_4),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_24),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_34),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_25),
.C(n_20),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_71),
.B(n_102),
.C(n_106),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_100),
.B1(n_105),
.B2(n_69),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_34),
.B1(n_25),
.B2(n_31),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_80),
.A2(n_81),
.B1(n_101),
.B2(n_110),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_38),
.B1(n_40),
.B2(n_36),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_84),
.B(n_85),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_29),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_24),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_88),
.B(n_89),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_113),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_44),
.B(n_22),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_53),
.A2(n_37),
.B1(n_33),
.B2(n_27),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_45),
.A2(n_62),
.B1(n_61),
.B2(n_55),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_57),
.B(n_4),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_62),
.A2(n_26),
.B1(n_31),
.B2(n_29),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_43),
.B(n_26),
.C(n_27),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_60),
.B(n_36),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_109),
.Y(n_132)
);

CKINVDCx12_ASAP7_75t_R g109 ( 
.A(n_47),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_49),
.A2(n_40),
.B1(n_32),
.B2(n_33),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_35),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_77),
.A2(n_92),
.B(n_90),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_114),
.A2(n_6),
.B(n_11),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_32),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_117),
.B(n_134),
.Y(n_171)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

OR2x2_ASAP7_75t_SL g119 ( 
.A(n_73),
.B(n_68),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_122),
.A2(n_145),
.B1(n_79),
.B2(n_111),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_76),
.A2(n_59),
.B1(n_65),
.B2(n_63),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_58),
.B1(n_52),
.B2(n_33),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_133),
.B1(n_144),
.B2(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_126),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_129),
.Y(n_157)
);

AND2x4_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_35),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_130),
.B(n_152),
.Y(n_179)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_80),
.A2(n_48),
.B1(n_46),
.B2(n_35),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_86),
.A2(n_35),
.B(n_37),
.C(n_33),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_135),
.B(n_139),
.Y(n_187)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_141),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_73),
.B(n_71),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_35),
.B1(n_68),
.B2(n_37),
.Y(n_144)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_73),
.B(n_37),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_78),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_99),
.A2(n_37),
.B1(n_33),
.B2(n_8),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_70),
.B1(n_99),
.B2(n_82),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_5),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_169),
.B1(n_172),
.B2(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_70),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_161),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_160),
.A2(n_168),
.B1(n_186),
.B2(n_170),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_104),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_93),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_112),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_164),
.A2(n_185),
.B(n_116),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_111),
.B1(n_79),
.B2(n_97),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_170),
.B1(n_184),
.B2(n_186),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_103),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_177),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_74),
.B1(n_103),
.B2(n_10),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_74),
.B1(n_9),
.B2(n_10),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_133),
.B1(n_114),
.B2(n_151),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_144),
.B(n_129),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_6),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_119),
.B(n_11),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_144),
.C(n_139),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_121),
.B(n_12),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_13),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_133),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_13),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_133),
.A2(n_14),
.B1(n_135),
.B2(n_144),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_164),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_193),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_215),
.B1(n_180),
.B2(n_155),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_145),
.B1(n_131),
.B2(n_129),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_126),
.B1(n_118),
.B2(n_120),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_209),
.B1(n_160),
.B2(n_158),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_200),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_115),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_203),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_128),
.Y(n_203)
);

INVx6_ASAP7_75t_SL g204 ( 
.A(n_158),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_207),
.Y(n_222)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_132),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_210),
.Y(n_225)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_140),
.B(n_138),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_159),
.B(n_14),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_153),
.B(n_137),
.C(n_125),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_217),
.C(n_179),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_153),
.B(n_125),
.C(n_127),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_220),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_127),
.B1(n_142),
.B2(n_161),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_221),
.B1(n_154),
.B2(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_162),
.A2(n_142),
.B1(n_167),
.B2(n_163),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_227),
.B1(n_240),
.B2(n_211),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_235),
.C(n_238),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_229),
.A2(n_224),
.B(n_246),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_179),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_243),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_179),
.C(n_174),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_174),
.C(n_155),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_209),
.A2(n_180),
.B1(n_157),
.B2(n_175),
.Y(n_240)
);

AO22x2_ASAP7_75t_L g242 ( 
.A1(n_210),
.A2(n_157),
.B1(n_183),
.B2(n_185),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_244),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_190),
.B(n_157),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_192),
.A2(n_196),
.B1(n_207),
.B2(n_189),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_196),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_246),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_191),
.B(n_221),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_239),
.B(n_214),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_250),
.B(n_254),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_216),
.C(n_217),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_256),
.C(n_257),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_241),
.B1(n_247),
.B2(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_214),
.C(n_219),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_194),
.C(n_198),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_225),
.A2(n_189),
.B(n_220),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_262),
.B(n_243),
.C(n_242),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_218),
.C(n_212),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_266),
.C(n_242),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_208),
.C(n_204),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_SL g271 ( 
.A(n_261),
.B(n_242),
.C(n_240),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_222),
.A2(n_201),
.B(n_205),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_238),
.C(n_244),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_233),
.Y(n_267)
);

BUFx12_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_241),
.B1(n_247),
.B2(n_228),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_282),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_272),
.Y(n_291)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_245),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_269),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_223),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_248),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_278),
.C(n_259),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_242),
.C(n_236),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_279),
.A2(n_262),
.B1(n_249),
.B2(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_263),
.B(n_254),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_270),
.B(n_275),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_293),
.C(n_295),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_291),
.B1(n_286),
.B2(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_296),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_256),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_260),
.B1(n_249),
.B2(n_268),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_279),
.B1(n_278),
.B2(n_277),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_275),
.Y(n_301)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_292),
.B(n_295),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_307),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_289),
.A2(n_264),
.B(n_275),
.C(n_284),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_306),
.Y(n_308)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_269),
.C(n_273),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_314),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_312),
.A2(n_305),
.B(n_304),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_237),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_237),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_311),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_306),
.B1(n_303),
.B2(n_307),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_303),
.Y(n_318)
);

OAI31xp33_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_312),
.A3(n_310),
.B(n_313),
.Y(n_321)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_319),
.B1(n_316),
.B2(n_290),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_323),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_325),
.Y(n_327)
);


endmodule