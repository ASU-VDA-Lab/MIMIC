module fake_netlist_5_2099_n_1597 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1597);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1597;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1557;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1564;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_5),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_88),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_109),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_86),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_108),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_61),
.Y(n_229)
);

BUFx8_ASAP7_75t_SL g230 ( 
.A(n_218),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_79),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_78),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_92),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_162),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_110),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_166),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_100),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_48),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_199),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_205),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_50),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_202),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_94),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_154),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_96),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_27),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_47),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_98),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_11),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_123),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_24),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_49),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_135),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_213),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_23),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_12),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_143),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_25),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_129),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_145),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_105),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_128),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_215),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_203),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_81),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_32),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_117),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_210),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_54),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_82),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_18),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_171),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_142),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_7),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_45),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_194),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_34),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_17),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_197),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_159),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_103),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_138),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_49),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_30),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_2),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_90),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_74),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_42),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_43),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_93),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_17),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_57),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_42),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_70),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_214),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_36),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_190),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_55),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_191),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_95),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_67),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_102),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_137),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_198),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_31),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_31),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_68),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_161),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_58),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_1),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_19),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_66),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_134),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_207),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_112),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_156),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_173),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_26),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_53),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_118),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_139),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_24),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_119),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_160),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_83),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_133),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_106),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_56),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_155),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_5),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_7),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_158),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_172),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_87),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_39),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_91),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_37),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_8),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_209),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_99),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_192),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_188),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_12),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_113),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_15),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_32),
.Y(n_352)
);

BUFx8_ASAP7_75t_SL g353 ( 
.A(n_126),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_183),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_8),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_111),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_174),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_148),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_36),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_45),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_141),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_73),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_167),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_115),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_279),
.B(n_51),
.Y(n_365)
);

BUFx8_ASAP7_75t_SL g366 ( 
.A(n_249),
.Y(n_366)
);

BUFx8_ASAP7_75t_SL g367 ( 
.A(n_249),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_279),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_250),
.A2(n_0),
.B(n_1),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_254),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_256),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_273),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_263),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_283),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_221),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_310),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_257),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_260),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_273),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_289),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_297),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_317),
.Y(n_383)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_273),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_355),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_240),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_240),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_273),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_337),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_341),
.A2(n_4),
.B(n_6),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_349),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_285),
.B(n_52),
.Y(n_396)
);

BUFx8_ASAP7_75t_L g397 ( 
.A(n_233),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_351),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_257),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_345),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_288),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_257),
.B(n_9),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_259),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_285),
.B(n_10),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_345),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_252),
.B(n_13),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_252),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_280),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_308),
.B(n_14),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_288),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_306),
.A2(n_16),
.B(n_18),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_222),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_226),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_284),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_227),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_306),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_290),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_291),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_315),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_325),
.B(n_16),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_294),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_239),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_315),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_308),
.B(n_19),
.Y(n_430)
);

BUFx12f_ASAP7_75t_L g431 ( 
.A(n_295),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_330),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_331),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_331),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_332),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_235),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_332),
.B(n_59),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_292),
.B(n_20),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_342),
.B(n_60),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_277),
.A2(n_359),
.B1(n_302),
.B2(n_311),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_237),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_299),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_241),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_342),
.B(n_20),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_244),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_262),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_267),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_271),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_312),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_316),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_276),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_425),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_R g454 ( 
.A(n_423),
.B(n_236),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_366),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_425),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_425),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_423),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_443),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_366),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_443),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_410),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_296),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_425),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_R g466 ( 
.A(n_431),
.B(n_236),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_425),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_367),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_378),
.B(n_243),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_373),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_373),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_429),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_367),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_420),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_431),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_420),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_397),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_429),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_397),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_397),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_429),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_429),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_376),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_378),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_428),
.B(n_419),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_401),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_401),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_424),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_429),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_424),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_R g492 ( 
.A(n_450),
.B(n_239),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_450),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_428),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_427),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_404),
.B(n_293),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_451),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_409),
.B(n_275),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_433),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_433),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_433),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_389),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_390),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_433),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_433),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_368),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_368),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_377),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_377),
.B(n_298),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_441),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_411),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_411),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_436),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_436),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_R g516 ( 
.A(n_370),
.B(n_243),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_370),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_383),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_370),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_R g520 ( 
.A(n_447),
.B(n_251),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_R g521 ( 
.A(n_447),
.B(n_251),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_365),
.Y(n_522)
);

INVxp33_ASAP7_75t_L g523 ( 
.A(n_412),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_498),
.B(n_486),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_517),
.B(n_519),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_453),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_517),
.B(n_414),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_396),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_494),
.B(n_430),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_406),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_508),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_457),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_458),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_516),
.B(n_396),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_484),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_522),
.B(n_396),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

INVxp33_ASAP7_75t_L g539 ( 
.A(n_454),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_470),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_522),
.B(n_365),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_470),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_510),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_463),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_459),
.B(n_460),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_467),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_464),
.B(n_365),
.Y(n_548)
);

AO221x1_ASAP7_75t_L g549 ( 
.A1(n_501),
.A2(n_379),
.B1(n_387),
.B2(n_447),
.C(n_436),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_472),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_512),
.B(n_513),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_479),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_512),
.B(n_438),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_509),
.B(n_439),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_482),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_520),
.B(n_438),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_483),
.B(n_438),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_485),
.B(n_417),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_513),
.B(n_445),
.C(n_421),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_490),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_487),
.B(n_418),
.Y(n_561)
);

NOR3xp33_ASAP7_75t_L g562 ( 
.A(n_504),
.B(n_413),
.C(n_408),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_463),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_499),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_488),
.B(n_437),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_521),
.B(n_440),
.Y(n_566)
);

NOR3xp33_ASAP7_75t_L g567 ( 
.A(n_469),
.B(n_321),
.C(n_343),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_474),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_523),
.B(n_452),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_470),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_511),
.B(n_442),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_492),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_500),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_502),
.B(n_440),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_505),
.B(n_440),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_474),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_518),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_511),
.B(n_444),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_477),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_506),
.B(n_514),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_515),
.B(n_404),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_477),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_496),
.B(n_404),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_503),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_495),
.A2(n_309),
.B1(n_329),
.B2(n_269),
.Y(n_585)
);

BUFx6f_ASAP7_75t_SL g586 ( 
.A(n_476),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_476),
.B(n_452),
.Y(n_587)
);

OAI21xp33_ASAP7_75t_L g588 ( 
.A1(n_497),
.A2(n_382),
.B(n_372),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_544),
.B(n_489),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_544),
.B(n_403),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_587),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_549),
.A2(n_524),
.B1(n_393),
.B2(n_369),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_541),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_525),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_525),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_569),
.B(n_374),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_538),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_569),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_530),
.B(n_483),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_557),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_557),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_557),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_582),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_571),
.Y(n_604)
);

AND3x2_ASAP7_75t_SL g605 ( 
.A(n_549),
.B(n_281),
.C(n_272),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_538),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_532),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_528),
.B(n_436),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_541),
.Y(n_609)
);

AND2x2_ASAP7_75t_SL g610 ( 
.A(n_567),
.B(n_416),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_582),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_556),
.A2(n_269),
.B1(n_329),
.B2(n_309),
.Y(n_612)
);

NOR2x2_ASAP7_75t_L g613 ( 
.A(n_585),
.B(n_484),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_532),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_536),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_551),
.B(n_476),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_556),
.B(n_436),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_548),
.B(n_493),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_545),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_529),
.B(n_491),
.Y(n_620)
);

BUFx12f_ASAP7_75t_L g621 ( 
.A(n_584),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_587),
.B(n_459),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_574),
.A2(n_400),
.B(n_384),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_566),
.B(n_535),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_SL g625 ( 
.A(n_539),
.B(n_535),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_584),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_542),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_446),
.Y(n_628)
);

NOR2x1p5_ASAP7_75t_L g629 ( 
.A(n_526),
.B(n_478),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_545),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_572),
.B(n_460),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_536),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_578),
.B(n_462),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_537),
.B(n_446),
.Y(n_634)
);

NAND3xp33_ASAP7_75t_SL g635 ( 
.A(n_531),
.B(n_462),
.C(n_358),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_563),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_558),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_553),
.B(n_340),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_554),
.B(n_446),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_563),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_561),
.B(n_446),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_559),
.A2(n_340),
.B1(n_362),
.B2(n_358),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_568),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_577),
.B(n_466),
.Y(n_644)
);

NOR2x2_ASAP7_75t_L g645 ( 
.A(n_562),
.B(n_272),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_527),
.B(n_374),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_541),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_577),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_575),
.A2(n_393),
.B1(n_369),
.B2(n_416),
.Y(n_649)
);

OR2x6_ASAP7_75t_L g650 ( 
.A(n_546),
.B(n_371),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_539),
.B(n_475),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_568),
.A2(n_393),
.B1(n_369),
.B2(n_416),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_565),
.B(n_533),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_R g654 ( 
.A(n_586),
.B(n_468),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_534),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_540),
.B(n_375),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_576),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_586),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_547),
.B(n_550),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_586),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_576),
.A2(n_434),
.B1(n_435),
.B2(n_415),
.Y(n_661)
);

BUFx12f_ASAP7_75t_SL g662 ( 
.A(n_588),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_552),
.B(n_446),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_579),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_555),
.B(n_473),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_581),
.A2(n_400),
.B(n_384),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_560),
.A2(n_362),
.B1(n_268),
.B2(n_224),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_579),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_564),
.B(n_448),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_573),
.A2(n_339),
.B1(n_225),
.B2(n_228),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_570),
.B(n_301),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_583),
.A2(n_346),
.B1(n_229),
.B2(n_231),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_541),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_580),
.A2(n_415),
.B1(n_434),
.B2(n_435),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_570),
.Y(n_675)
);

OAI21xp33_ASAP7_75t_SL g676 ( 
.A1(n_624),
.A2(n_305),
.B(n_303),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_SL g677 ( 
.A1(n_616),
.A2(n_570),
.B(n_350),
.C(n_318),
.Y(n_677)
);

AO21x1_ASAP7_75t_L g678 ( 
.A1(n_625),
.A2(n_334),
.B(n_449),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_606),
.Y(n_679)
);

BUFx12f_ASAP7_75t_L g680 ( 
.A(n_621),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_600),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_617),
.A2(n_543),
.B(n_541),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_610),
.A2(n_448),
.B1(n_344),
.B2(n_281),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_593),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_604),
.B(n_480),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_604),
.B(n_543),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_606),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_601),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_633),
.B(n_481),
.Y(n_689)
);

AO32x2_ASAP7_75t_L g690 ( 
.A1(n_612),
.A2(n_398),
.A3(n_371),
.B1(n_543),
.B2(n_344),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_SL g691 ( 
.A1(n_633),
.A2(n_461),
.B1(n_456),
.B2(n_360),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_598),
.B(n_385),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_634),
.A2(n_400),
.B(n_384),
.Y(n_693)
);

AO21x2_ASAP7_75t_L g694 ( 
.A1(n_628),
.A2(n_392),
.B(n_385),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_638),
.A2(n_335),
.B(n_232),
.C(n_234),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_637),
.B(n_456),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_616),
.B(n_461),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_639),
.B(n_223),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_627),
.B(n_238),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_608),
.A2(n_400),
.B(n_384),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_638),
.A2(n_347),
.B1(n_242),
.B2(n_247),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_594),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_615),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_622),
.B(n_230),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_SL g705 ( 
.A1(n_599),
.A2(n_412),
.B(n_392),
.C(n_395),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_652),
.A2(n_400),
.B(n_384),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_593),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_602),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_610),
.A2(n_448),
.B1(n_422),
.B2(n_405),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_626),
.B(n_245),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_591),
.B(n_230),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_592),
.A2(n_338),
.B1(n_248),
.B2(n_253),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_591),
.B(n_246),
.Y(n_713)
);

AOI222xp33_ASAP7_75t_L g714 ( 
.A1(n_635),
.A2(n_395),
.B1(n_398),
.B2(n_386),
.C1(n_388),
.C2(n_381),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_641),
.B(n_255),
.Y(n_715)
);

BUFx8_ASAP7_75t_L g716 ( 
.A(n_632),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_648),
.B(n_375),
.Y(n_717)
);

NAND2x1p5_ASAP7_75t_L g718 ( 
.A(n_607),
.B(n_470),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_593),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_631),
.B(n_353),
.Y(n_720)
);

AND2x6_ASAP7_75t_L g721 ( 
.A(n_590),
.B(n_381),
.Y(n_721)
);

AOI21xp33_ASAP7_75t_L g722 ( 
.A1(n_620),
.A2(n_261),
.B(n_258),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_SL g723 ( 
.A(n_593),
.B(n_609),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_596),
.B(n_264),
.Y(n_724)
);

NAND2x1p5_ASAP7_75t_L g725 ( 
.A(n_596),
.B(n_471),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_648),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_609),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_603),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_SL g729 ( 
.A(n_642),
.B(n_266),
.C(n_265),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_635),
.B(n_353),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_652),
.A2(n_649),
.B(n_647),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_649),
.A2(n_471),
.B(n_380),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_609),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_620),
.B(n_618),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_630),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_590),
.B(n_386),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_650),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_614),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_595),
.Y(n_739)
);

CKINVDCx8_ASAP7_75t_R g740 ( 
.A(n_650),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_653),
.A2(n_618),
.B(n_592),
.C(n_589),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_597),
.A2(n_422),
.B(n_405),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_644),
.B(n_388),
.Y(n_743)
);

O2A1O1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_653),
.A2(n_405),
.B(n_422),
.C(n_432),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_609),
.A2(n_471),
.B(n_380),
.Y(n_745)
);

AOI21x1_ASAP7_75t_L g746 ( 
.A1(n_623),
.A2(n_669),
.B(n_663),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_667),
.A2(n_333),
.B1(n_274),
.B2(n_278),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_647),
.A2(n_471),
.B(n_373),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_589),
.Y(n_749)
);

BUFx12f_ASAP7_75t_L g750 ( 
.A(n_650),
.Y(n_750)
);

O2A1O1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_611),
.A2(n_432),
.B(n_322),
.C(n_364),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_662),
.B(n_270),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_651),
.B(n_282),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_659),
.A2(n_354),
.B(n_287),
.C(n_300),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_SL g755 ( 
.A(n_658),
.B(n_286),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_655),
.A2(n_643),
.B(n_640),
.C(n_657),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_646),
.Y(n_757)
);

BUFx12f_ASAP7_75t_L g758 ( 
.A(n_629),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_665),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_670),
.B(n_304),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_646),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_672),
.B(n_307),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_675),
.A2(n_647),
.B1(n_673),
.B2(n_668),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_647),
.A2(n_373),
.B(n_380),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_656),
.B(n_313),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_673),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_673),
.A2(n_636),
.B(n_619),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_664),
.A2(n_432),
.B(n_348),
.C(n_363),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_656),
.A2(n_327),
.B(n_361),
.C(n_357),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_673),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_666),
.A2(n_314),
.B(n_319),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_671),
.A2(n_320),
.B1(n_323),
.B2(n_356),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_671),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_681),
.B(n_658),
.Y(n_774)
);

AO21x2_ASAP7_75t_L g775 ( 
.A1(n_678),
.A2(n_605),
.B(n_660),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_738),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_680),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_735),
.Y(n_778)
);

OAI21x1_ASAP7_75t_L g779 ( 
.A1(n_746),
.A2(n_661),
.B(n_674),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_688),
.B(n_660),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_726),
.Y(n_781)
);

BUFx2_ASAP7_75t_R g782 ( 
.A(n_740),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_716),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_703),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_743),
.B(n_674),
.Y(n_785)
);

OAI21x1_ASAP7_75t_L g786 ( 
.A1(n_731),
.A2(n_661),
.B(n_671),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_684),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_716),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_735),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_728),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_702),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_708),
.Y(n_792)
);

BUFx4_ASAP7_75t_SL g793 ( 
.A(n_757),
.Y(n_793)
);

AOI22x1_ASAP7_75t_L g794 ( 
.A1(n_732),
.A2(n_605),
.B1(n_448),
.B2(n_645),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_684),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_684),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_707),
.Y(n_797)
);

AOI22x1_ASAP7_75t_L g798 ( 
.A1(n_767),
.A2(n_739),
.B1(n_708),
.B2(n_679),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_761),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_707),
.Y(n_800)
);

OA21x2_ASAP7_75t_L g801 ( 
.A1(n_742),
.A2(n_671),
.B(n_448),
.Y(n_801)
);

INVx8_ASAP7_75t_L g802 ( 
.A(n_721),
.Y(n_802)
);

OAI21x1_ASAP7_75t_L g803 ( 
.A1(n_682),
.A2(n_671),
.B(n_140),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_687),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_734),
.B(n_654),
.Y(n_805)
);

INVx8_ASAP7_75t_L g806 ( 
.A(n_721),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_750),
.Y(n_807)
);

AO21x1_ASAP7_75t_L g808 ( 
.A1(n_741),
.A2(n_21),
.B(n_22),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_758),
.Y(n_809)
);

OAI21x1_ASAP7_75t_SL g810 ( 
.A1(n_756),
.A2(n_136),
.B(n_220),
.Y(n_810)
);

OAI21x1_ASAP7_75t_L g811 ( 
.A1(n_763),
.A2(n_132),
.B(n_193),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_770),
.Y(n_812)
);

BUFx2_ASAP7_75t_R g813 ( 
.A(n_710),
.Y(n_813)
);

BUFx12f_ASAP7_75t_L g814 ( 
.A(n_737),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_694),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_717),
.B(n_654),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_707),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_721),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_736),
.B(n_749),
.Y(n_819)
);

INVx6_ASAP7_75t_L g820 ( 
.A(n_719),
.Y(n_820)
);

AO21x2_ASAP7_75t_L g821 ( 
.A1(n_694),
.A2(n_613),
.B(n_407),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_766),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_723),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_719),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_759),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_686),
.B(n_21),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_752),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_766),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_L g829 ( 
.A(n_721),
.B(n_373),
.Y(n_829)
);

OR2x6_ASAP7_75t_L g830 ( 
.A(n_773),
.B(n_380),
.Y(n_830)
);

AO21x2_ASAP7_75t_L g831 ( 
.A1(n_698),
.A2(n_402),
.B(n_399),
.Y(n_831)
);

OAI21x1_ASAP7_75t_L g832 ( 
.A1(n_706),
.A2(n_748),
.B(n_745),
.Y(n_832)
);

CKINVDCx14_ASAP7_75t_R g833 ( 
.A(n_691),
.Y(n_833)
);

CKINVDCx14_ASAP7_75t_R g834 ( 
.A(n_696),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_719),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_727),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_727),
.Y(n_837)
);

CKINVDCx6p67_ASAP7_75t_R g838 ( 
.A(n_736),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_765),
.Y(n_839)
);

BUFx12f_ASAP7_75t_L g840 ( 
.A(n_692),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_718),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_692),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_727),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_733),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_733),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_733),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_725),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_773),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_690),
.B(n_62),
.Y(n_849)
);

OAI21x1_ASAP7_75t_L g850 ( 
.A1(n_700),
.A2(n_131),
.B(n_219),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_753),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_689),
.B(n_22),
.Y(n_852)
);

AO21x2_ASAP7_75t_L g853 ( 
.A1(n_715),
.A2(n_677),
.B(n_695),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_724),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_764),
.A2(n_130),
.B(n_216),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_713),
.Y(n_856)
);

BUFx8_ASAP7_75t_SL g857 ( 
.A(n_699),
.Y(n_857)
);

OA21x2_ASAP7_75t_L g858 ( 
.A1(n_709),
.A2(n_407),
.B(n_402),
.Y(n_858)
);

BUFx12f_ASAP7_75t_L g859 ( 
.A(n_755),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_754),
.A2(n_127),
.B(n_189),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_711),
.Y(n_861)
);

BUFx12f_ASAP7_75t_L g862 ( 
.A(n_714),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_744),
.A2(n_693),
.B(n_768),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_704),
.Y(n_864)
);

NAND2x1p5_ASAP7_75t_L g865 ( 
.A(n_772),
.B(n_407),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_690),
.B(n_63),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_697),
.Y(n_867)
);

BUFx12f_ASAP7_75t_L g868 ( 
.A(n_685),
.Y(n_868)
);

CKINVDCx16_ASAP7_75t_R g869 ( 
.A(n_729),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_789),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_781),
.Y(n_871)
);

BUFx8_ASAP7_75t_SL g872 ( 
.A(n_783),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_778),
.Y(n_873)
);

OAI22xp33_ASAP7_75t_L g874 ( 
.A1(n_862),
.A2(n_730),
.B1(n_720),
.B2(n_760),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_778),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_817),
.Y(n_876)
);

AO21x2_ASAP7_75t_L g877 ( 
.A1(n_815),
.A2(n_705),
.B(n_771),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_789),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_784),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_785),
.B(n_690),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_790),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_784),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_840),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_785),
.B(n_683),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_790),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_848),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_848),
.Y(n_887)
);

BUFx8_ASAP7_75t_L g888 ( 
.A(n_788),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_825),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_792),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_792),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_862),
.A2(n_762),
.B1(n_701),
.B2(n_747),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_791),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_852),
.A2(n_722),
.B1(n_712),
.B2(n_676),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_856),
.B(n_769),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_776),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_791),
.Y(n_897)
);

OAI21xp33_ASAP7_75t_L g898 ( 
.A1(n_842),
.A2(n_751),
.B(n_407),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_822),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_819),
.B(n_849),
.Y(n_900)
);

INVx4_ASAP7_75t_L g901 ( 
.A(n_817),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_794),
.A2(n_407),
.B1(n_402),
.B2(n_399),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_826),
.A2(n_786),
.B(n_779),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_812),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_782),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_819),
.B(n_64),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_812),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_832),
.A2(n_147),
.B(n_212),
.Y(n_908)
);

CKINVDCx11_ASAP7_75t_R g909 ( 
.A(n_783),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_822),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_815),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_798),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_804),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_804),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_798),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_828),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_840),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_859),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_854),
.B(n_23),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_779),
.Y(n_920)
);

OA21x2_ASAP7_75t_L g921 ( 
.A1(n_808),
.A2(n_811),
.B(n_803),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_799),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_819),
.B(n_65),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_828),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_794),
.A2(n_402),
.B1(n_399),
.B2(n_394),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_837),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_832),
.A2(n_149),
.B(n_211),
.Y(n_927)
);

AO21x1_ASAP7_75t_L g928 ( 
.A1(n_849),
.A2(n_866),
.B(n_860),
.Y(n_928)
);

NAND2x1p5_ASAP7_75t_L g929 ( 
.A(n_848),
.B(n_380),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_837),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_866),
.B(n_69),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_859),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_805),
.A2(n_402),
.B1(n_399),
.B2(n_394),
.Y(n_933)
);

INVx4_ASAP7_75t_SL g934 ( 
.A(n_848),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_845),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_848),
.B(n_818),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_851),
.A2(n_399),
.B1(n_394),
.B2(n_391),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_845),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_816),
.B(n_71),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_801),
.Y(n_940)
);

CKINVDCx11_ASAP7_75t_R g941 ( 
.A(n_788),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_801),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_SL g943 ( 
.A1(n_867),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_801),
.Y(n_944)
);

BUFx12f_ASAP7_75t_L g945 ( 
.A(n_777),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_786),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_858),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_827),
.B(n_28),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_858),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_836),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_817),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_858),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_803),
.A2(n_150),
.B(n_208),
.Y(n_953)
);

INVx6_ASAP7_75t_L g954 ( 
.A(n_795),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_777),
.Y(n_955)
);

AO21x2_ASAP7_75t_L g956 ( 
.A1(n_808),
.A2(n_125),
.B(n_206),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_816),
.B(n_72),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_836),
.Y(n_958)
);

INVx6_ASAP7_75t_L g959 ( 
.A(n_795),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_820),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_851),
.B(n_75),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_869),
.A2(n_394),
.B1(n_391),
.B2(n_30),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_823),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_774),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_818),
.A2(n_394),
.B1(n_391),
.B2(n_33),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_775),
.B(n_151),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_865),
.A2(n_124),
.B(n_201),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_774),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_839),
.A2(n_391),
.B1(n_29),
.B2(n_33),
.Y(n_969)
);

INVx5_ASAP7_75t_L g970 ( 
.A(n_802),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_774),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_867),
.B(n_28),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_780),
.B(n_29),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_780),
.Y(n_974)
);

OAI21x1_ASAP7_75t_SL g975 ( 
.A1(n_810),
.A2(n_153),
.B(n_200),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_858),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_780),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_821),
.A2(n_391),
.B1(n_35),
.B2(n_37),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_787),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_873),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_900),
.B(n_821),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_889),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_876),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_SL g984 ( 
.A1(n_892),
.A2(n_833),
.B(n_834),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_884),
.A2(n_861),
.B1(n_868),
.B2(n_864),
.Y(n_985)
);

CKINVDCx6p67_ASAP7_75t_R g986 ( 
.A(n_945),
.Y(n_986)
);

OR2x6_ASAP7_75t_L g987 ( 
.A(n_936),
.B(n_802),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_936),
.B(n_802),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_881),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_900),
.B(n_821),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_884),
.B(n_775),
.Y(n_991)
);

NOR3xp33_ASAP7_75t_SL g992 ( 
.A(n_874),
.B(n_932),
.C(n_918),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_895),
.A2(n_868),
.B1(n_864),
.B2(n_861),
.Y(n_993)
);

CKINVDCx16_ASAP7_75t_R g994 ( 
.A(n_945),
.Y(n_994)
);

XOR2x2_ASAP7_75t_SL g995 ( 
.A(n_943),
.B(n_969),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_879),
.B(n_775),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_964),
.B(n_838),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_878),
.B(n_853),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_873),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_878),
.B(n_853),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_928),
.A2(n_857),
.B1(n_814),
.B2(n_838),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_880),
.B(n_875),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_885),
.Y(n_1003)
);

CKINVDCx11_ASAP7_75t_R g1004 ( 
.A(n_955),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_904),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_907),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_SL g1007 ( 
.A1(n_962),
.A2(n_865),
.B(n_813),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_968),
.B(n_841),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_879),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_971),
.B(n_841),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_928),
.A2(n_814),
.B1(n_810),
.B2(n_853),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_R g1012 ( 
.A(n_918),
.B(n_787),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_974),
.B(n_847),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_870),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_882),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_R g1016 ( 
.A(n_932),
.B(n_787),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_872),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_872),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_R g1019 ( 
.A(n_909),
.B(n_809),
.Y(n_1019)
);

BUFx10_ASAP7_75t_L g1020 ( 
.A(n_961),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_894),
.A2(n_829),
.B(n_811),
.C(n_802),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_936),
.B(n_806),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_977),
.B(n_847),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_906),
.B(n_807),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_934),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_931),
.A2(n_830),
.B1(n_865),
.B2(n_806),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_909),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_939),
.B(n_796),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_893),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_R g1030 ( 
.A(n_882),
.B(n_809),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_897),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_939),
.B(n_796),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_875),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_913),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_890),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_914),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_871),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_957),
.B(n_796),
.Y(n_1038)
);

CKINVDCx16_ASAP7_75t_R g1039 ( 
.A(n_955),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_931),
.A2(n_830),
.B1(n_806),
.B2(n_843),
.Y(n_1040)
);

AO31x2_ASAP7_75t_L g1041 ( 
.A1(n_912),
.A2(n_795),
.A3(n_824),
.B(n_831),
.Y(n_1041)
);

BUFx4f_ASAP7_75t_SL g1042 ( 
.A(n_888),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_L g1043 ( 
.A(n_963),
.B(n_824),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_890),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_896),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_916),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_908),
.A2(n_863),
.B(n_850),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_924),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_957),
.B(n_797),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_899),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_922),
.B(n_797),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_941),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_899),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_966),
.A2(n_807),
.B1(n_806),
.B2(n_829),
.Y(n_1054)
);

AND2x4_ASAP7_75t_SL g1055 ( 
.A(n_961),
.B(n_824),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_891),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_910),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_973),
.B(n_797),
.Y(n_1058)
);

CKINVDCx16_ASAP7_75t_R g1059 ( 
.A(n_917),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_880),
.B(n_891),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_908),
.A2(n_863),
.B(n_850),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_972),
.A2(n_830),
.B1(n_846),
.B2(n_817),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_910),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_966),
.A2(n_844),
.B1(n_800),
.B2(n_820),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_911),
.B(n_800),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_950),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_958),
.Y(n_1067)
);

AO22x2_ASAP7_75t_L g1068 ( 
.A1(n_920),
.A2(n_844),
.B1(n_800),
.B2(n_793),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_926),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_923),
.B(n_844),
.Y(n_1070)
);

OAI21xp33_ASAP7_75t_L g1071 ( 
.A1(n_919),
.A2(n_855),
.B(n_830),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_876),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_998),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_1068),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_991),
.B(n_946),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_991),
.B(n_920),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_1068),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_998),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_996),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1000),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_1066),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1002),
.B(n_911),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1000),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_985),
.A2(n_948),
.B1(n_956),
.B2(n_978),
.Y(n_1084)
);

OAI31xp33_ASAP7_75t_L g1085 ( 
.A1(n_1007),
.A2(n_898),
.A3(n_965),
.B(n_961),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_981),
.B(n_946),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1002),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1047),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_987),
.B(n_903),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1061),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1014),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_990),
.B(n_956),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1060),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1060),
.B(n_956),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_987),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_989),
.B(n_906),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_987),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_988),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_1011),
.B(n_921),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_988),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1003),
.B(n_921),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1005),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1006),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1046),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_1009),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1048),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_988),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1029),
.B(n_906),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1031),
.B(n_921),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1034),
.B(n_947),
.Y(n_1110)
);

AND2x2_ASAP7_75t_SL g1111 ( 
.A(n_1001),
.B(n_1025),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1022),
.B(n_927),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1036),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_985),
.B(n_912),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_980),
.B(n_930),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1069),
.B(n_947),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1041),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1050),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1053),
.B(n_949),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_1041),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1041),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1022),
.B(n_927),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1067),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1057),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1063),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_999),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1033),
.B(n_949),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_1022),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1035),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1044),
.B(n_952),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1056),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_1037),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1065),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1065),
.B(n_952),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1058),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_983),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_983),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_1015),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1111),
.B(n_993),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_1123),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1106),
.Y(n_1141)
);

AND2x4_ASAP7_75t_SL g1142 ( 
.A(n_1123),
.B(n_1020),
.Y(n_1142)
);

NOR3xp33_ASAP7_75t_SL g1143 ( 
.A(n_1085),
.B(n_1016),
.C(n_1012),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1106),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_SL g1145 ( 
.A(n_1074),
.Y(n_1145)
);

OAI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_1084),
.A2(n_1007),
.B(n_984),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1092),
.B(n_1028),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1092),
.B(n_1032),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1092),
.B(n_1086),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_1079),
.B(n_1076),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1135),
.B(n_1045),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1086),
.B(n_1038),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1079),
.B(n_1062),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1079),
.B(n_1062),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1091),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1085),
.A2(n_967),
.B1(n_1024),
.B2(n_975),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1086),
.B(n_1049),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1091),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1091),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1075),
.B(n_1079),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_SL g1161 ( 
.A1(n_1084),
.A2(n_984),
.B(n_1054),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1106),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1075),
.B(n_1071),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1112),
.B(n_1021),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_1107),
.B(n_1025),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1075),
.B(n_1101),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1135),
.B(n_1045),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1113),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1111),
.B(n_992),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1091),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1076),
.B(n_982),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1102),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1135),
.B(n_1051),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1101),
.B(n_1070),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1138),
.B(n_905),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1113),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1112),
.B(n_953),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1101),
.B(n_877),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1076),
.B(n_915),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1080),
.B(n_915),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1112),
.B(n_1122),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1132),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1109),
.B(n_877),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1135),
.B(n_1024),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1113),
.Y(n_1185)
);

AND2x2_ASAP7_75t_SL g1186 ( 
.A(n_1107),
.B(n_1055),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1132),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1109),
.B(n_877),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1102),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1102),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1143),
.A2(n_1111),
.B1(n_1077),
.B2(n_1074),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1141),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1149),
.B(n_1109),
.Y(n_1193)
);

AOI31xp33_ASAP7_75t_L g1194 ( 
.A1(n_1169),
.A2(n_1027),
.A3(n_1052),
.B(n_1017),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1149),
.B(n_1094),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1181),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1141),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_L g1198 ( 
.A(n_1146),
.B(n_1030),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1155),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1151),
.B(n_1081),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1167),
.B(n_1081),
.Y(n_1201)
);

AND2x4_ASAP7_75t_SL g1202 ( 
.A(n_1182),
.B(n_1107),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1166),
.B(n_1094),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1181),
.B(n_1074),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1144),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1155),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1166),
.B(n_1094),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1187),
.B(n_1105),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1144),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1150),
.B(n_1080),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1173),
.B(n_1105),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1160),
.B(n_1080),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1160),
.B(n_1080),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_L g1214 ( 
.A(n_1171),
.B(n_1138),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1162),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1147),
.B(n_1083),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1150),
.B(n_1083),
.Y(n_1217)
);

NOR2xp67_ASAP7_75t_L g1218 ( 
.A(n_1171),
.B(n_1107),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1140),
.B(n_1083),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1140),
.B(n_1147),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1148),
.B(n_1181),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1148),
.B(n_1083),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1181),
.B(n_1099),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1162),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1163),
.B(n_1089),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1163),
.B(n_1089),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1184),
.B(n_1087),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1168),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1158),
.B(n_1099),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1174),
.B(n_1089),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1152),
.B(n_1087),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1158),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1168),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1174),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1152),
.B(n_1093),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1178),
.B(n_1089),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1176),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1178),
.B(n_1089),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1176),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1177),
.B(n_1074),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1175),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1185),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1157),
.B(n_1093),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1159),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1183),
.B(n_1089),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1157),
.B(n_1093),
.Y(n_1246)
);

AOI32xp33_ASAP7_75t_L g1247 ( 
.A1(n_1198),
.A2(n_1146),
.A3(n_1191),
.B1(n_1139),
.B2(n_1214),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1211),
.B(n_1179),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1220),
.B(n_1153),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1205),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1205),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1241),
.A2(n_1161),
.B1(n_1145),
.B2(n_1156),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1200),
.B(n_1179),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1241),
.A2(n_1111),
.B1(n_1077),
.B2(n_1186),
.Y(n_1254)
);

INVx5_ASAP7_75t_L g1255 ( 
.A(n_1196),
.Y(n_1255)
);

INVxp67_ASAP7_75t_SL g1256 ( 
.A(n_1229),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1209),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1199),
.Y(n_1258)
);

XNOR2xp5_ASAP7_75t_L g1259 ( 
.A(n_1204),
.B(n_1018),
.Y(n_1259)
);

OAI32xp33_ASAP7_75t_L g1260 ( 
.A1(n_1223),
.A2(n_1077),
.A3(n_1201),
.B1(n_1220),
.B2(n_1208),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1221),
.B(n_1164),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1199),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1206),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_R g1264 ( 
.A(n_1196),
.B(n_1019),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1218),
.B(n_1186),
.Y(n_1265)
);

NOR2x1_ASAP7_75t_L g1266 ( 
.A(n_1198),
.B(n_1185),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1227),
.B(n_1102),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1206),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1221),
.B(n_1164),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1232),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1223),
.B(n_1153),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1209),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1215),
.Y(n_1273)
);

NAND2xp33_ASAP7_75t_R g1274 ( 
.A(n_1219),
.B(n_1240),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1215),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1231),
.B(n_1235),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1228),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1240),
.B(n_1164),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1210),
.B(n_1154),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1247),
.A2(n_1077),
.B1(n_1154),
.B2(n_1186),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1250),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1266),
.A2(n_1240),
.B(n_1164),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1252),
.A2(n_1264),
.B1(n_1254),
.B2(n_1274),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1265),
.A2(n_1108),
.B(n_1096),
.Y(n_1284)
);

OAI221xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1259),
.A2(n_995),
.B1(n_1099),
.B2(n_1114),
.C(n_986),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1251),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1257),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1261),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1264),
.A2(n_1204),
.B1(n_1107),
.B2(n_1098),
.Y(n_1289)
);

INVxp33_ASAP7_75t_L g1290 ( 
.A(n_1253),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1269),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1272),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1265),
.A2(n_1100),
.B1(n_1095),
.B2(n_1128),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1273),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1255),
.Y(n_1295)
);

XOR2x2_ASAP7_75t_L g1296 ( 
.A(n_1248),
.B(n_1194),
.Y(n_1296)
);

INVxp67_ASAP7_75t_SL g1297 ( 
.A(n_1258),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1278),
.A2(n_1204),
.B1(n_1098),
.B2(n_1100),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1271),
.A2(n_1096),
.B1(n_1108),
.B2(n_1128),
.Y(n_1299)
);

AOI211x1_ASAP7_75t_L g1300 ( 
.A1(n_1260),
.A2(n_1246),
.B(n_1243),
.C(n_1225),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1275),
.Y(n_1301)
);

AOI211xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1278),
.A2(n_1042),
.B(n_1177),
.C(n_1114),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1278),
.A2(n_1097),
.B1(n_1100),
.B2(n_1095),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1277),
.Y(n_1304)
);

OAI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1274),
.A2(n_1100),
.B1(n_1128),
.B2(n_1095),
.Y(n_1305)
);

XOR2xp5_ASAP7_75t_L g1306 ( 
.A(n_1249),
.B(n_994),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1258),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1279),
.Y(n_1308)
);

XNOR2x1_ASAP7_75t_SL g1309 ( 
.A(n_1255),
.B(n_1004),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1262),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1255),
.B(n_1202),
.Y(n_1311)
);

NAND2xp33_ASAP7_75t_L g1312 ( 
.A(n_1280),
.B(n_1255),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1283),
.B(n_1276),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1283),
.A2(n_975),
.B(n_917),
.C(n_883),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1293),
.A2(n_1267),
.B(n_1256),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1311),
.B(n_1095),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1281),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1296),
.A2(n_1256),
.B(n_1226),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1287),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1306),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1289),
.A2(n_1098),
.B1(n_1177),
.B2(n_1097),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1305),
.A2(n_1177),
.B1(n_1097),
.B2(n_1128),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1309),
.Y(n_1323)
);

AO22x1_ASAP7_75t_L g1324 ( 
.A1(n_1309),
.A2(n_888),
.B1(n_1234),
.B2(n_1263),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1288),
.B(n_1203),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1295),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1292),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1294),
.Y(n_1328)
);

NOR2x1_ASAP7_75t_L g1329 ( 
.A(n_1311),
.B(n_1262),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1286),
.Y(n_1330)
);

NAND3xp33_ASAP7_75t_L g1331 ( 
.A(n_1285),
.B(n_1114),
.C(n_1229),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1291),
.B(n_1203),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1300),
.B(n_1284),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1290),
.B(n_1207),
.Y(n_1334)
);

NOR3xp33_ASAP7_75t_SL g1335 ( 
.A(n_1285),
.B(n_1039),
.C(n_1059),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1308),
.A2(n_1282),
.B1(n_1305),
.B2(n_1303),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1298),
.A2(n_1097),
.B1(n_1226),
.B2(n_1225),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1299),
.A2(n_1165),
.B1(n_1202),
.B2(n_1230),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1299),
.A2(n_1301),
.B1(n_1304),
.B2(n_1230),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1302),
.B(n_1207),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1297),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1297),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1307),
.B(n_1195),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1310),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1281),
.Y(n_1345)
);

NOR3x1_ASAP7_75t_L g1346 ( 
.A(n_1323),
.B(n_883),
.C(n_941),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1330),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1316),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1323),
.A2(n_1165),
.B1(n_1142),
.B2(n_1219),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1333),
.B(n_1195),
.Y(n_1350)
);

AOI211xp5_ASAP7_75t_L g1351 ( 
.A1(n_1318),
.A2(n_1026),
.B(n_1040),
.C(n_1122),
.Y(n_1351)
);

AOI221xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1313),
.A2(n_1224),
.B1(n_1237),
.B2(n_1197),
.C(n_1233),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1331),
.A2(n_1268),
.B(n_1263),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1326),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_1329),
.Y(n_1355)
);

NOR3x1_ASAP7_75t_L g1356 ( 
.A(n_1324),
.B(n_888),
.C(n_1192),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1320),
.B(n_1334),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1317),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1312),
.A2(n_1142),
.B1(n_1245),
.B2(n_1236),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1327),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1339),
.B(n_1193),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1340),
.B(n_1319),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_SL g1363 ( 
.A(n_1335),
.B(n_1165),
.C(n_1210),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_SL g1364 ( 
.A(n_1335),
.B(n_1217),
.C(n_1236),
.Y(n_1364)
);

AOI211xp5_ASAP7_75t_L g1365 ( 
.A1(n_1314),
.A2(n_1026),
.B(n_1040),
.C(n_1122),
.Y(n_1365)
);

NOR3xp33_ASAP7_75t_L g1366 ( 
.A(n_1314),
.B(n_997),
.C(n_1043),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1319),
.B(n_1268),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1316),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1315),
.B(n_1104),
.C(n_1103),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1328),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1336),
.A2(n_1270),
.B(n_1239),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1344),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1338),
.A2(n_1270),
.B(n_1239),
.Y(n_1373)
);

AOI21xp33_ASAP7_75t_L g1374 ( 
.A1(n_1341),
.A2(n_1342),
.B(n_1345),
.Y(n_1374)
);

XOR2x2_ASAP7_75t_L g1375 ( 
.A(n_1337),
.B(n_34),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1343),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1344),
.B(n_1193),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1355),
.A2(n_1322),
.B(n_1321),
.Y(n_1378)
);

OAI21xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1374),
.A2(n_1332),
.B(n_1325),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_SL g1380 ( 
.A1(n_1362),
.A2(n_1228),
.B(n_1242),
.C(n_1217),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1347),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1346),
.B(n_1216),
.Y(n_1382)
);

NAND4xp75_ASAP7_75t_L g1383 ( 
.A(n_1356),
.B(n_923),
.C(n_1245),
.D(n_1238),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1357),
.A2(n_970),
.B1(n_1064),
.B2(n_1122),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1354),
.B(n_1216),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1358),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1359),
.B(n_1222),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1350),
.B(n_1222),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1375),
.B(n_1238),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1364),
.B(n_35),
.Y(n_1390)
);

OAI211xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1374),
.A2(n_1242),
.B(n_1124),
.C(n_1118),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1360),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1363),
.A2(n_1112),
.B(n_1122),
.C(n_1213),
.Y(n_1393)
);

OA22x2_ASAP7_75t_L g1394 ( 
.A1(n_1353),
.A2(n_1370),
.B1(n_1372),
.B2(n_1348),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1367),
.Y(n_1395)
);

NOR3xp33_ASAP7_75t_L g1396 ( 
.A(n_1366),
.B(n_1008),
.C(n_1010),
.Y(n_1396)
);

NOR3xp33_ASAP7_75t_SL g1397 ( 
.A(n_1349),
.B(n_1115),
.C(n_1118),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1376),
.A2(n_1122),
.B1(n_1112),
.B2(n_1183),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1371),
.A2(n_1103),
.B(n_1104),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1369),
.B(n_38),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1352),
.B(n_1212),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1351),
.A2(n_1112),
.B1(n_1188),
.B2(n_1103),
.Y(n_1402)
);

NOR3x1_ASAP7_75t_L g1403 ( 
.A(n_1349),
.B(n_960),
.C(n_1115),
.Y(n_1403)
);

AO22x1_ASAP7_75t_L g1404 ( 
.A1(n_1368),
.A2(n_970),
.B1(n_1104),
.B2(n_1103),
.Y(n_1404)
);

AOI211xp5_ASAP7_75t_L g1405 ( 
.A1(n_1373),
.A2(n_1124),
.B(n_1104),
.C(n_1136),
.Y(n_1405)
);

OAI221xp5_ASAP7_75t_L g1406 ( 
.A1(n_1361),
.A2(n_1244),
.B1(n_1232),
.B2(n_1189),
.C(n_1190),
.Y(n_1406)
);

NOR3xp33_ASAP7_75t_L g1407 ( 
.A(n_1367),
.B(n_1137),
.C(n_1136),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1377),
.B(n_1212),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1377),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1365),
.B(n_1213),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1381),
.Y(n_1411)
);

AOI222xp33_ASAP7_75t_L g1412 ( 
.A1(n_1390),
.A2(n_1189),
.B1(n_1190),
.B2(n_40),
.C1(n_41),
.C2(n_43),
.Y(n_1412)
);

NOR2x1_ASAP7_75t_L g1413 ( 
.A(n_1400),
.B(n_901),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1394),
.A2(n_1244),
.B(n_1082),
.Y(n_1414)
);

AOI221xp5_ASAP7_75t_L g1415 ( 
.A1(n_1395),
.A2(n_1073),
.B1(n_1078),
.B2(n_1023),
.C(n_1013),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1410),
.B(n_38),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1386),
.A2(n_1023),
.B(n_1013),
.C(n_1136),
.Y(n_1417)
);

AOI322xp5_ASAP7_75t_L g1418 ( 
.A1(n_1389),
.A2(n_1188),
.A3(n_902),
.B1(n_925),
.B2(n_1073),
.C1(n_1078),
.C2(n_1159),
.Y(n_1418)
);

AOI221xp5_ASAP7_75t_L g1419 ( 
.A1(n_1392),
.A2(n_1078),
.B1(n_1073),
.B2(n_1170),
.C(n_1172),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1382),
.B(n_39),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1409),
.Y(n_1421)
);

NAND3xp33_ASAP7_75t_L g1422 ( 
.A(n_1397),
.B(n_1137),
.C(n_1136),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1388),
.B(n_40),
.Y(n_1423)
);

OAI211xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1379),
.A2(n_1137),
.B(n_1126),
.C(n_1129),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1393),
.B(n_1170),
.Y(n_1425)
);

OAI211xp5_ASAP7_75t_L g1426 ( 
.A1(n_1402),
.A2(n_1137),
.B(n_44),
.C(n_46),
.Y(n_1426)
);

NOR4xp25_ASAP7_75t_L g1427 ( 
.A(n_1380),
.B(n_41),
.C(n_44),
.D(n_46),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1378),
.A2(n_953),
.B(n_855),
.C(n_1172),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1396),
.A2(n_1405),
.B(n_1401),
.C(n_1391),
.Y(n_1429)
);

NAND4xp25_ASAP7_75t_L g1430 ( 
.A(n_1403),
.B(n_47),
.C(n_48),
.D(n_937),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1385),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1394),
.Y(n_1432)
);

AOI211xp5_ASAP7_75t_L g1433 ( 
.A1(n_1384),
.A2(n_1126),
.B(n_1131),
.C(n_1129),
.Y(n_1433)
);

NAND5xp2_ASAP7_75t_L g1434 ( 
.A(n_1407),
.B(n_1131),
.C(n_1129),
.D(n_1126),
.E(n_935),
.Y(n_1434)
);

AOI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1406),
.A2(n_1131),
.B1(n_1125),
.B2(n_938),
.C(n_1082),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1383),
.B(n_960),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1387),
.Y(n_1437)
);

AOI221xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1399),
.A2(n_1121),
.B1(n_1117),
.B2(n_1180),
.C(n_1125),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1408),
.B(n_1125),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1408),
.A2(n_933),
.B(n_979),
.C(n_1125),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1398),
.A2(n_1180),
.B1(n_1120),
.B2(n_1117),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1404),
.A2(n_1020),
.B1(n_1133),
.B2(n_1110),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1389),
.B(n_76),
.Y(n_1443)
);

AOI221x1_ASAP7_75t_L g1444 ( 
.A1(n_1390),
.A2(n_901),
.B1(n_951),
.B2(n_876),
.C(n_983),
.Y(n_1444)
);

NOR3xp33_ASAP7_75t_L g1445 ( 
.A(n_1381),
.B(n_901),
.C(n_887),
.Y(n_1445)
);

OAI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1390),
.A2(n_1133),
.B1(n_1090),
.B2(n_1088),
.C(n_1120),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_SL g1447 ( 
.A(n_1390),
.B(n_970),
.Y(n_1447)
);

XNOR2x1_ASAP7_75t_L g1448 ( 
.A(n_1383),
.B(n_77),
.Y(n_1448)
);

A2O1A1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1390),
.A2(n_970),
.B(n_1133),
.C(n_1120),
.Y(n_1449)
);

A2O1A1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1390),
.A2(n_970),
.B(n_1133),
.C(n_1120),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1432),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1431),
.B(n_1110),
.Y(n_1452)
);

AOI221xp5_ASAP7_75t_L g1453 ( 
.A1(n_1427),
.A2(n_1110),
.B1(n_1116),
.B2(n_1134),
.C(n_1120),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1411),
.Y(n_1454)
);

AO22x1_ASAP7_75t_L g1455 ( 
.A1(n_1413),
.A2(n_1072),
.B1(n_876),
.B2(n_951),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1423),
.Y(n_1456)
);

NOR2x1_ASAP7_75t_L g1457 ( 
.A(n_1420),
.B(n_817),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1421),
.Y(n_1458)
);

NOR2x1_ASAP7_75t_L g1459 ( 
.A(n_1448),
.B(n_835),
.Y(n_1459)
);

NOR2x1_ASAP7_75t_L g1460 ( 
.A(n_1416),
.B(n_835),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1443),
.B(n_1442),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1439),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1436),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1437),
.A2(n_1116),
.B1(n_1134),
.B2(n_959),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1440),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1434),
.B(n_80),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1422),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1430),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1417),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1426),
.A2(n_1447),
.B1(n_1412),
.B2(n_1430),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1429),
.B(n_84),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1445),
.Y(n_1472)
);

NOR2x1_ASAP7_75t_L g1473 ( 
.A(n_1424),
.B(n_835),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1444),
.Y(n_1474)
);

NOR2x1_ASAP7_75t_L g1475 ( 
.A(n_1449),
.B(n_835),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1450),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1425),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1414),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1415),
.A2(n_1116),
.B1(n_1134),
.B2(n_959),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1433),
.Y(n_1480)
);

NOR2xp67_ASAP7_75t_L g1481 ( 
.A(n_1446),
.B(n_85),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1435),
.Y(n_1482)
);

OAI211xp5_ASAP7_75t_L g1483 ( 
.A1(n_1418),
.A2(n_1072),
.B(n_1088),
.C(n_1090),
.Y(n_1483)
);

INVxp67_ASAP7_75t_SL g1484 ( 
.A(n_1419),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1441),
.A2(n_959),
.B1(n_954),
.B2(n_1072),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1428),
.Y(n_1486)
);

OA22x2_ASAP7_75t_L g1487 ( 
.A1(n_1438),
.A2(n_1121),
.B1(n_1117),
.B2(n_1090),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1411),
.B(n_89),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1468),
.B(n_97),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1456),
.Y(n_1490)
);

NOR3xp33_ASAP7_75t_SL g1491 ( 
.A(n_1471),
.B(n_101),
.C(n_104),
.Y(n_1491)
);

NOR2xp67_ASAP7_75t_L g1492 ( 
.A(n_1477),
.B(n_107),
.Y(n_1492)
);

NOR3x1_ASAP7_75t_L g1493 ( 
.A(n_1451),
.B(n_1463),
.C(n_1454),
.Y(n_1493)
);

NAND4xp75_ASAP7_75t_L g1494 ( 
.A(n_1451),
.B(n_934),
.C(n_1119),
.D(n_1130),
.Y(n_1494)
);

NAND4xp25_ASAP7_75t_L g1495 ( 
.A(n_1470),
.B(n_886),
.C(n_887),
.D(n_1090),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1460),
.B(n_934),
.Y(n_1496)
);

AOI31xp33_ASAP7_75t_L g1497 ( 
.A1(n_1457),
.A2(n_929),
.A3(n_934),
.B(n_954),
.Y(n_1497)
);

NOR2xp67_ASAP7_75t_L g1498 ( 
.A(n_1467),
.B(n_114),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_R g1499 ( 
.A(n_1458),
.B(n_116),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1488),
.B(n_120),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1469),
.B(n_121),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1466),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1462),
.Y(n_1503)
);

AOI31xp33_ASAP7_75t_L g1504 ( 
.A1(n_1472),
.A2(n_929),
.A3(n_954),
.B(n_959),
.Y(n_1504)
);

NAND4xp75_ASAP7_75t_L g1505 ( 
.A(n_1474),
.B(n_1119),
.C(n_1127),
.D(n_1130),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1465),
.B(n_122),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1475),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1482),
.B(n_152),
.Y(n_1508)
);

NOR3xp33_ASAP7_75t_L g1509 ( 
.A(n_1476),
.B(n_886),
.C(n_887),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1452),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1473),
.Y(n_1511)
);

AOI222xp33_ASAP7_75t_L g1512 ( 
.A1(n_1484),
.A2(n_1478),
.B1(n_1482),
.B2(n_1480),
.C1(n_1453),
.C2(n_1483),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_L g1513 ( 
.A(n_1459),
.B(n_835),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1481),
.B(n_1119),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1486),
.B(n_1127),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1461),
.Y(n_1516)
);

OA22x2_ASAP7_75t_L g1517 ( 
.A1(n_1464),
.A2(n_1121),
.B1(n_1117),
.B2(n_1088),
.Y(n_1517)
);

CKINVDCx6p67_ASAP7_75t_R g1518 ( 
.A(n_1455),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1479),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1487),
.Y(n_1520)
);

NAND4xp75_ASAP7_75t_L g1521 ( 
.A(n_1485),
.B(n_1130),
.C(n_1127),
.D(n_954),
.Y(n_1521)
);

OAI22x1_ASAP7_75t_L g1522 ( 
.A1(n_1516),
.A2(n_886),
.B1(n_929),
.B2(n_1121),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1499),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1492),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1490),
.B(n_157),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1503),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1502),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1489),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1507),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1493),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1506),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1508),
.Y(n_1532)
);

CKINVDCx6p67_ASAP7_75t_R g1533 ( 
.A(n_1501),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1498),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1510),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1491),
.Y(n_1536)
);

AOI22x1_ASAP7_75t_L g1537 ( 
.A1(n_1512),
.A2(n_951),
.B1(n_876),
.B2(n_846),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1500),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1518),
.A2(n_1520),
.B1(n_1514),
.B2(n_1519),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1496),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1519),
.B(n_163),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1511),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1514),
.Y(n_1543)
);

XNOR2x1_ASAP7_75t_L g1544 ( 
.A(n_1527),
.B(n_1494),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1529),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1524),
.Y(n_1546)
);

AO22x2_ASAP7_75t_L g1547 ( 
.A1(n_1530),
.A2(n_1509),
.B1(n_1496),
.B2(n_1515),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1542),
.Y(n_1548)
);

AO22x2_ASAP7_75t_L g1549 ( 
.A1(n_1539),
.A2(n_1515),
.B1(n_1521),
.B2(n_1505),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1543),
.Y(n_1550)
);

OAI22x1_ASAP7_75t_L g1551 ( 
.A1(n_1537),
.A2(n_1513),
.B1(n_1495),
.B2(n_1504),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1527),
.A2(n_1497),
.B1(n_1517),
.B2(n_1088),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1535),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1540),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_1523),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1528),
.B(n_951),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1536),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1525),
.B(n_164),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1536),
.A2(n_820),
.B1(n_951),
.B2(n_846),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1526),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1541),
.Y(n_1561)
);

AOI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1538),
.A2(n_820),
.B1(n_846),
.B2(n_831),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1538),
.A2(n_846),
.B1(n_976),
.B2(n_169),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1532),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1550),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1545),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1555),
.A2(n_1532),
.B1(n_1531),
.B2(n_1533),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1548),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1546),
.A2(n_1531),
.B1(n_1533),
.B2(n_1522),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1554),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1557),
.A2(n_831),
.B1(n_976),
.B2(n_942),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1564),
.A2(n_944),
.B1(n_942),
.B2(n_940),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1553),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1560),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1547),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1561),
.B(n_165),
.Y(n_1576)
);

AND3x4_ASAP7_75t_L g1577 ( 
.A(n_1570),
.B(n_1544),
.C(n_1547),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1565),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1575),
.Y(n_1579)
);

OAI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1567),
.A2(n_1569),
.B1(n_1566),
.B2(n_1568),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1573),
.B(n_1559),
.C(n_1556),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1576),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1574),
.A2(n_1549),
.B1(n_1563),
.B2(n_1551),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1571),
.Y(n_1584)
);

AOI22x1_ASAP7_75t_L g1585 ( 
.A1(n_1572),
.A2(n_1549),
.B1(n_1552),
.B2(n_1562),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1578),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1577),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1583),
.A2(n_1558),
.B1(n_170),
.B2(n_175),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1579),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1580),
.A2(n_168),
.B(n_176),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1587),
.A2(n_1581),
.B(n_1585),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1590),
.A2(n_1586),
.B(n_1589),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1591),
.A2(n_1588),
.B1(n_1582),
.B2(n_1584),
.Y(n_1593)
);

OAI222xp33_ASAP7_75t_L g1594 ( 
.A1(n_1592),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.C1(n_180),
.C2(n_182),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1593),
.B(n_184),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1594),
.B(n_185),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1596),
.A2(n_1595),
.B1(n_944),
.B2(n_940),
.Y(n_1597)
);


endmodule