module fake_jpeg_26602_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx5_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_4),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

A2O1A1Ixp33_ASAP7_75t_L g13 ( 
.A1(n_8),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_13),
.B(n_15),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_18),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_6),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_17),
.A2(n_19),
.B1(n_9),
.B2(n_7),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_3),
.Y(n_18)
);

NAND2x1_ASAP7_75t_SL g19 ( 
.A(n_9),
.B(n_4),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_15),
.A2(n_12),
.B1(n_6),
.B2(n_8),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_23),
.B(n_19),
.Y(n_28)
);

NOR2x1_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_24),
.Y(n_32)
);

A2O1A1O1Ixp25_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_19),
.B(n_18),
.C(n_13),
.D(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_18),
.B2(n_23),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_18),
.A3(n_14),
.B1(n_11),
.B2(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_24),
.C(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_25),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_34),
.B(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_36),
.B(n_33),
.Y(n_37)
);


endmodule