module fake_jpeg_2435_n_72 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_72);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_72;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_1),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_31),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_11),
.Y(n_44)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_22),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g46 ( 
.A(n_38),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_26),
.B1(n_20),
.B2(n_25),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_43),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_23),
.B1(n_20),
.B2(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_14),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_32),
.C(n_36),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_40),
.C(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_16),
.C(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_49),
.B1(n_46),
.B2(n_40),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_54),
.B1(n_4),
.B2(n_5),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_7),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_61),
.B(n_62),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_60),
.B(n_67),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_54),
.Y(n_72)
);


endmodule