module fake_jpeg_22605_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_2),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_14),
.B1(n_20),
.B2(n_28),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.C(n_43),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_14),
.B1(n_20),
.B2(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_17),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_25),
.C(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_20),
.B1(n_18),
.B2(n_26),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_22),
.B1(n_16),
.B2(n_36),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_53),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_58),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_25),
.B(n_23),
.C(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_62),
.B1(n_39),
.B2(n_22),
.Y(n_73)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_17),
.B(n_27),
.C(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_27),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_23),
.Y(n_83)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_24),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_74),
.B1(n_77),
.B2(n_57),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_41),
.B1(n_51),
.B2(n_53),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_51),
.B1(n_47),
.B2(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_40),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_43),
.C(n_40),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_68),
.B(n_59),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_45),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_23),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_87),
.C(n_90),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_89),
.B1(n_92),
.B2(n_57),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_91),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_57),
.B1(n_58),
.B2(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_61),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_57),
.B1(n_40),
.B2(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_83),
.C(n_80),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_85),
.C(n_87),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_8),
.C(n_11),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_105),
.B(n_106),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_78),
.B1(n_76),
.B2(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_78),
.B(n_79),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_79),
.B1(n_76),
.B2(n_75),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_19),
.B(n_81),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_8),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_6),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_115),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_116),
.C(n_117),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_9),
.C(n_12),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_9),
.C(n_12),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_119),
.B(n_121),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_124),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_99),
.B(n_105),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_115),
.C(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_126),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_125),
.B(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_120),
.C(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_3),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_103),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_136),
.B(n_5),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_131),
.B(n_3),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_139),
.Y(n_140)
);


endmodule