module fake_jpeg_11701_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_5),
.B(n_16),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_58),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_20),
.B1(n_30),
.B2(n_27),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_66),
.B1(n_23),
.B2(n_35),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_63),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_20),
.B1(n_27),
.B2(n_26),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_27),
.C(n_40),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_70),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_42),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_41),
.B(n_20),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_38),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_22),
.B1(n_71),
.B2(n_28),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_20),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_35),
.Y(n_88)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_79),
.B(n_92),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_23),
.B(n_35),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_77),
.A2(n_28),
.B(n_32),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_43),
.B1(n_42),
.B2(n_21),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_78),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_22),
.B(n_35),
.C(n_23),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_22),
.B1(n_19),
.B2(n_34),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_22),
.B1(n_21),
.B2(n_26),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_103),
.B1(n_92),
.B2(n_102),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_21),
.B1(n_26),
.B2(n_22),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_21),
.B1(n_26),
.B2(n_22),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_88),
.B(n_32),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_67),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_65),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_23),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_94),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_22),
.B1(n_29),
.B2(n_17),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_67),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_102),
.B1(n_28),
.B2(n_33),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_22),
.B1(n_29),
.B2(n_17),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_101),
.B1(n_104),
.B2(n_106),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_53),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_19),
.B1(n_34),
.B2(n_33),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_19),
.B1(n_34),
.B2(n_33),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_65),
.A2(n_36),
.B1(n_17),
.B2(n_29),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_36),
.B1(n_31),
.B2(n_32),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_50),
.A2(n_34),
.B1(n_33),
.B2(n_19),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_61),
.B1(n_53),
.B2(n_50),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_109),
.B1(n_110),
.B2(n_121),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_119),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_50),
.B1(n_62),
.B2(n_61),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_61),
.B1(n_56),
.B2(n_68),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_68),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_84),
.C(n_86),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_78),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_28),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_125),
.B(n_134),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_56),
.B1(n_64),
.B2(n_62),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_98),
.B1(n_101),
.B2(n_106),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_131),
.B(n_93),
.Y(n_142)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_64),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_117),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_79),
.A2(n_75),
.B(n_77),
.C(n_76),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_90),
.B1(n_95),
.B2(n_79),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_138),
.B1(n_140),
.B2(n_145),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_95),
.B1(n_77),
.B2(n_81),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_75),
.B1(n_100),
.B2(n_78),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_144),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_142),
.B(n_156),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_75),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_80),
.B1(n_103),
.B2(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_112),
.B(n_83),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_158),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_160),
.C(n_162),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_155),
.B1(n_164),
.B2(n_139),
.Y(n_183)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_101),
.B1(n_56),
.B2(n_85),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_161),
.B1(n_0),
.B2(n_1),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_104),
.B1(n_85),
.B2(n_62),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_86),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_89),
.Y(n_158)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_31),
.B1(n_89),
.B2(n_60),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_16),
.C(n_15),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_109),
.B1(n_108),
.B2(n_107),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_31),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_124),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_131),
.B(n_16),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_124),
.Y(n_176)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_179),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_164),
.A2(n_126),
.B1(n_118),
.B2(n_111),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_182),
.B1(n_183),
.B2(n_186),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_176),
.B(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_133),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_133),
.B1(n_110),
.B2(n_129),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_181),
.A2(n_184),
.B(n_187),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_139),
.A2(n_118),
.B1(n_111),
.B2(n_125),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_125),
.B(n_133),
.C(n_114),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_142),
.B(n_121),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_146),
.A2(n_130),
.B1(n_132),
.B2(n_60),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_114),
.B(n_130),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_135),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_190),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_130),
.B(n_135),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_189),
.A2(n_197),
.B(n_201),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_141),
.A2(n_130),
.B1(n_60),
.B2(n_15),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_195),
.B1(n_153),
.B2(n_145),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_14),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_198),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_60),
.B1(n_14),
.B2(n_2),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_0),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_136),
.B(n_0),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_143),
.B(n_14),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_149),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_3),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_60),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_4),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_144),
.A2(n_0),
.B(n_1),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_160),
.C(n_148),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_208),
.C(n_213),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_140),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_216),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_138),
.B1(n_165),
.B2(n_150),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_163),
.C(n_152),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_172),
.A2(n_137),
.B1(n_151),
.B2(n_149),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_137),
.C(n_162),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_217),
.C(n_219),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_159),
.B1(n_3),
.B2(n_4),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_159),
.C(n_3),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_195),
.B1(n_191),
.B2(n_206),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_228),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_200),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_170),
.B(n_6),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_201),
.C(n_171),
.Y(n_253)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_199),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_232),
.A2(n_234),
.B1(n_246),
.B2(n_247),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_180),
.B1(n_177),
.B2(n_186),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_235),
.A2(n_236),
.B(n_248),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_224),
.A2(n_180),
.B1(n_177),
.B2(n_175),
.Y(n_236)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_210),
.A2(n_175),
.B1(n_197),
.B2(n_170),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_238),
.A2(n_218),
.B1(n_228),
.B2(n_225),
.Y(n_277)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_208),
.B(n_207),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_244),
.B(n_222),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_176),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_252),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_205),
.B1(n_189),
.B2(n_209),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_197),
.B1(n_185),
.B2(n_181),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_212),
.A2(n_184),
.B(n_187),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_188),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_196),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_256),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_222),
.A2(n_184),
.B(n_174),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_255),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_174),
.C(n_178),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_206),
.B(n_168),
.Y(n_257)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_239),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_264),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_239),
.B(n_215),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_267),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_205),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_217),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_271),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_230),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_219),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_260),
.C(n_266),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_204),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_240),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_276),
.Y(n_279)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_246),
.B1(n_233),
.B2(n_216),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_251),
.B(n_235),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_287),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_234),
.B1(n_249),
.B2(n_247),
.Y(n_284)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_232),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_286),
.A2(n_262),
.B1(n_220),
.B2(n_204),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_249),
.B1(n_202),
.B2(n_254),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_242),
.B1(n_250),
.B2(n_238),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_253),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_295),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_242),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_265),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_251),
.C(n_248),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_267),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_7),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_306),
.B1(n_298),
.B2(n_302),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_SL g303 ( 
.A1(n_279),
.A2(n_264),
.A3(n_278),
.B1(n_269),
.B2(n_272),
.C1(n_271),
.C2(n_168),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_308),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_283),
.A2(n_278),
.B1(n_231),
.B2(n_8),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_6),
.C(n_7),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_292),
.C(n_287),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_291),
.Y(n_311)
);

AOI31xp33_ASAP7_75t_L g330 ( 
.A1(n_311),
.A2(n_315),
.A3(n_13),
.B(n_11),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_302),
.A2(n_285),
.B1(n_294),
.B2(n_295),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_313),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_292),
.Y(n_315)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_316),
.Y(n_327)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_281),
.C(n_280),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_281),
.C(n_10),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_320),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_305),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_10),
.B(n_11),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_321),
.A2(n_307),
.B1(n_296),
.B2(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_326),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_314),
.B1(n_317),
.B2(n_319),
.Y(n_332)
);

AOI31xp67_ASAP7_75t_L g328 ( 
.A1(n_310),
.A2(n_10),
.A3(n_11),
.B(n_12),
.Y(n_328)
);

OAI21x1_ASAP7_75t_L g336 ( 
.A1(n_328),
.A2(n_330),
.B(n_13),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_10),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_12),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_332),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_316),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_335),
.C(n_334),
.Y(n_337)
);

AND2x2_ASAP7_75t_SL g335 ( 
.A(n_322),
.B(n_313),
.Y(n_335)
);

A2O1A1O1Ixp25_ASAP7_75t_L g339 ( 
.A1(n_336),
.A2(n_328),
.B(n_327),
.C(n_325),
.D(n_13),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_337),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_338),
.C(n_326),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_318),
.C(n_339),
.Y(n_343)
);


endmodule