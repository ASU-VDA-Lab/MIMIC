module fake_jpeg_15753_n_294 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_0),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_36),
.B(n_23),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_31),
.B1(n_27),
.B2(n_30),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_53),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_57),
.Y(n_79)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_31),
.B1(n_29),
.B2(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_66),
.B(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_68),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_20),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_70),
.B(n_76),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_74),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_34),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_81),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_22),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_38),
.C(n_40),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_88),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_34),
.C(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_101),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_22),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_52),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_21),
.B1(n_24),
.B2(n_19),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_90),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_30),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_92),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_96),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_45),
.B(n_23),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_23),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_97),
.A2(n_27),
.B1(n_57),
.B2(n_49),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_17),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_111),
.B1(n_112),
.B2(n_88),
.Y(n_147)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_13),
.Y(n_105)
);

OAI221xp5_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_18),
.B1(n_25),
.B2(n_21),
.C(n_3),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_27),
.B1(n_40),
.B2(n_28),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_120),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_24),
.B1(n_19),
.B2(n_18),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_28),
.B1(n_21),
.B2(n_25),
.Y(n_112)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_118),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_71),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_71),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_124),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_78),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_76),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_78),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_77),
.B1(n_68),
.B2(n_84),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_70),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_87),
.B1(n_64),
.B2(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_114),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_160),
.B(n_122),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_108),
.A2(n_87),
.B1(n_64),
.B2(n_86),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_147),
.A2(n_149),
.B1(n_153),
.B2(n_159),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_108),
.A2(n_64),
.B1(n_79),
.B2(n_91),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_92),
.B1(n_98),
.B2(n_79),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_122),
.B1(n_119),
.B2(n_118),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_156),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_65),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_106),
.B(n_120),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_103),
.C(n_117),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_111),
.A2(n_89),
.B1(n_93),
.B2(n_2),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_0),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_117),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_162),
.C(n_172),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_130),
.B(n_127),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_174),
.B1(n_185),
.B2(n_160),
.Y(n_201)
);

XOR2x2_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_105),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_175),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_127),
.C(n_130),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_173),
.B(n_153),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_105),
.B(n_0),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_112),
.C(n_113),
.Y(n_175)
);

AOI32xp33_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_124),
.A3(n_104),
.B1(n_113),
.B2(n_100),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_180),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_124),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_181),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_65),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_55),
.C(n_121),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_139),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_1),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_135),
.A2(n_121),
.B1(n_104),
.B2(n_2),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_150),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_183),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_197),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_189),
.A2(n_148),
.B1(n_151),
.B2(n_147),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_203),
.B1(n_207),
.B2(n_170),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_194),
.A2(n_198),
.B(n_170),
.Y(n_226)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_163),
.B(n_133),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_168),
.B1(n_164),
.B2(n_177),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_135),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_171),
.A2(n_146),
.B1(n_154),
.B2(n_156),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_104),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_142),
.B1(n_1),
.B2(n_0),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_212),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_1),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_99),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_161),
.C(n_172),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_216),
.C(n_220),
.Y(n_247)
);

XOR2x2_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_175),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_215),
.A2(n_217),
.B(n_198),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_181),
.C(n_182),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_174),
.B(n_165),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_55),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_206),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_230),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_199),
.B(n_205),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_167),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_207),
.B1(n_168),
.B2(n_173),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_195),
.B(n_198),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_233),
.A2(n_238),
.B1(n_240),
.B2(n_214),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_234),
.B(n_244),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_236),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_222),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_194),
.B(n_191),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_226),
.A2(n_210),
.B(n_192),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_225),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_227),
.B(n_197),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_245),
.Y(n_258)
);

OAI321xp33_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_212),
.A3(n_211),
.B1(n_203),
.B2(n_201),
.C(n_209),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_8),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_230),
.B(n_229),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_248),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_216),
.B1(n_223),
.B2(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_255),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_239),
.C(n_233),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_225),
.B1(n_4),
.B2(n_5),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_12),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_9),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_238),
.A2(n_6),
.B(n_7),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_9),
.B(n_10),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_10),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_14),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_235),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_261),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_239),
.B(n_247),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_272),
.B(n_256),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_270),
.A2(n_254),
.B(n_250),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_257),
.B1(n_15),
.B2(n_16),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_12),
.B(n_13),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_255),
.C(n_251),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_277),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_253),
.B(n_14),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_265),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_271),
.B(n_267),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_279),
.B(n_280),
.Y(n_282)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_284),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_276),
.C(n_253),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_275),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_287),
.A2(n_283),
.B(n_15),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_289),
.B(n_288),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_291),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);


endmodule