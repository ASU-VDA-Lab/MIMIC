module fake_jpeg_28612_n_409 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_409);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_25),
.B(n_23),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_58),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_11),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_27),
.B(n_11),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_82),
.Y(n_89)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_75),
.Y(n_90)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_11),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx5_ASAP7_75t_SL g113 ( 
.A(n_83),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_47),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_119),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_46),
.B1(n_42),
.B2(n_31),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_105),
.A2(n_77),
.B1(n_79),
.B2(n_67),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_33),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_37),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_69),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_115),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_45),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_36),
.B1(n_34),
.B2(n_40),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_34),
.B1(n_40),
.B2(n_39),
.Y(n_149)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_31),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_45),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_145),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_57),
.B1(n_55),
.B2(n_61),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_153),
.B1(n_157),
.B2(n_164),
.Y(n_173)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_142),
.Y(n_189)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_152),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_148),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_89),
.A2(n_44),
.B(n_43),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_147),
.Y(n_168)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_151),
.B1(n_158),
.B2(n_160),
.Y(n_170)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_95),
.B(n_33),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_155),
.B(n_161),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_95),
.B(n_30),
.C(n_62),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_115),
.C(n_24),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_66),
.B1(n_64),
.B2(n_46),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_36),
.B1(n_40),
.B2(n_46),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_113),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_37),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_88),
.B(n_44),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_165),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_110),
.A2(n_42),
.B1(n_28),
.B2(n_32),
.Y(n_164)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_110),
.B1(n_118),
.B2(n_124),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_124),
.B1(n_129),
.B2(n_166),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_181),
.Y(n_197)
);

INVx2_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_91),
.C(n_32),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_120),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_97),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_101),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_106),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_176),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_192),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_157),
.B(n_153),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_199),
.B(n_207),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_204),
.B1(n_189),
.B2(n_175),
.Y(n_217)
);

NOR2x1p5_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_164),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_205),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_154),
.B1(n_143),
.B2(n_93),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_201),
.A2(n_207),
.B1(n_189),
.B2(n_190),
.Y(n_214)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_129),
.B1(n_111),
.B2(n_132),
.Y(n_204)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_165),
.B1(n_151),
.B2(n_134),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_209),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_145),
.B1(n_117),
.B2(n_133),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_169),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_169),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_174),
.B1(n_186),
.B2(n_187),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_175),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_215),
.B(n_229),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_220),
.B1(n_223),
.B2(n_195),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_178),
.B(n_184),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_205),
.A2(n_179),
.B1(n_171),
.B2(n_148),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_198),
.B1(n_159),
.B2(n_90),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_217),
.A2(n_194),
.B1(n_210),
.B2(n_193),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_181),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_219),
.B(n_211),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_201),
.A2(n_172),
.B1(n_182),
.B2(n_168),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_225),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_172),
.B1(n_185),
.B2(n_191),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_199),
.A2(n_186),
.B1(n_183),
.B2(n_171),
.Y(n_229)
);

OAI32xp33_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_198),
.A3(n_205),
.B1(n_175),
.B2(n_179),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_196),
.B(n_176),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_200),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_183),
.C(n_135),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_211),
.C(n_210),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_227),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_234),
.B(n_243),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_249),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_208),
.C(n_196),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_229),
.Y(n_270)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_179),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_239),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_248),
.B1(n_255),
.B2(n_222),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_227),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_225),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_246),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_218),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_205),
.B(n_204),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_216),
.B(n_230),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_213),
.A2(n_200),
.B1(n_193),
.B2(n_211),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_214),
.A2(n_211),
.B1(n_193),
.B2(n_205),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_250),
.A2(n_252),
.B1(n_217),
.B2(n_175),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_212),
.A2(n_228),
.B1(n_223),
.B2(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_141),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_256),
.B(n_125),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_278),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_261),
.A2(n_273),
.B(n_275),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_212),
.Y(n_263)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_252),
.A2(n_229),
.B1(n_232),
.B2(n_218),
.Y(n_265)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_265),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_266),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_232),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_279),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_274),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_277),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_240),
.B1(n_248),
.B2(n_254),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_242),
.A2(n_163),
.B(n_134),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_179),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_242),
.A2(n_163),
.B(n_123),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_247),
.A2(n_123),
.B1(n_116),
.B2(n_131),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_250),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_226),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_244),
.B1(n_233),
.B2(n_241),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_304),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_293),
.B1(n_262),
.B2(n_28),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_226),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_285),
.B(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_236),
.Y(n_286)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_258),
.B(n_237),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_288),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_290),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_271),
.B1(n_272),
.B2(n_261),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_251),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_292),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_256),
.B1(n_234),
.B2(n_235),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_249),
.C(n_253),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_298),
.C(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_136),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_275),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_125),
.C(n_112),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_24),
.Y(n_299)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

INVx3_ASAP7_75t_SL g300 ( 
.A(n_266),
.Y(n_300)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_264),
.B(n_38),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_277),
.B(n_25),
.CI(n_38),
.CON(n_304),
.SN(n_304)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_305),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_322),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_312),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_291),
.B1(n_292),
.B2(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_316),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_297),
.C(n_294),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_318),
.C(n_326),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_260),
.B1(n_264),
.B2(n_280),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_317),
.A2(n_282),
.B1(n_296),
.B2(n_287),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_262),
.C(n_136),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_281),
.A2(n_136),
.B(n_1),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_321),
.B(n_323),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_40),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_281),
.A2(n_13),
.B(n_1),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_90),
.C(n_98),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_292),
.A2(n_12),
.B(n_3),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_304),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_329),
.Y(n_351)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_333),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_308),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_337),
.Y(n_359)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_336),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_301),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_340),
.Y(n_353)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

FAx1_ASAP7_75t_SL g341 ( 
.A(n_308),
.B(n_284),
.CI(n_290),
.CON(n_341),
.SN(n_341)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_341),
.B(n_342),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_300),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_307),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_345),
.A2(n_305),
.B1(n_304),
.B2(n_326),
.Y(n_358)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_327),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_346),
.A2(n_312),
.B1(n_3),
.B2(n_4),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_314),
.C(n_306),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_349),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_318),
.C(n_316),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_337),
.A2(n_328),
.B1(n_320),
.B2(n_313),
.Y(n_350)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_350),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_344),
.A2(n_310),
.B1(n_328),
.B2(n_311),
.Y(n_354)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_354),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_335),
.A2(n_301),
.B(n_315),
.Y(n_357)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_357),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_347),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_360),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_330),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_362),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_333),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_338),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_367),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_347),
.A2(n_341),
.B1(n_332),
.B2(n_338),
.Y(n_366)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_366),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_330),
.C(n_5),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_370),
.B(n_371),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_355),
.C(n_357),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_372),
.B(n_14),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_368),
.B(n_356),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_375),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_353),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_354),
.C(n_350),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_377),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_353),
.Y(n_377)
);

NAND3xp33_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_14),
.C(n_5),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_378),
.A2(n_381),
.B(n_25),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_380),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_369),
.A2(n_14),
.B(n_5),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_384),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_15),
.Y(n_384)
);

AOI21x1_ASAP7_75t_SL g385 ( 
.A1(n_378),
.A2(n_15),
.B(n_6),
.Y(n_385)
);

NOR3xp33_ASAP7_75t_L g396 ( 
.A(n_385),
.B(n_7),
.C(n_9),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_391),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_374),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_390),
.A2(n_7),
.B(n_9),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_382),
.B(n_13),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_17),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_393),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_389),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_398),
.C(n_399),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_396),
.B(n_397),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_18),
.C(n_19),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_395),
.A2(n_390),
.B(n_386),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_401),
.B(n_21),
.Y(n_404)
);

OAI31xp33_ASAP7_75t_SL g403 ( 
.A1(n_402),
.A2(n_18),
.A3(n_19),
.B(n_20),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_403),
.B(n_404),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_405),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_400),
.C(n_19),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_407),
.B(n_21),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_0),
.B(n_406),
.Y(n_409)
);


endmodule