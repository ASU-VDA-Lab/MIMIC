module fake_jpeg_3669_n_215 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_215);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_10),
.B(n_11),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_0),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_55),
.B1(n_66),
.B2(n_64),
.Y(n_83)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_60),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_71),
.B1(n_53),
.B2(n_69),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_65),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_53),
.B1(n_71),
.B2(n_69),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_94),
.B1(n_62),
.B2(n_64),
.Y(n_109)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_69),
.B1(n_71),
.B2(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_97),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_81),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_106),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_80),
.B1(n_54),
.B2(n_59),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_89),
.B1(n_88),
.B2(n_80),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_62),
.B(n_70),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_102),
.B(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_58),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_72),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_63),
.Y(n_124)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_93),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_132),
.B1(n_122),
.B2(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_123),
.Y(n_135)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_33),
.Y(n_156)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_130),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_0),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_77),
.B1(n_55),
.B2(n_90),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_77),
.B1(n_86),
.B2(n_67),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_67),
.B1(n_73),
.B2(n_50),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_134),
.B(n_48),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_137),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_110),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_146),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_77),
.B(n_67),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_150),
.B1(n_4),
.B2(n_5),
.Y(n_164)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_155),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_47),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_51),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_36),
.C(n_35),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_1),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_51),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_153),
.B1(n_146),
.B2(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_46),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_25),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_119),
.B(n_1),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_51),
.B(n_45),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_159),
.B(n_168),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_43),
.B(n_40),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_157),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_154),
.B1(n_139),
.B2(n_9),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_173),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_169),
.B1(n_19),
.B2(n_13),
.Y(n_189)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_27),
.B(n_26),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_178),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_24),
.B(n_23),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_20),
.C(n_7),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_147),
.C(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_179),
.B(n_163),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_187),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_6),
.C(n_8),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_182),
.C(n_184),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_188),
.A2(n_189),
.B1(n_166),
.B2(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_191),
.B(n_193),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_196),
.Y(n_200)
);

AO221x1_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_172),
.B1(n_175),
.B2(n_174),
.C(n_15),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_175),
.B(n_171),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_197),
.A2(n_188),
.B(n_13),
.Y(n_203)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_177),
.C(n_173),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_188),
.B1(n_181),
.B2(n_14),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_203),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_204),
.A2(n_195),
.B1(n_199),
.B2(n_15),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_200),
.Y(n_210)
);

OAI321xp33_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_206),
.A3(n_202),
.B1(n_201),
.B2(n_18),
.C(n_12),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_212),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_209),
.B1(n_14),
.B2(n_16),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_12),
.Y(n_215)
);


endmodule