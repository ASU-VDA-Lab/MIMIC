module fake_ibex_502_n_5014 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_5014);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_5014;

wire n_4557;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_4204;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_962;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_3479;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_2343;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_4423;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3472;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_4801;
wire n_3639;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_4569;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_4567;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1306;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_3565;
wire n_3883;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_2147;
wire n_2253;
wire n_4479;
wire n_3858;
wire n_4173;
wire n_1078;
wire n_4422;
wire n_1865;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_1653;
wire n_1375;
wire n_1118;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_3060;
wire n_4124;
wire n_971;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_3293;
wire n_2550;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_1108;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_1209;
wire n_3732;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_1121;
wire n_4823;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_4757;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_1042;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_1987;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_4374;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3529;
wire n_3222;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_1008;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_1210;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_1246;
wire n_4231;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_2361;
wire n_4128;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_3119;
wire n_2590;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_3544;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_2046;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_4679;
wire n_1345;
wire n_4456;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_1471;
wire n_3441;
wire n_4559;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_2010;
wire n_2733;
wire n_3796;
wire n_1836;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_4024;
wire n_3975;
wire n_3164;
wire n_1448;
wire n_3034;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_1967;
wire n_1095;
wire n_3834;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_3428;
wire n_2427;
wire n_1127;
wire n_947;
wire n_1004;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_2422;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_972;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_3339;
wire n_3673;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_1340;
wire n_2562;
wire n_3269;
wire n_2223;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_4339;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3686;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_1517;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_977;
wire n_1895;
wire n_1860;
wire n_1763;
wire n_3912;
wire n_1607;
wire n_2959;
wire n_2420;
wire n_2380;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1021;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_4729;
wire n_1617;
wire n_2639;
wire n_3099;
wire n_1001;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_1017;
wire n_2049;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_4417;
wire n_1550;
wire n_1169;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1072;
wire n_2194;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_3096;
wire n_2059;
wire n_1278;
wire n_4730;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_950;
wire n_4282;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_4919;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_2871;
wire n_2764;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_985;
wire n_4611;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_1459;
wire n_4032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_995;
wire n_1303;
wire n_1994;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_946;
wire n_4895;
wire n_3354;
wire n_4069;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_2574;
wire n_1887;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_2228;
wire n_4474;
wire n_1518;
wire n_4350;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_1010;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_4911;
wire n_1329;
wire n_2409;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_3742;
wire n_3532;
wire n_4686;
wire n_4682;
wire n_2914;
wire n_1833;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_4733;
wire n_987;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_1166;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_4962;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_4644;
wire n_1012;
wire n_960;
wire n_4412;
wire n_4266;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_1230;
wire n_3622;
wire n_3857;
wire n_2357;
wire n_4354;
wire n_2937;
wire n_3728;
wire n_4401;
wire n_4727;
wire n_4296;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1033;
wire n_990;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_4539;
wire n_1205;
wire n_2969;
wire n_3550;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_1002;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_3662;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_3789;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_984;
wire n_2978;
wire n_3502;
wire n_3935;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_4926;
wire n_4688;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_1930;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_969;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_3484;
wire n_2485;
wire n_4477;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_948;
wire n_3726;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_4433;
wire n_3030;
wire n_4503;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_3221;
wire n_3210;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_1301;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_4610;
wire n_4067;
wire n_4997;
wire n_4393;
wire n_3777;
wire n_4553;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_2257;
wire n_4856;
wire n_1467;
wire n_3217;
wire n_2511;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_4649;
wire n_3832;
wire n_3508;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_3633;
wire n_1731;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_2076;
wire n_974;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_959;
wire n_1312;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_965;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_2176;
wire n_2805;
wire n_2319;
wire n_3757;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_3787;
wire n_3445;
wire n_2080;
wire n_2554;
wire n_1676;
wire n_1013;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_1014;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_3394;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_3488;
wire n_2832;
wire n_4991;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_2142;
wire n_3703;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_954;
wire n_4734;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_1729;
wire n_998;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_4579;
wire n_943;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1775;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_3074;
wire n_4640;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_2170;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_997;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_3350;
wire n_4873;
wire n_945;
wire n_3936;
wire n_1560;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_4636;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_4609;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_1011;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_2442;
wire n_1067;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_1894;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_4699;
wire n_1331;
wire n_1223;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_1294;
wire n_1351;
wire n_1380;
wire n_3336;
wire n_1291;
wire n_3763;
wire n_4284;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_1662;
wire n_3443;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_1660;
wire n_4000;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_1962;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_2309;
wire n_2274;
wire n_3712;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_4643;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_1241;
wire n_2589;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_1238;
wire n_3959;
wire n_976;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_1644;
wire n_4586;
wire n_3860;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_1149;
wire n_4905;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_1261;
wire n_3327;
wire n_1114;
wire n_3647;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1018;
wire n_1669;
wire n_1885;
wire n_1989;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_4408;
wire n_1175;
wire n_1221;
wire n_3875;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_4565;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_1507;
wire n_1206;
wire n_3576;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_956;
wire n_4597;
wire n_1812;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_1798;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_941;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_3050;
wire n_2666;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_4516;
wire n_2913;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_4196;
wire n_2371;
wire n_3898;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_5013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_2671;
wire n_3296;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_3207;
wire n_953;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_3036;
wire n_5012;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_3332;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_3861;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_955;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3738;
wire n_1640;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_1355;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_4590;
wire n_4602;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_1780;
wire n_1091;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_1743;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_4883;
wire n_1079;
wire n_3559;
wire n_4943;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_3750;
wire n_3838;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_4159;
wire n_4372;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_1233;
wire n_4360;
wire n_3653;
wire n_4897;
wire n_963;
wire n_2139;
wire n_3693;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_1829;
wire n_1338;
wire n_1327;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_2565;
wire n_4201;
wire n_1636;
wire n_1687;
wire n_4584;
wire n_3184;
wire n_4155;
wire n_3890;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1680;
wire n_1195;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_3641;
wire n_4887;
wire n_3996;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_1841;
wire n_2685;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_3722;
wire n_3802;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_4806;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_1007;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_3765;
wire n_2216;
wire n_4259;
wire n_1620;
wire n_3518;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_2899;
wire n_3351;
wire n_2008;
wire n_2859;
wire n_2564;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_1764;
wire n_1019;
wire n_1250;
wire n_1190;
wire n_4598;
wire n_3259;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_2114;
wire n_1609;
wire n_3530;
wire n_1132;
wire n_4548;
wire n_1803;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_4999;
wire n_2660;
wire n_5006;
wire n_4604;
wire n_3467;
wire n_4240;
wire n_2219;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_2539;
wire n_1701;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_3282;
wire n_1003;
wire n_2708;
wire n_2748;
wire n_2224;
wire n_2233;
wire n_2499;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_1553;
wire n_3542;
wire n_1090;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_3171;
wire n_1733;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_1189;
wire n_4995;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_4205;
wire n_3790;
wire n_2404;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_4504;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_1236;
wire n_3412;
wire n_1712;
wire n_4537;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_4184;
wire n_2468;
wire n_3248;
wire n_2606;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_4876;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_4747;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_2481;
wire n_4409;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_3396;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_2977;
wire n_1682;
wire n_3599;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_4152;
wire n_1352;
wire n_2328;
wire n_4587;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_4500;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_2419;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_951;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_4496;
wire n_1528;
wire n_3840;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_1413;
wire n_2464;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_2414;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_4316;
wire n_3328;
wire n_2763;
wire n_994;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_4306;
wire n_2997;
wire n_3735;
wire n_961;
wire n_2127;
wire n_3028;
wire n_3228;
wire n_3706;
wire n_1432;
wire n_3322;
wire n_996;
wire n_1174;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_2694;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_982;
wire n_2180;
wire n_3376;
wire n_2617;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_2086;
wire n_4832;
wire n_3666;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_2108;
wire n_2535;
wire n_2945;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_2196;
wire n_1538;
wire n_3773;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_1124;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_1642;
wire n_2447;
wire n_3358;
wire n_2894;
wire n_2587;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_3410;
wire n_975;
wire n_4900;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_2299;
wire n_2078;
wire n_3709;
wire n_3011;
wire n_2315;
wire n_3623;
wire n_2157;
wire n_3446;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_4334;
wire n_2211;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_1501;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_2893;
wire n_2009;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_1005;
wire n_4581;
wire n_4618;
wire n_1105;
wire n_2898;
wire n_2519;
wire n_2231;
wire n_1000;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_4670;
wire n_4982;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_1939;
wire n_4053;
wire n_4279;
wire n_3937;
wire n_3303;
wire n_4555;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_1693;
wire n_2081;
wire n_2993;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_3989;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_967;
wire n_4263;
wire n_3725;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_1336;
wire n_1358;
wire n_3318;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_3430;
wire n_1685;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_1074;
wire n_1462;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_1398;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_1692;
wire n_4796;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_3837;
wire n_4841;
wire n_3076;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2855;
wire n_2653;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_2331;
wire n_1600;
wire n_4701;
wire n_4088;
wire n_2136;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_4972;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_1822;
wire n_1804;
wire n_1581;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_2262;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_4327;
wire n_2656;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_1016;
wire n_4465;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_983;
wire n_4224;
wire n_4868;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_4387;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_992;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_4967;
wire n_1080;
wire n_2290;
wire n_957;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_4668;
wire n_2383;
wire n_2640;
wire n_1492;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_2230;
wire n_3033;
wire n_2151;
wire n_4912;
wire n_1971;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_2571;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_989;
wire n_1668;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_4311;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_1606;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_4650;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_979;
wire n_1999;
wire n_3810;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_2826;
wire n_2112;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_4671;
wire n_1326;
wire n_4981;
wire n_978;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_3618;
wire n_2727;
wire n_2719;
wire n_2213;
wire n_3521;
wire n_2723;
wire n_4054;
wire n_1569;
wire n_4012;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_2292;
wire n_3560;
wire n_1742;
wire n_1818;
wire n_3847;
wire n_2203;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_2646;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_4755;
wire n_3827;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_4996;
wire n_4136;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1360;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_1036;
wire n_1106;
wire n_4655;
wire n_1634;
wire n_1452;
wire n_4953;
wire n_4570;
wire n_3966;
wire n_4293;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_2819;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_3436;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_4527;
wire n_2877;
wire n_1996;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_4407;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_3680;
wire n_3624;
wire n_4989;
wire n_2467;
wire n_4292;
wire n_3145;
wire n_2662;
wire n_3872;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_1566;
wire n_1464;
wire n_944;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_4929;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_1009;
wire n_2160;
wire n_2991;
wire n_2699;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_942;
wire n_4042;
wire n_2525;
wire n_4624;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_4958;
wire n_4297;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_2095;
wire n_2486;
wire n_2521;
wire n_1574;
wire n_4764;
wire n_4899;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_1357;
wire n_4566;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_2117;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_3638;
wire n_2106;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_964;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_4133;
wire n_3985;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_2745;
wire n_2110;
wire n_3747;
wire n_991;
wire n_1323;
wire n_3710;
wire n_1429;
wire n_3209;
wire n_2026;
wire n_3588;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_2642;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_4048;
wire n_4084;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_2849;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_4860;
wire n_4438;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_3047;
wire n_2610;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_4383;
wire n_2709;
wire n_2244;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_2665;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_993;
wire n_2581;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_1406;
wire n_3591;
wire n_2137;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_3139;
wire n_4715;
wire n_4222;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_1167;
wire n_3231;
wire n_3138;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_3454;
wire n_4143;
wire n_4410;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_1513;
wire n_1788;
wire n_2348;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_2248;
wire n_958;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_3846;
wire n_4328;
wire n_1433;
wire n_1907;
wire n_3994;
wire n_2135;
wire n_1088;
wire n_1102;
wire n_4487;
wire n_1165;
wire n_4148;
wire n_3066;
wire n_2869;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_2667;
wire n_1565;
wire n_2325;
wire n_3346;
wire n_3391;
wire n_1547;
wire n_1542;
wire n_1362;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_3045;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_2021;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_2061;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_3042;
wire n_2561;
wire n_2491;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_4811;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_1759;
wire n_2096;
wire n_2296;
wire n_1911;
wire n_2870;
wire n_4869;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_1419;
wire n_4738;
wire n_980;
wire n_1193;
wire n_3557;
wire n_2928;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_4086;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_999;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_1499;
wire n_2155;
wire n_966;
wire n_3938;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_3053;
wire n_1039;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_1762;
wire n_940;
wire n_4944;
wire n_4468;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_1791;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_1164;
wire n_3749;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_4280;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_1665;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_4978;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_1417;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_1410;
wire n_988;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_857),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_621),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_315),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_229),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_832),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_874),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_521),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_260),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_840),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_128),
.Y(n_949)
);

BUFx10_ASAP7_75t_L g950 ( 
.A(n_919),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_788),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_672),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_885),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_536),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_59),
.Y(n_955)
);

CKINVDCx14_ASAP7_75t_R g956 ( 
.A(n_835),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_871),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_727),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_780),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_446),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_543),
.Y(n_961)
);

BUFx5_ASAP7_75t_L g962 ( 
.A(n_934),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_368),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_851),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_526),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_331),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_854),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_548),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_858),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_841),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_614),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_444),
.Y(n_972)
);

CKINVDCx16_ASAP7_75t_R g973 ( 
.A(n_151),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_343),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_897),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_130),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_527),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_685),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_269),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_325),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_656),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_884),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_3),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_206),
.Y(n_984)
);

CKINVDCx16_ASAP7_75t_R g985 ( 
.A(n_54),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_535),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_75),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_457),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_16),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_241),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_270),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_913),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_817),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_477),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_538),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_769),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_763),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_922),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_657),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_906),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_587),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_836),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_490),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_722),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_522),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_875),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_80),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_4),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_557),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_491),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_914),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_18),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_927),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_491),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_111),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_343),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_444),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_930),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_298),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_197),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_929),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_460),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_514),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_63),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_821),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_779),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_682),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_804),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_483),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_385),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_136),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_34),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_864),
.Y(n_1033)
);

BUFx5_ASAP7_75t_L g1034 ( 
.A(n_860),
.Y(n_1034)
);

BUFx8_ASAP7_75t_SL g1035 ( 
.A(n_920),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_62),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_932),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_119),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_23),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_445),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_56),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_639),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_846),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_523),
.Y(n_1044)
);

BUFx10_ASAP7_75t_L g1045 ( 
.A(n_790),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_684),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_577),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_567),
.Y(n_1048)
);

CKINVDCx14_ASAP7_75t_R g1049 ( 
.A(n_88),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_237),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_6),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_928),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_750),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_903),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_84),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_76),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_231),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_898),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_619),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_140),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_870),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_879),
.Y(n_1062)
);

CKINVDCx16_ASAP7_75t_R g1063 ( 
.A(n_834),
.Y(n_1063)
);

CKINVDCx16_ASAP7_75t_R g1064 ( 
.A(n_645),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_165),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_432),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_353),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_843),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_563),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_597),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_508),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_96),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_706),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_304),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_238),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_405),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_480),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_851),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_839),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_856),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_292),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_359),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_805),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_760),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_901),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_402),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_806),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_81),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_343),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_775),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_799),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_859),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_456),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_570),
.Y(n_1094)
);

BUFx10_ASAP7_75t_L g1095 ( 
.A(n_853),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_633),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_70),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_540),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_926),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_753),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_131),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_726),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_913),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_597),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_933),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_890),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_268),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_532),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_305),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_848),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_622),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_588),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_207),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_223),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_679),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_296),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_475),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_246),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_470),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_685),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_285),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_634),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_749),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_565),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_403),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_108),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_920),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_360),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_456),
.Y(n_1129)
);

INVxp67_ASAP7_75t_SL g1130 ( 
.A(n_918),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_874),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_279),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_900),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_305),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_916),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_382),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_9),
.Y(n_1137)
);

CKINVDCx16_ASAP7_75t_R g1138 ( 
.A(n_67),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_822),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_423),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_195),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_551),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_72),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_654),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_282),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_935),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_333),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_847),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_182),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_937),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_815),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_807),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_684),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_900),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_93),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_292),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_899),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_289),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_459),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_846),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_476),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_669),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_886),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_601),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_566),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_936),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_434),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_31),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_818),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_896),
.Y(n_1171)
);

CKINVDCx16_ASAP7_75t_R g1172 ( 
.A(n_114),
.Y(n_1172)
);

BUFx5_ASAP7_75t_L g1173 ( 
.A(n_555),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_77),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_395),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_667),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_551),
.Y(n_1177)
);

CKINVDCx14_ASAP7_75t_R g1178 ( 
.A(n_637),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_72),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_830),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_712),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_530),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_812),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_534),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_803),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_451),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_272),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_98),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_910),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_924),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_379),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_124),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_902),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_596),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_328),
.Y(n_1195)
);

CKINVDCx16_ASAP7_75t_R g1196 ( 
.A(n_828),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_893),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_800),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_86),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_814),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_37),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_334),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_820),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_750),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_71),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_509),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_755),
.Y(n_1207)
);

BUFx2_ASAP7_75t_SL g1208 ( 
.A(n_552),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_36),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_933),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_712),
.Y(n_1211)
);

BUFx10_ASAP7_75t_L g1212 ( 
.A(n_24),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_582),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_891),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_669),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_262),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_278),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_159),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_619),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_178),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_813),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_203),
.Y(n_1222)
);

BUFx10_ASAP7_75t_L g1223 ( 
.A(n_49),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_714),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_289),
.Y(n_1225)
);

BUFx10_ASAP7_75t_L g1226 ( 
.A(n_880),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_492),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_178),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_16),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_260),
.Y(n_1230)
);

INVx4_ASAP7_75t_R g1231 ( 
.A(n_179),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_14),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_731),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_660),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_707),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_60),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_931),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_554),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_17),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_45),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_274),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_274),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_173),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_508),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_435),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_372),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_726),
.Y(n_1247)
);

BUFx2_ASAP7_75t_SL g1248 ( 
.A(n_798),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_530),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_501),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_429),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_867),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_465),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_41),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_191),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_15),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_769),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_763),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_109),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_863),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_352),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_707),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_845),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_827),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_811),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_90),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_888),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_270),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_801),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_87),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_909),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_614),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_661),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_782),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_0),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_221),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_545),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_592),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_315),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_473),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_827),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_440),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_925),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_623),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_826),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_859),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_895),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_888),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_555),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_476),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_824),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_283),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_264),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_917),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_500),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_197),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_892),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_862),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_322),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_825),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_345),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_95),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_646),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_849),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_790),
.Y(n_1305)
);

BUFx10_ASAP7_75t_L g1306 ( 
.A(n_538),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_782),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_70),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_444),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_866),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_514),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_861),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_877),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_863),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_903),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_659),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_869),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_717),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_186),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_627),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_32),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_912),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_624),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_578),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_838),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_311),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_245),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_818),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_429),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_844),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_280),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_222),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_224),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_248),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_683),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_181),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_628),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_789),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_234),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_883),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_725),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_415),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_775),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_209),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_492),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_651),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_445),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_883),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_558),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_376),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_369),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_850),
.Y(n_1352)
);

BUFx8_ASAP7_75t_SL g1353 ( 
.A(n_865),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_269),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_297),
.Y(n_1355)
);

CKINVDCx16_ASAP7_75t_R g1356 ( 
.A(n_795),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_615),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_572),
.Y(n_1358)
);

BUFx10_ASAP7_75t_L g1359 ( 
.A(n_465),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_606),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_626),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_509),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_298),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_50),
.Y(n_1364)
);

CKINVDCx11_ASAP7_75t_R g1365 ( 
.A(n_447),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_709),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_887),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_872),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_320),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_876),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_781),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_715),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_833),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_857),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_930),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_921),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_417),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_761),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_776),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_285),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_337),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_808),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_137),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_809),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_598),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_816),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_881),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_320),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_617),
.Y(n_1389)
);

BUFx8_ASAP7_75t_SL g1390 ( 
.A(n_567),
.Y(n_1390)
);

INVxp67_ASAP7_75t_SL g1391 ( 
.A(n_567),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_470),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_28),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_912),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_770),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_451),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_528),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_617),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_353),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_228),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_882),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_716),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_536),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_223),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_802),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_359),
.Y(n_1406)
);

CKINVDCx16_ASAP7_75t_R g1407 ( 
.A(n_830),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_590),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_550),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_455),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_819),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_713),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_904),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_367),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_831),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_563),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_26),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_672),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_303),
.Y(n_1419)
);

INVxp33_ASAP7_75t_SL g1420 ( 
.A(n_506),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_378),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_938),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_695),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_114),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_703),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_407),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_333),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_923),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_668),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_855),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_741),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_613),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_630),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_540),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_30),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_474),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_568),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_270),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_301),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_635),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_710),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_931),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_435),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_70),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_67),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_797),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_622),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_460),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_11),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_87),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_810),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_132),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_899),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_878),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_180),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_577),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_486),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_894),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_917),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_695),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_873),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_579),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_82),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_166),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_83),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_74),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_110),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_829),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_504),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_477),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_915),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_566),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_36),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_697),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_339),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_812),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_63),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_641),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_908),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_305),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_394),
.Y(n_1481)
);

BUFx10_ASAP7_75t_L g1482 ( 
.A(n_473),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_97),
.Y(n_1483)
);

INVxp67_ASAP7_75t_SL g1484 ( 
.A(n_667),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_500),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_126),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_631),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_696),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_374),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_907),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_443),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_320),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_852),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_589),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_82),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_905),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_768),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_758),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_868),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_683),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_837),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_747),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_813),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_825),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_928),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_260),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_397),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_57),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_16),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_823),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_832),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_37),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_703),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_679),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_307),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_105),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_826),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_58),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_198),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_439),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_413),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_480),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_564),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_713),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_638),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_349),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_266),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_602),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_383),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_699),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_873),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_700),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_889),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_842),
.Y(n_1534)
);

CKINVDCx14_ASAP7_75t_R g1535 ( 
.A(n_911),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_889),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1365),
.Y(n_1537)
);

INVxp33_ASAP7_75t_SL g1538 ( 
.A(n_1129),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1372),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1372),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1365),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1420),
.B(n_0),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1049),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1049),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_973),
.B(n_0),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_969),
.B(n_1),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1411),
.Y(n_1547)
);

INVxp33_ASAP7_75t_SL g1548 ( 
.A(n_1160),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1411),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1069),
.B(n_2),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1111),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1178),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_1390),
.Y(n_1553)
);

NOR2xp67_ASAP7_75t_L g1554 ( 
.A(n_988),
.B(n_1),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1364),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1166),
.B(n_2),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1397),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_982),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_988),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1390),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1494),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1361),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1178),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_956),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1276),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1219),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1475),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1535),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_956),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_1276),
.Y(n_1570)
);

CKINVDCx16_ASAP7_75t_R g1571 ( 
.A(n_985),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1110),
.B(n_2),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_963),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_1303),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_965),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1535),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1212),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_974),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_962),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_1303),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_1346),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1212),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_980),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1052),
.B(n_3),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1035),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1035),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1003),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_962),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1007),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1353),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_977),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1008),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_962),
.Y(n_1593)
);

INVxp33_ASAP7_75t_SL g1594 ( 
.A(n_1271),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1064),
.B(n_4),
.Y(n_1595)
);

CKINVDCx16_ASAP7_75t_R g1596 ( 
.A(n_1138),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_1346),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1353),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1172),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1357),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1017),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1331),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1149),
.B(n_1158),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_943),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1357),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1024),
.Y(n_1606)
);

NOR2xp67_ASAP7_75t_L g1607 ( 
.A(n_1193),
.B(n_1371),
.Y(n_1607)
);

INVxp67_ASAP7_75t_SL g1608 ( 
.A(n_972),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1030),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1038),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1039),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1042),
.Y(n_1612)
);

CKINVDCx20_ASAP7_75t_R g1613 ( 
.A(n_1414),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_946),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1414),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1533),
.B(n_3),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1048),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_1417),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1417),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1426),
.Y(n_1620)
);

INVxp67_ASAP7_75t_SL g1621 ( 
.A(n_972),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_947),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1051),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_949),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_954),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1057),
.Y(n_1626)
);

INVxp33_ASAP7_75t_L g1627 ( 
.A(n_1313),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1060),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1212),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_955),
.Y(n_1630)
);

INVxp67_ASAP7_75t_L g1631 ( 
.A(n_1223),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1065),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1479),
.B(n_4),
.Y(n_1633)
);

NOR2xp67_ASAP7_75t_L g1634 ( 
.A(n_1461),
.B(n_5),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_960),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1426),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1445),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_981),
.Y(n_1638)
);

CKINVDCx20_ASAP7_75t_R g1639 ( 
.A(n_1445),
.Y(n_1639)
);

CKINVDCx20_ASAP7_75t_R g1640 ( 
.A(n_941),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_961),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1071),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_966),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1072),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_968),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1223),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_962),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1082),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1086),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_981),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1094),
.Y(n_1651)
);

CKINVDCx20_ASAP7_75t_R g1652 ( 
.A(n_942),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_971),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1101),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_976),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1112),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_979),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1279),
.B(n_5),
.Y(n_1658)
);

INVxp33_ASAP7_75t_SL g1659 ( 
.A(n_983),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1223),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_984),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1113),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1118),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_987),
.Y(n_1664)
);

CKINVDCx14_ASAP7_75t_R g1665 ( 
.A(n_1306),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1122),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_989),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1159),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1569),
.B(n_1063),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1638),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1591),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1558),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1563),
.B(n_990),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1638),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1650),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1665),
.B(n_1306),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1559),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1539),
.Y(n_1678)
);

OAI22x1_ASAP7_75t_SL g1679 ( 
.A1(n_1640),
.A2(n_1067),
.B1(n_1077),
.B2(n_986),
.Y(n_1679)
);

INVx6_ASAP7_75t_L g1680 ( 
.A(n_1550),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1551),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1579),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1571),
.A2(n_994),
.B1(n_995),
.B2(n_991),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1588),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1593),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1563),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1647),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1540),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1537),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1555),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1591),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1547),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1549),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1608),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1621),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1629),
.B(n_999),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1604),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1614),
.Y(n_1698)
);

AND2x6_ASAP7_75t_L g1699 ( 
.A(n_1577),
.B(n_1089),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1557),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1561),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1631),
.B(n_1001),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1646),
.B(n_1005),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1627),
.B(n_1306),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1633),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1582),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1573),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1660),
.B(n_1538),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1575),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1578),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1583),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1587),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1589),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1592),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1591),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1601),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1606),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1609),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1610),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1611),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1612),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1617),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1623),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1626),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1628),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1622),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1596),
.B(n_1359),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1632),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1642),
.Y(n_1729)
);

AND2x6_ASAP7_75t_L g1730 ( 
.A(n_1566),
.B(n_1089),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1644),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1648),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1649),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1624),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1651),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1654),
.A2(n_1047),
.B(n_1012),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1656),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1548),
.B(n_1009),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1562),
.B(n_982),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_SL g1740 ( 
.A(n_1659),
.B(n_1359),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1662),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1541),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1594),
.A2(n_1603),
.B1(n_1543),
.B2(n_1552),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1564),
.B(n_1196),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1663),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1666),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1568),
.B(n_1356),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1668),
.Y(n_1748)
);

INVx6_ASAP7_75t_L g1749 ( 
.A(n_1591),
.Y(n_1749)
);

INVx6_ASAP7_75t_L g1750 ( 
.A(n_1595),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1554),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1544),
.B(n_1010),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1567),
.B(n_1173),
.Y(n_1753)
);

BUFx8_ASAP7_75t_L g1754 ( 
.A(n_1553),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1584),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1584),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1607),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1658),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1658),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1556),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1556),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1625),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1630),
.B(n_1359),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_1635),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1641),
.B(n_1482),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1643),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1634),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1576),
.B(n_1014),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1545),
.B(n_1103),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1667),
.B(n_1173),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1645),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1546),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1572),
.B(n_1103),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1653),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1616),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_L g1776 ( 
.A(n_1655),
.B(n_1173),
.Y(n_1776)
);

NAND2xp33_ASAP7_75t_L g1777 ( 
.A(n_1657),
.B(n_1173),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1542),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1661),
.B(n_1015),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1664),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1599),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1602),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1585),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1586),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1590),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1598),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1560),
.B(n_1482),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1652),
.B(n_1407),
.Y(n_1788)
);

BUFx3_ASAP7_75t_L g1789 ( 
.A(n_1565),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1570),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1574),
.B(n_1135),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1580),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1581),
.Y(n_1793)
);

CKINVDCx11_ASAP7_75t_R g1794 ( 
.A(n_1597),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1600),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1605),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1613),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1615),
.B(n_1173),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1618),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1619),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1620),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1636),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1637),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1639),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1638),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1558),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1558),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1638),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1563),
.B(n_1016),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1665),
.B(n_1482),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1558),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1665),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1638),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1665),
.B(n_1104),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1638),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1665),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1563),
.B(n_1135),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1665),
.B(n_1104),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1577),
.B(n_1173),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1638),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1577),
.B(n_1173),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1558),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1591),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1665),
.B(n_1119),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1558),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1650),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1638),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1638),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1638),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1558),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1558),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1638),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1569),
.B(n_1334),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1563),
.B(n_1151),
.Y(n_1834)
);

AND2x2_ASAP7_75t_SL g1835 ( 
.A(n_1571),
.B(n_944),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1558),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1665),
.B(n_1119),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1591),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1558),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1638),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1638),
.Y(n_1841)
);

AND2x2_ASAP7_75t_SL g1842 ( 
.A(n_1571),
.B(n_944),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1558),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1569),
.B(n_1019),
.Y(n_1844)
);

OAI21x1_ASAP7_75t_L g1845 ( 
.A1(n_1579),
.A2(n_1047),
.B(n_1012),
.Y(n_1845)
);

BUFx6f_ASAP7_75t_L g1846 ( 
.A(n_1591),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1563),
.B(n_1151),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1591),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1569),
.B(n_1022),
.Y(n_1849)
);

AND3x2_ASAP7_75t_L g1850 ( 
.A(n_1563),
.B(n_1130),
.C(n_1391),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1558),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1638),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1638),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1638),
.Y(n_1854)
);

BUFx6f_ASAP7_75t_L g1855 ( 
.A(n_1591),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1638),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1591),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1638),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1638),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1638),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1665),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1638),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1558),
.Y(n_1863)
);

BUFx2_ASAP7_75t_L g1864 ( 
.A(n_1563),
.Y(n_1864)
);

INVx3_ASAP7_75t_L g1865 ( 
.A(n_1558),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1638),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1577),
.B(n_962),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1665),
.B(n_1126),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1665),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1591),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1665),
.Y(n_1871)
);

OAI21x1_ASAP7_75t_L g1872 ( 
.A1(n_1579),
.A2(n_1132),
.B(n_1075),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1563),
.B(n_1029),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1558),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1558),
.Y(n_1875)
);

BUFx6f_ASAP7_75t_L g1876 ( 
.A(n_1591),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1577),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1577),
.B(n_962),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1558),
.Y(n_1879)
);

CKINVDCx6p67_ASAP7_75t_R g1880 ( 
.A(n_1571),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1571),
.A2(n_1031),
.B1(n_1036),
.B2(n_1032),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1638),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1558),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1558),
.Y(n_1884)
);

OR2x6_ASAP7_75t_L g1885 ( 
.A(n_1812),
.B(n_1248),
.Y(n_1885)
);

OR2x2_ASAP7_75t_SL g1886 ( 
.A(n_1816),
.B(n_1025),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1760),
.A2(n_1761),
.B1(n_1705),
.B2(n_1778),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1706),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1701),
.Y(n_1889)
);

INVx4_ASAP7_75t_SL g1890 ( 
.A(n_1730),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1845),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1690),
.Y(n_1892)
);

INVx3_ASAP7_75t_L g1893 ( 
.A(n_1877),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1872),
.Y(n_1894)
);

OR2x6_ASAP7_75t_L g1895 ( 
.A(n_1861),
.B(n_1208),
.Y(n_1895)
);

INVxp67_ASAP7_75t_SL g1896 ( 
.A(n_1686),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1736),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1717),
.B(n_1040),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1758),
.A2(n_1126),
.B1(n_1222),
.B2(n_1184),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1736),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1722),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1723),
.Y(n_1902)
);

INVx2_ASAP7_75t_SL g1903 ( 
.A(n_1676),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1672),
.Y(n_1904)
);

INVx3_ASAP7_75t_L g1905 ( 
.A(n_1806),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1741),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1700),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1822),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1794),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1810),
.B(n_1075),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1769),
.B(n_1041),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1825),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1769),
.B(n_1044),
.Y(n_1913)
);

CKINVDCx11_ASAP7_75t_R g1914 ( 
.A(n_1880),
.Y(n_1914)
);

OR2x6_ASAP7_75t_L g1915 ( 
.A(n_1869),
.B(n_1107),
.Y(n_1915)
);

OR2x6_ASAP7_75t_L g1916 ( 
.A(n_1871),
.B(n_1157),
.Y(n_1916)
);

OR2x6_ASAP7_75t_L g1917 ( 
.A(n_1697),
.B(n_1232),
.Y(n_1917)
);

INVx3_ASAP7_75t_L g1918 ( 
.A(n_1807),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1830),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1678),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1864),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1755),
.B(n_1050),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1688),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1704),
.B(n_1864),
.Y(n_1924)
);

AOI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1680),
.A2(n_1056),
.B1(n_1059),
.B2(n_1055),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1756),
.B(n_1066),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1692),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1680),
.A2(n_1074),
.B1(n_1076),
.B2(n_1070),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1693),
.Y(n_1929)
);

OA22x2_ASAP7_75t_L g1930 ( 
.A1(n_1791),
.A2(n_1850),
.B1(n_1743),
.B2(n_1800),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1694),
.Y(n_1931)
);

NOR3xp33_ASAP7_75t_L g1932 ( 
.A(n_1708),
.B(n_1484),
.C(n_1109),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1695),
.B(n_1759),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1759),
.B(n_1132),
.Y(n_1934)
);

OAI21xp33_ASAP7_75t_SL g1935 ( 
.A1(n_1772),
.A2(n_1176),
.B(n_1169),
.Y(n_1935)
);

AOI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1740),
.A2(n_1093),
.B1(n_1096),
.B2(n_1081),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1814),
.B(n_1150),
.Y(n_1937)
);

INVx2_ASAP7_75t_SL g1938 ( 
.A(n_1818),
.Y(n_1938)
);

INVx6_ASAP7_75t_L g1939 ( 
.A(n_1764),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1831),
.Y(n_1940)
);

INVx4_ASAP7_75t_L g1941 ( 
.A(n_1730),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1836),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1727),
.B(n_950),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1824),
.B(n_1097),
.Y(n_1944)
);

INVx5_ASAP7_75t_L g1945 ( 
.A(n_1730),
.Y(n_1945)
);

OR2x6_ASAP7_75t_L g1946 ( 
.A(n_1697),
.B(n_1256),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1677),
.Y(n_1947)
);

INVx5_ASAP7_75t_L g1948 ( 
.A(n_1782),
.Y(n_1948)
);

AND2x6_ASAP7_75t_L g1949 ( 
.A(n_1837),
.B(n_1184),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1839),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1681),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1868),
.B(n_1098),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1843),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1851),
.Y(n_1954)
);

AND2x6_ASAP7_75t_L g1955 ( 
.A(n_1763),
.B(n_1222),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1811),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1707),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1709),
.Y(n_1958)
);

NAND3xp33_ASAP7_75t_L g1959 ( 
.A(n_1738),
.B(n_1114),
.C(n_1108),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1863),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1874),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1712),
.Y(n_1962)
);

BUFx10_ASAP7_75t_L g1963 ( 
.A(n_1742),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1775),
.A2(n_1450),
.B1(n_1478),
.B2(n_1332),
.Y(n_1964)
);

AO22x2_ASAP7_75t_L g1965 ( 
.A1(n_1791),
.A2(n_1125),
.B1(n_1128),
.B2(n_1020),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_SL g1966 ( 
.A(n_1779),
.B(n_1150),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1713),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1765),
.B(n_1174),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1673),
.B(n_1116),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1875),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1879),
.Y(n_1971)
);

OR2x6_ASAP7_75t_L g1972 ( 
.A(n_1726),
.B(n_1266),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1883),
.Y(n_1973)
);

INVx2_ASAP7_75t_SL g1974 ( 
.A(n_1826),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1670),
.A2(n_1121),
.B1(n_1124),
.B2(n_1117),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1696),
.B(n_1174),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1721),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1729),
.Y(n_1978)
);

CKINVDCx20_ASAP7_75t_R g1979 ( 
.A(n_1726),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1731),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1689),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1865),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1733),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1884),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1745),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1809),
.B(n_1134),
.Y(n_1986)
);

NAND3xp33_ASAP7_75t_L g1987 ( 
.A(n_1833),
.B(n_1849),
.C(n_1844),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1873),
.B(n_1136),
.Y(n_1988)
);

INVx2_ASAP7_75t_SL g1989 ( 
.A(n_1750),
.Y(n_1989)
);

INVx4_ASAP7_75t_L g1990 ( 
.A(n_1699),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1710),
.B(n_1137),
.Y(n_1991)
);

INVx1_ASAP7_75t_SL g1992 ( 
.A(n_1750),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1674),
.A2(n_1450),
.B1(n_1478),
.B2(n_1332),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1751),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1702),
.B(n_1228),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1805),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1762),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1711),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1703),
.B(n_1140),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1808),
.Y(n_2000)
);

AO21x2_ASAP7_75t_L g2001 ( 
.A1(n_1770),
.A2(n_1187),
.B(n_1179),
.Y(n_2001)
);

OAI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1762),
.A2(n_1477),
.B1(n_1520),
.B2(n_1282),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1714),
.B(n_1141),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1716),
.B(n_1142),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1718),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1813),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1815),
.Y(n_2007)
);

INVx2_ASAP7_75t_SL g2008 ( 
.A(n_1817),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1683),
.B(n_1881),
.Y(n_2009)
);

INVxp67_ASAP7_75t_L g2010 ( 
.A(n_1698),
.Y(n_2010)
);

NAND2xp33_ASAP7_75t_SL g2011 ( 
.A(n_1764),
.B(n_1144),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1752),
.B(n_1228),
.Y(n_2012)
);

AND2x6_ASAP7_75t_L g2013 ( 
.A(n_1780),
.B(n_1766),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_SL g2014 ( 
.A(n_1734),
.B(n_1025),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1768),
.B(n_1146),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1820),
.B(n_1148),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_1827),
.B(n_1156),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1828),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1719),
.Y(n_2019)
);

BUFx2_ASAP7_75t_L g2020 ( 
.A(n_1774),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1829),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1832),
.Y(n_2022)
);

XOR2xp5_ASAP7_75t_R g2023 ( 
.A(n_1679),
.B(n_5),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1840),
.Y(n_2024)
);

BUFx4f_ASAP7_75t_L g2025 ( 
.A(n_1782),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1720),
.B(n_1162),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1766),
.B(n_1028),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1841),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1724),
.B(n_1725),
.Y(n_2029)
);

INVxp67_ASAP7_75t_L g2030 ( 
.A(n_1787),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1852),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1754),
.Y(n_2032)
);

INVx2_ASAP7_75t_SL g2033 ( 
.A(n_1817),
.Y(n_2033)
);

OAI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_1853),
.A2(n_1028),
.B1(n_1168),
.B2(n_1165),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1771),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_1799),
.B(n_1143),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1728),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1854),
.Y(n_2038)
);

INVx4_ASAP7_75t_L g2039 ( 
.A(n_1699),
.Y(n_2039)
);

INVxp67_ASAP7_75t_SL g2040 ( 
.A(n_1834),
.Y(n_2040)
);

INVx3_ASAP7_75t_L g2041 ( 
.A(n_1739),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1856),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1732),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1735),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1858),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1737),
.B(n_1175),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_1859),
.A2(n_1182),
.B1(n_1186),
.B2(n_1177),
.Y(n_2047)
);

NAND3xp33_ASAP7_75t_L g2048 ( 
.A(n_1860),
.B(n_1194),
.C(n_1192),
.Y(n_2048)
);

OR2x6_ASAP7_75t_L g2049 ( 
.A(n_1789),
.B(n_953),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1746),
.B(n_1195),
.Y(n_2050)
);

INVx3_ASAP7_75t_L g2051 ( 
.A(n_1739),
.Y(n_2051)
);

INVxp33_ASAP7_75t_L g2052 ( 
.A(n_1788),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1862),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1748),
.B(n_1199),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1866),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1682),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1682),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1834),
.B(n_1202),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1882),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1847),
.B(n_1205),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1847),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1675),
.A2(n_1842),
.B1(n_1835),
.B2(n_1798),
.Y(n_2062)
);

AND2x6_ASAP7_75t_L g2063 ( 
.A(n_1771),
.B(n_1245),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1773),
.B(n_1206),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1767),
.Y(n_2065)
);

INVxp33_ASAP7_75t_L g2066 ( 
.A(n_1803),
.Y(n_2066)
);

BUFx10_ASAP7_75t_L g2067 ( 
.A(n_1786),
.Y(n_2067)
);

AO22x2_ASAP7_75t_L g2068 ( 
.A1(n_1797),
.A2(n_1216),
.B1(n_1381),
.B2(n_1188),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1684),
.Y(n_2069)
);

INVx2_ASAP7_75t_SL g2070 ( 
.A(n_1699),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1773),
.Y(n_2071)
);

BUFx4f_ASAP7_75t_L g2072 ( 
.A(n_1786),
.Y(n_2072)
);

INVx2_ASAP7_75t_SL g2073 ( 
.A(n_1757),
.Y(n_2073)
);

AND2x6_ASAP7_75t_L g2074 ( 
.A(n_1781),
.B(n_1245),
.Y(n_2074)
);

BUFx2_ASAP7_75t_L g2075 ( 
.A(n_1801),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1684),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1819),
.B(n_1821),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1753),
.Y(n_2078)
);

NAND2xp33_ASAP7_75t_SL g2079 ( 
.A(n_1783),
.B(n_1209),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1867),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1878),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1685),
.Y(n_2082)
);

OR2x6_ASAP7_75t_L g2083 ( 
.A(n_1792),
.B(n_953),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1685),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1687),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1669),
.B(n_1217),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1687),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_1776),
.A2(n_1201),
.B1(n_1213),
.B2(n_1191),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1749),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1749),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1671),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1744),
.B(n_950),
.Y(n_2092)
);

INVx1_ASAP7_75t_SL g2093 ( 
.A(n_1801),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1747),
.B(n_1249),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1777),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1671),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1784),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1691),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1691),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_L g2100 ( 
.A(n_1785),
.B(n_1218),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1715),
.Y(n_2101)
);

AND2x6_ASAP7_75t_L g2102 ( 
.A(n_1793),
.B(n_1249),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_1797),
.A2(n_1227),
.B1(n_1230),
.B2(n_1220),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_1715),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1823),
.Y(n_2105)
);

NAND3xp33_ASAP7_75t_L g2106 ( 
.A(n_1800),
.B(n_1229),
.C(n_1225),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1823),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1838),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1838),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1802),
.B(n_1259),
.Y(n_2110)
);

INVxp67_ASAP7_75t_L g2111 ( 
.A(n_1790),
.Y(n_2111)
);

AOI22xp33_ASAP7_75t_L g2112 ( 
.A1(n_1802),
.A2(n_1241),
.B1(n_1250),
.B2(n_1234),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1795),
.B(n_1236),
.Y(n_2113)
);

AOI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_1796),
.A2(n_1239),
.B1(n_1240),
.B2(n_1238),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1846),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_1804),
.B(n_948),
.Y(n_2116)
);

NAND2xp33_ASAP7_75t_L g2117 ( 
.A(n_1846),
.B(n_962),
.Y(n_2117)
);

NAND2xp33_ASAP7_75t_SL g2118 ( 
.A(n_1848),
.B(n_1523),
.Y(n_2118)
);

INVxp67_ASAP7_75t_SL g2119 ( 
.A(n_1754),
.Y(n_2119)
);

BUFx6f_ASAP7_75t_L g2120 ( 
.A(n_1848),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1855),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1855),
.B(n_1526),
.Y(n_2122)
);

INVxp67_ASAP7_75t_SL g2123 ( 
.A(n_1857),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1857),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1870),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_1870),
.B(n_1259),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_1876),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1876),
.Y(n_2128)
);

NOR2xp33_ASAP7_75t_L g2129 ( 
.A(n_1705),
.B(n_1242),
.Y(n_2129)
);

BUFx4f_ASAP7_75t_L g2130 ( 
.A(n_1880),
.Y(n_2130)
);

BUFx6f_ASAP7_75t_L g2131 ( 
.A(n_1736),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_1736),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1705),
.B(n_1527),
.Y(n_2133)
);

BUFx2_ASAP7_75t_L g2134 ( 
.A(n_1877),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1845),
.Y(n_2135)
);

INVx2_ASAP7_75t_SL g2136 ( 
.A(n_1676),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_1697),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1845),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1845),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1736),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1877),
.B(n_950),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1701),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_1877),
.B(n_967),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_1697),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1701),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1845),
.Y(n_2146)
);

BUFx10_ASAP7_75t_L g2147 ( 
.A(n_1742),
.Y(n_2147)
);

BUFx2_ASAP7_75t_L g2148 ( 
.A(n_1877),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1845),
.Y(n_2149)
);

INVx5_ASAP7_75t_L g2150 ( 
.A(n_1730),
.Y(n_2150)
);

INVx4_ASAP7_75t_L g2151 ( 
.A(n_1706),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_1676),
.B(n_1301),
.Y(n_2152)
);

INVx5_ASAP7_75t_L g2153 ( 
.A(n_1690),
.Y(n_2153)
);

INVx5_ASAP7_75t_L g2154 ( 
.A(n_1690),
.Y(n_2154)
);

BUFx10_ASAP7_75t_L g2155 ( 
.A(n_1742),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1705),
.B(n_1243),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1736),
.Y(n_2157)
);

INVx2_ASAP7_75t_SL g2158 ( 
.A(n_1676),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1845),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1705),
.B(n_1244),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_SL g2161 ( 
.A(n_1676),
.B(n_1301),
.Y(n_2161)
);

INVxp67_ASAP7_75t_L g2162 ( 
.A(n_1877),
.Y(n_2162)
);

BUFx3_ASAP7_75t_L g2163 ( 
.A(n_1697),
.Y(n_2163)
);

NAND3xp33_ASAP7_75t_L g2164 ( 
.A(n_1738),
.B(n_1253),
.C(n_1246),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1676),
.B(n_1389),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1705),
.B(n_1254),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1845),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1705),
.B(n_1516),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1676),
.B(n_1389),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1701),
.Y(n_2170)
);

BUFx3_ASAP7_75t_L g2171 ( 
.A(n_1697),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1701),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1845),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1705),
.B(n_1519),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1845),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_1736),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1701),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1845),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1705),
.B(n_1522),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1705),
.B(n_1529),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1701),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1845),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2129),
.B(n_1255),
.Y(n_2183)
);

AOI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_1924),
.A2(n_2162),
.B1(n_1896),
.B2(n_1932),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1887),
.B(n_1261),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1947),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_2052),
.B(n_1943),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_1893),
.B(n_1280),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_1914),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2056),
.Y(n_2190)
);

AOI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2134),
.A2(n_1272),
.B1(n_1289),
.B2(n_1268),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_1903),
.B(n_1292),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_2148),
.B(n_1350),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2133),
.B(n_1293),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1931),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_2097),
.B(n_957),
.Y(n_2196)
);

NAND2xp33_ASAP7_75t_L g2197 ( 
.A(n_2131),
.B(n_1296),
.Y(n_2197)
);

NAND2xp33_ASAP7_75t_L g2198 ( 
.A(n_2131),
.B(n_1308),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1933),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2156),
.B(n_1515),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1945),
.B(n_1326),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2057),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1945),
.B(n_1347),
.Y(n_2203)
);

BUFx12f_ASAP7_75t_L g2204 ( 
.A(n_2032),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2160),
.B(n_1295),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2166),
.B(n_1299),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1907),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2029),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_1945),
.B(n_1320),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2168),
.B(n_1316),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2069),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_2136),
.B(n_2158),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_1996),
.B(n_959),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2000),
.B(n_996),
.Y(n_2214)
);

BUFx3_ASAP7_75t_L g2215 ( 
.A(n_2130),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2174),
.B(n_1323),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2076),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2082),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_2087),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1998),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_2006),
.B(n_1004),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2005),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2179),
.B(n_1336),
.Y(n_2223)
);

BUFx5_ASAP7_75t_L g2224 ( 
.A(n_2084),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2019),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1897),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2137),
.B(n_1045),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2180),
.B(n_1337),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_2150),
.B(n_1351),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2007),
.B(n_1339),
.Y(n_2230)
);

INVxp67_ASAP7_75t_L g2231 ( 
.A(n_1997),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1900),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2018),
.B(n_1342),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_SL g2234 ( 
.A(n_2150),
.B(n_1355),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2021),
.B(n_1344),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2022),
.B(n_1362),
.Y(n_2236)
);

INVx2_ASAP7_75t_SL g2237 ( 
.A(n_2144),
.Y(n_2237)
);

INVxp67_ASAP7_75t_L g2238 ( 
.A(n_2163),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_1987),
.B(n_1363),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2037),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2043),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_2132),
.Y(n_2242)
);

NOR2xp67_ASAP7_75t_L g2243 ( 
.A(n_2010),
.B(n_1948),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2132),
.Y(n_2244)
);

O2A1O1Ixp33_ASAP7_75t_L g2245 ( 
.A1(n_1935),
.A2(n_1452),
.B(n_1455),
.C(n_1404),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_2030),
.B(n_1369),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2140),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2024),
.B(n_1380),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2028),
.B(n_2031),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2044),
.Y(n_2250)
);

INVx8_ASAP7_75t_L g2251 ( 
.A(n_1895),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2038),
.B(n_1383),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2140),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2061),
.Y(n_2254)
);

AOI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2040),
.A2(n_1392),
.B1(n_1393),
.B2(n_1388),
.Y(n_2255)
);

NAND2xp33_ASAP7_75t_L g2256 ( 
.A(n_2157),
.B(n_1424),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2042),
.B(n_1396),
.Y(n_2257)
);

INVxp67_ASAP7_75t_L g2258 ( 
.A(n_2171),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_2151),
.B(n_1408),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_2150),
.B(n_1416),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_1969),
.A2(n_1410),
.B1(n_1419),
.B2(n_1409),
.Y(n_2261)
);

AOI22xp33_ASAP7_75t_L g2262 ( 
.A1(n_1922),
.A2(n_1422),
.B1(n_1504),
.B2(n_1300),
.Y(n_2262)
);

AOI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_1988),
.A2(n_1427),
.B1(n_1432),
.B2(n_1421),
.Y(n_2263)
);

BUFx3_ASAP7_75t_L g2264 ( 
.A(n_1948),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2045),
.B(n_1434),
.Y(n_2265)
);

NAND2xp33_ASAP7_75t_L g2266 ( 
.A(n_2157),
.B(n_2176),
.Y(n_2266)
);

NAND3xp33_ASAP7_75t_L g2267 ( 
.A(n_2015),
.B(n_1438),
.C(n_1437),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_1921),
.B(n_1045),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2053),
.B(n_1439),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_1992),
.B(n_1443),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2055),
.B(n_1444),
.Y(n_2271)
);

OAI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2059),
.A2(n_1037),
.B1(n_1073),
.B2(n_1033),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_1999),
.B(n_1456),
.Y(n_2273)
);

BUFx3_ASAP7_75t_L g2274 ( 
.A(n_2067),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_1921),
.B(n_1457),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1926),
.B(n_1463),
.Y(n_2276)
);

OAI22xp33_ASAP7_75t_L g2277 ( 
.A1(n_2014),
.A2(n_1946),
.B1(n_1972),
.B2(n_1917),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2176),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1986),
.B(n_1466),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1911),
.B(n_1467),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_1913),
.B(n_1469),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1889),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2085),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_1991),
.B(n_1470),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2003),
.B(n_1472),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2004),
.B(n_1481),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2142),
.Y(n_2287)
);

INVxp67_ASAP7_75t_L g2288 ( 
.A(n_2020),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2026),
.B(n_1483),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2145),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2170),
.Y(n_2291)
);

A2O1A1Ixp33_ASAP7_75t_L g2292 ( 
.A1(n_2016),
.A2(n_1422),
.B(n_1504),
.C(n_1300),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2046),
.B(n_1489),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_1941),
.B(n_1491),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2050),
.B(n_1495),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2054),
.B(n_1506),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1908),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2172),
.B(n_1508),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_1888),
.B(n_1509),
.Y(n_2299)
);

AOI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2062),
.A2(n_951),
.B1(n_952),
.B2(n_940),
.Y(n_2300)
);

NAND2xp33_ASAP7_75t_L g2301 ( 
.A(n_1949),
.B(n_1034),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_R g2302 ( 
.A(n_1979),
.B(n_1139),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_1912),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_R g2304 ( 
.A(n_1909),
.B(n_1147),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2086),
.B(n_1115),
.Y(n_2305)
);

BUFx3_ASAP7_75t_L g2306 ( 
.A(n_1939),
.Y(n_2306)
);

NAND2xp33_ASAP7_75t_L g2307 ( 
.A(n_1949),
.B(n_1034),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2177),
.B(n_2181),
.Y(n_2308)
);

BUFx4_ASAP7_75t_L g2309 ( 
.A(n_1917),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_1890),
.B(n_964),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2017),
.B(n_1270),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2064),
.B(n_1273),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_2104),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1955),
.B(n_1275),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_1890),
.B(n_970),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1955),
.B(n_1277),
.Y(n_2316)
);

AOI22xp33_ASAP7_75t_L g2317 ( 
.A1(n_2071),
.A2(n_1284),
.B1(n_1290),
.B2(n_1278),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1919),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_2153),
.B(n_975),
.Y(n_2319)
);

INVxp67_ASAP7_75t_L g2320 ( 
.A(n_2143),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1955),
.B(n_1518),
.Y(n_2321)
);

NOR3xp33_ASAP7_75t_L g2322 ( 
.A(n_2002),
.B(n_2034),
.C(n_2009),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1957),
.B(n_1521),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1958),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1962),
.B(n_1525),
.Y(n_2325)
);

BUFx2_ASAP7_75t_L g2326 ( 
.A(n_1946),
.Y(n_2326)
);

INVx2_ASAP7_75t_SL g2327 ( 
.A(n_1895),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1967),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_1977),
.B(n_1528),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1978),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_L g2331 ( 
.A(n_1989),
.B(n_1968),
.Y(n_2331)
);

AND2x6_ASAP7_75t_L g2332 ( 
.A(n_2095),
.B(n_1512),
.Y(n_2332)
);

INVxp67_ASAP7_75t_L g2333 ( 
.A(n_1972),
.Y(n_2333)
);

NOR2xp67_ASAP7_75t_SL g2334 ( 
.A(n_1974),
.B(n_978),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1940),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1980),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2008),
.B(n_1197),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1983),
.Y(n_2338)
);

OAI22xp5_ASAP7_75t_SL g2339 ( 
.A1(n_1886),
.A2(n_1235),
.B1(n_1446),
.B2(n_1233),
.Y(n_2339)
);

NAND2x1_ASAP7_75t_L g2340 ( 
.A(n_1990),
.B(n_1231),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_1942),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_2104),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_L g2343 ( 
.A(n_2033),
.B(n_1476),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_1985),
.B(n_1302),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2047),
.B(n_1309),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_1920),
.Y(n_2346)
);

NAND2xp33_ASAP7_75t_SL g2347 ( 
.A(n_2039),
.B(n_1513),
.Y(n_2347)
);

INVx2_ASAP7_75t_SL g2348 ( 
.A(n_2153),
.Y(n_2348)
);

NOR2xp67_ASAP7_75t_L g2349 ( 
.A(n_2106),
.B(n_6),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_2154),
.B(n_992),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1950),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_1953),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_1898),
.B(n_1311),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_2154),
.B(n_993),
.Y(n_2354)
);

NAND2xp33_ASAP7_75t_SL g2355 ( 
.A(n_2070),
.B(n_1517),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_1944),
.B(n_1319),
.Y(n_2356)
);

AOI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_1891),
.A2(n_1512),
.B(n_1324),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2141),
.B(n_997),
.Y(n_2358)
);

INVxp67_ASAP7_75t_SL g2359 ( 
.A(n_2027),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1923),
.Y(n_2360)
);

NOR2xp67_ASAP7_75t_L g2361 ( 
.A(n_1936),
.B(n_6),
.Y(n_2361)
);

NOR2x1p5_ASAP7_75t_L g2362 ( 
.A(n_2119),
.B(n_1531),
.Y(n_2362)
);

NAND2x1_ASAP7_75t_L g2363 ( 
.A(n_2063),
.B(n_977),
.Y(n_2363)
);

INVxp67_ASAP7_75t_L g2364 ( 
.A(n_1915),
.Y(n_2364)
);

AOI22xp5_ASAP7_75t_L g2365 ( 
.A1(n_2060),
.A2(n_1000),
.B1(n_1002),
.B2(n_998),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_1954),
.Y(n_2366)
);

NAND3xp33_ASAP7_75t_L g2367 ( 
.A(n_2100),
.B(n_1013),
.C(n_1011),
.Y(n_2367)
);

AOI21xp5_ASAP7_75t_L g2368 ( 
.A1(n_1894),
.A2(n_1327),
.B(n_1321),
.Y(n_2368)
);

INVx3_ASAP7_75t_L g2369 ( 
.A(n_1960),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_1952),
.B(n_1329),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_1925),
.B(n_1021),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_1965),
.B(n_1045),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_1927),
.B(n_1333),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1929),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2041),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2051),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2058),
.B(n_1345),
.Y(n_2377)
);

INVx4_ASAP7_75t_L g2378 ( 
.A(n_2063),
.Y(n_2378)
);

NAND2xp33_ASAP7_75t_L g2379 ( 
.A(n_1949),
.B(n_1034),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_2066),
.B(n_1026),
.Y(n_2380)
);

HB1xp67_ASAP7_75t_L g2381 ( 
.A(n_1915),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_1934),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_1964),
.B(n_1349),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_1928),
.B(n_1354),
.Y(n_2384)
);

INVx8_ASAP7_75t_L g2385 ( 
.A(n_1885),
.Y(n_2385)
);

AOI22xp33_ASAP7_75t_L g2386 ( 
.A1(n_2074),
.A2(n_2048),
.B1(n_1965),
.B2(n_1959),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2092),
.B(n_1027),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1961),
.Y(n_2388)
);

AOI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_1975),
.A2(n_1046),
.B1(n_1061),
.B2(n_1043),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_1994),
.B(n_1358),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2068),
.B(n_1095),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_1970),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2074),
.B(n_1360),
.Y(n_2393)
);

INVx8_ASAP7_75t_L g2394 ( 
.A(n_1885),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_SL g2395 ( 
.A(n_2088),
.B(n_1078),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_SL g2396 ( 
.A(n_2164),
.B(n_1079),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2074),
.B(n_1377),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_1951),
.B(n_1006),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1901),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2079),
.B(n_1084),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_1902),
.Y(n_2401)
);

NOR2xp33_ASAP7_75t_L g2402 ( 
.A(n_2111),
.B(n_1087),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_1892),
.B(n_1100),
.Y(n_2403)
);

INVxp67_ASAP7_75t_SL g2404 ( 
.A(n_2035),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_1981),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2065),
.B(n_1385),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1899),
.B(n_1398),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_1906),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_1993),
.B(n_1399),
.Y(n_2409)
);

AOI22x1_ASAP7_75t_SL g2410 ( 
.A1(n_2023),
.A2(n_1105),
.B1(n_1106),
.B2(n_1102),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_SL g2411 ( 
.A(n_1938),
.B(n_1120),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1971),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_1910),
.B(n_1123),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_1976),
.B(n_1400),
.Y(n_2414)
);

AOI22xp5_ASAP7_75t_L g2415 ( 
.A1(n_2114),
.A2(n_1133),
.B1(n_1154),
.B2(n_1131),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2068),
.B(n_1095),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_1973),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_1937),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2122),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2110),
.Y(n_2420)
);

INVxp67_ASAP7_75t_L g2421 ( 
.A(n_1916),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_1995),
.B(n_1403),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_SL g2423 ( 
.A(n_2113),
.B(n_1155),
.Y(n_2423)
);

AOI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2152),
.A2(n_2165),
.B1(n_2169),
.B2(n_2161),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2012),
.B(n_1406),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1984),
.Y(n_2426)
);

OR2x2_ASAP7_75t_L g2427 ( 
.A(n_1916),
.B(n_945),
.Y(n_2427)
);

BUFx3_ASAP7_75t_L g2428 ( 
.A(n_1939),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_1966),
.B(n_1429),
.Y(n_2429)
);

NAND2xp33_ASAP7_75t_SL g2430 ( 
.A(n_2036),
.B(n_1524),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2103),
.B(n_1433),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_L g2432 ( 
.A(n_2094),
.B(n_1170),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2073),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_L g2434 ( 
.A(n_1904),
.B(n_1905),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_1963),
.B(n_1095),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_1918),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_1956),
.B(n_1185),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1982),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_2112),
.B(n_1203),
.Y(n_2439)
);

INVx2_ASAP7_75t_SL g2440 ( 
.A(n_2025),
.Y(n_2440)
);

AOI22xp5_ASAP7_75t_L g2441 ( 
.A1(n_1930),
.A2(n_1207),
.B1(n_1210),
.B2(n_1204),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2135),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2013),
.B(n_1435),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_L g2444 ( 
.A(n_2116),
.B(n_1214),
.Y(n_2444)
);

OAI22x1_ASAP7_75t_L g2445 ( 
.A1(n_2023),
.A2(n_1221),
.B1(n_1224),
.B2(n_1215),
.Y(n_2445)
);

CKINVDCx5p33_ASAP7_75t_R g2446 ( 
.A(n_2147),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2013),
.B(n_1436),
.Y(n_2447)
);

INVx3_ASAP7_75t_L g2448 ( 
.A(n_2127),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2083),
.B(n_1237),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2080),
.B(n_1247),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2081),
.B(n_1252),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2078),
.B(n_2011),
.Y(n_2452)
);

INVx2_ASAP7_75t_SL g2453 ( 
.A(n_2072),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_SL g2454 ( 
.A(n_2077),
.B(n_1257),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2138),
.Y(n_2455)
);

BUFx3_ASAP7_75t_L g2456 ( 
.A(n_2075),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2013),
.B(n_1440),
.Y(n_2457)
);

BUFx6f_ASAP7_75t_L g2458 ( 
.A(n_2120),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2139),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2063),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2102),
.B(n_1447),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2102),
.B(n_1448),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2102),
.B(n_1449),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2001),
.B(n_1462),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2146),
.B(n_1464),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_2155),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_2049),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2149),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2159),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_2167),
.B(n_1262),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2173),
.B(n_1465),
.Y(n_2471)
);

OAI22xp5_ASAP7_75t_L g2472 ( 
.A1(n_1886),
.A2(n_1485),
.B1(n_1486),
.B2(n_1480),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2175),
.Y(n_2473)
);

NAND3xp33_ASAP7_75t_L g2474 ( 
.A(n_2083),
.B(n_2049),
.C(n_2118),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2178),
.B(n_1487),
.Y(n_2475)
);

OR2x2_ASAP7_75t_L g2476 ( 
.A(n_2093),
.B(n_958),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2182),
.B(n_1492),
.Y(n_2477)
);

NAND2xp33_ASAP7_75t_L g2478 ( 
.A(n_2120),
.B(n_1034),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2126),
.Y(n_2479)
);

OAI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2123),
.A2(n_1018),
.B1(n_1054),
.B2(n_1053),
.Y(n_2480)
);

NOR3xp33_ASAP7_75t_L g2481 ( 
.A(n_2117),
.B(n_1183),
.C(n_1180),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2089),
.B(n_1263),
.Y(n_2482)
);

BUFx4_ASAP7_75t_L g2483 ( 
.A(n_2101),
.Y(n_2483)
);

AOI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_2090),
.A2(n_1281),
.B1(n_1285),
.B2(n_1267),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2107),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2108),
.B(n_1286),
.Y(n_2486)
);

AND2x4_ASAP7_75t_L g2487 ( 
.A(n_2109),
.B(n_1058),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2115),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_2121),
.B(n_1062),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2091),
.B(n_1287),
.Y(n_2490)
);

NOR3xp33_ASAP7_75t_L g2491 ( 
.A(n_2096),
.B(n_1425),
.C(n_1264),
.Y(n_2491)
);

BUFx5_ASAP7_75t_L g2492 ( 
.A(n_2098),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2099),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_L g2494 ( 
.A(n_2105),
.B(n_1288),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2124),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2125),
.B(n_1294),
.Y(n_2496)
);

NAND2x1_ASAP7_75t_L g2497 ( 
.A(n_2128),
.B(n_977),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2129),
.B(n_1297),
.Y(n_2498)
);

NOR2xp67_ASAP7_75t_L g2499 ( 
.A(n_2162),
.B(n_7),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2056),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2129),
.B(n_1298),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_2162),
.B(n_1304),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_1947),
.Y(n_2503)
);

NOR2x1p5_ASAP7_75t_L g2504 ( 
.A(n_2119),
.B(n_1315),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_1947),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2056),
.Y(n_2506)
);

INVx2_ASAP7_75t_SL g2507 ( 
.A(n_2134),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2129),
.B(n_1307),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_2162),
.B(n_1310),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2129),
.B(n_1314),
.Y(n_2510)
);

INVx3_ASAP7_75t_L g2511 ( 
.A(n_1941),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2129),
.B(n_1317),
.Y(n_2512)
);

XOR2xp5_ASAP7_75t_L g2513 ( 
.A(n_2032),
.B(n_1325),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2134),
.B(n_1226),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_2162),
.B(n_1328),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2129),
.B(n_1330),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2056),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2129),
.B(n_1335),
.Y(n_2518)
);

INVx2_ASAP7_75t_SL g2519 ( 
.A(n_2134),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_SL g2520 ( 
.A(n_2162),
.B(n_1338),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_1947),
.Y(n_2521)
);

NOR2xp33_ASAP7_75t_L g2522 ( 
.A(n_2162),
.B(n_1340),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_1947),
.Y(n_2523)
);

AO22x1_ASAP7_75t_L g2524 ( 
.A1(n_2134),
.A2(n_1348),
.B1(n_1352),
.B2(n_1341),
.Y(n_2524)
);

BUFx6f_ASAP7_75t_L g2525 ( 
.A(n_2131),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2129),
.B(n_1366),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2056),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2056),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2162),
.B(n_1367),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2129),
.B(n_1368),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2056),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2056),
.Y(n_2532)
);

BUFx6f_ASAP7_75t_L g2533 ( 
.A(n_2131),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2134),
.B(n_1226),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2162),
.B(n_1374),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2056),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2056),
.Y(n_2537)
);

INVx8_ASAP7_75t_L g2538 ( 
.A(n_1895),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2056),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_1947),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2134),
.B(n_1226),
.Y(n_2541)
);

AOI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_1924),
.A2(n_1375),
.B1(n_1376),
.B2(n_1370),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2129),
.B(n_1378),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2162),
.B(n_1384),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2056),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_1947),
.Y(n_2546)
);

INVx2_ASAP7_75t_SL g2547 ( 
.A(n_2134),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_L g2548 ( 
.A(n_2162),
.B(n_1386),
.Y(n_2548)
);

AOI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_1924),
.A2(n_1395),
.B1(n_1405),
.B2(n_1379),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_L g2550 ( 
.A(n_2162),
.B(n_1412),
.Y(n_2550)
);

OR2x2_ASAP7_75t_L g2551 ( 
.A(n_2134),
.B(n_1458),
.Y(n_2551)
);

INVx2_ASAP7_75t_SL g2552 ( 
.A(n_2134),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_SL g2553 ( 
.A(n_2162),
.B(n_1413),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2056),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_1947),
.Y(n_2555)
);

NOR3xp33_ASAP7_75t_L g2556 ( 
.A(n_2002),
.B(n_1500),
.C(n_1423),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2056),
.Y(n_2557)
);

NAND3xp33_ASAP7_75t_L g2558 ( 
.A(n_2015),
.B(n_1428),
.C(n_1415),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2129),
.B(n_1430),
.Y(n_2559)
);

OR2x2_ASAP7_75t_L g2560 ( 
.A(n_2272),
.B(n_2507),
.Y(n_2560)
);

OAI21xp5_ASAP7_75t_L g2561 ( 
.A1(n_2368),
.A2(n_1083),
.B(n_1068),
.Y(n_2561)
);

OAI21xp5_ASAP7_75t_L g2562 ( 
.A1(n_2357),
.A2(n_1090),
.B(n_1085),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_2519),
.B(n_1505),
.Y(n_2563)
);

INVx4_ASAP7_75t_L g2564 ( 
.A(n_2251),
.Y(n_2564)
);

AO22x1_ASAP7_75t_L g2565 ( 
.A1(n_2309),
.A2(n_1454),
.B1(n_1460),
.B2(n_1453),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_2547),
.B(n_2552),
.Y(n_2566)
);

AOI21xp5_ASAP7_75t_L g2567 ( 
.A1(n_2468),
.A2(n_1092),
.B(n_1091),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2208),
.B(n_1471),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2288),
.B(n_1488),
.Y(n_2569)
);

BUFx2_ASAP7_75t_L g2570 ( 
.A(n_2302),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2249),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2199),
.B(n_1490),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2186),
.B(n_1493),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2469),
.Y(n_2574)
);

BUFx6f_ASAP7_75t_L g2575 ( 
.A(n_2313),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2226),
.Y(n_2576)
);

BUFx6f_ASAP7_75t_L g2577 ( 
.A(n_2313),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2195),
.B(n_1496),
.Y(n_2578)
);

NOR3xp33_ASAP7_75t_L g2579 ( 
.A(n_2277),
.B(n_1514),
.C(n_1499),
.Y(n_2579)
);

AOI21xp5_ASAP7_75t_L g2580 ( 
.A1(n_2442),
.A2(n_1152),
.B(n_1127),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2503),
.B(n_1497),
.Y(n_2581)
);

OAI21xp33_ASAP7_75t_L g2582 ( 
.A1(n_2246),
.A2(n_1501),
.B(n_1498),
.Y(n_2582)
);

AOI22xp5_ASAP7_75t_L g2583 ( 
.A1(n_2322),
.A2(n_1503),
.B1(n_1510),
.B2(n_1502),
.Y(n_2583)
);

BUFx3_ASAP7_75t_L g2584 ( 
.A(n_2274),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2505),
.Y(n_2585)
);

AOI21xp5_ASAP7_75t_L g2586 ( 
.A1(n_2455),
.A2(n_1161),
.B(n_1153),
.Y(n_2586)
);

OAI21xp33_ASAP7_75t_L g2587 ( 
.A1(n_2194),
.A2(n_1511),
.B(n_1164),
.Y(n_2587)
);

BUFx6f_ASAP7_75t_L g2588 ( 
.A(n_2313),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2232),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2521),
.B(n_1163),
.Y(n_2590)
);

AOI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2472),
.A2(n_1171),
.B1(n_1190),
.B2(n_1181),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_SL g2592 ( 
.A(n_2231),
.B(n_977),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2523),
.B(n_1442),
.Y(n_2593)
);

AND2x4_ASAP7_75t_L g2594 ( 
.A(n_2540),
.B(n_1198),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_2305),
.B(n_1468),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2546),
.B(n_1474),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_SL g2597 ( 
.A(n_2430),
.B(n_1023),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2555),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_SL g2599 ( 
.A(n_2224),
.B(n_1023),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2283),
.Y(n_2600)
);

AOI22xp33_ASAP7_75t_L g2601 ( 
.A1(n_2556),
.A2(n_1088),
.B1(n_1145),
.B2(n_1023),
.Y(n_2601)
);

AND2x4_ASAP7_75t_L g2602 ( 
.A(n_2419),
.B(n_1211),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_SL g2603 ( 
.A(n_2224),
.B(n_1023),
.Y(n_2603)
);

AOI21xp5_ASAP7_75t_L g2604 ( 
.A1(n_2459),
.A2(n_1265),
.B(n_1260),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_SL g2605 ( 
.A(n_2224),
.B(n_1088),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2483),
.Y(n_2606)
);

NOR2xp67_ASAP7_75t_SL g2607 ( 
.A(n_2446),
.B(n_1088),
.Y(n_2607)
);

AOI21xp5_ASAP7_75t_L g2608 ( 
.A1(n_2473),
.A2(n_1274),
.B(n_1269),
.Y(n_2608)
);

OR2x6_ASAP7_75t_L g2609 ( 
.A(n_2251),
.B(n_1080),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2207),
.B(n_2239),
.Y(n_2610)
);

AO21x2_ASAP7_75t_L g2611 ( 
.A1(n_2266),
.A2(n_1305),
.B(n_1291),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2317),
.B(n_2345),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2356),
.B(n_1387),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2370),
.B(n_1401),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2311),
.B(n_1402),
.Y(n_2615)
);

INVx11_ASAP7_75t_L g2616 ( 
.A(n_2204),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2391),
.B(n_1418),
.Y(n_2617)
);

AOI22xp5_ASAP7_75t_L g2618 ( 
.A1(n_2361),
.A2(n_1318),
.B1(n_1343),
.B2(n_1322),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2220),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_SL g2620 ( 
.A(n_2224),
.B(n_1088),
.Y(n_2620)
);

BUFx2_ASAP7_75t_L g2621 ( 
.A(n_2238),
.Y(n_2621)
);

AOI21xp5_ASAP7_75t_L g2622 ( 
.A1(n_2465),
.A2(n_1431),
.B(n_1382),
.Y(n_2622)
);

INVx3_ASAP7_75t_L g2623 ( 
.A(n_2378),
.Y(n_2623)
);

AOI21xp5_ASAP7_75t_L g2624 ( 
.A1(n_2471),
.A2(n_2477),
.B(n_2475),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2196),
.B(n_2213),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_SL g2626 ( 
.A(n_2224),
.B(n_1145),
.Y(n_2626)
);

A2O1A1Ixp33_ASAP7_75t_L g2627 ( 
.A1(n_2245),
.A2(n_1532),
.B(n_1536),
.C(n_1530),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2200),
.A2(n_1099),
.B(n_1080),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_SL g2629 ( 
.A(n_2237),
.B(n_1145),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2190),
.Y(n_2630)
);

INVx1_ASAP7_75t_SL g2631 ( 
.A(n_2551),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2196),
.B(n_1099),
.Y(n_2632)
);

AND2x4_ASAP7_75t_L g2633 ( 
.A(n_2327),
.B(n_1167),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2416),
.B(n_1167),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2202),
.Y(n_2635)
);

A2O1A1Ixp33_ASAP7_75t_L g2636 ( 
.A1(n_2292),
.A2(n_1258),
.B(n_1283),
.C(n_1189),
.Y(n_2636)
);

NOR2xp33_ASAP7_75t_L g2637 ( 
.A(n_2187),
.B(n_1189),
.Y(n_2637)
);

AOI21xp5_ASAP7_75t_L g2638 ( 
.A1(n_2205),
.A2(n_1283),
.B(n_1258),
.Y(n_2638)
);

AOI21xp5_ASAP7_75t_L g2639 ( 
.A1(n_2206),
.A2(n_2216),
.B(n_2210),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2213),
.B(n_2214),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2214),
.B(n_1312),
.Y(n_2641)
);

AOI21xp5_ASAP7_75t_L g2642 ( 
.A1(n_2223),
.A2(n_1373),
.B(n_1312),
.Y(n_2642)
);

AOI21xp5_ASAP7_75t_L g2643 ( 
.A1(n_2228),
.A2(n_1373),
.B(n_1251),
.Y(n_2643)
);

AOI21xp5_ASAP7_75t_L g2644 ( 
.A1(n_2284),
.A2(n_1251),
.B(n_1145),
.Y(n_2644)
);

AOI21xp5_ASAP7_75t_L g2645 ( 
.A1(n_2285),
.A2(n_1473),
.B(n_1251),
.Y(n_2645)
);

AOI21xp5_ASAP7_75t_L g2646 ( 
.A1(n_2286),
.A2(n_1473),
.B(n_1251),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2221),
.B(n_1034),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2221),
.B(n_1034),
.Y(n_2648)
);

AOI21xp5_ASAP7_75t_L g2649 ( 
.A1(n_2289),
.A2(n_1507),
.B(n_1473),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2211),
.Y(n_2650)
);

AOI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_2293),
.A2(n_1507),
.B(n_1473),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2222),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2217),
.Y(n_2653)
);

OAI21xp5_ASAP7_75t_L g2654 ( 
.A1(n_2464),
.A2(n_1034),
.B(n_1507),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_2342),
.B(n_1507),
.Y(n_2655)
);

AOI21xp5_ASAP7_75t_L g2656 ( 
.A1(n_2295),
.A2(n_2296),
.B(n_2276),
.Y(n_2656)
);

AND2x2_ASAP7_75t_SL g2657 ( 
.A(n_2326),
.B(n_1394),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2384),
.B(n_7),
.Y(n_2658)
);

CKINVDCx10_ASAP7_75t_R g2659 ( 
.A(n_2189),
.Y(n_2659)
);

BUFx2_ASAP7_75t_L g2660 ( 
.A(n_2258),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2218),
.Y(n_2661)
);

BUFx4f_ASAP7_75t_L g2662 ( 
.A(n_2538),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2219),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2500),
.Y(n_2664)
);

AND2x4_ASAP7_75t_L g2665 ( 
.A(n_2243),
.B(n_7),
.Y(n_2665)
);

INVxp67_ASAP7_75t_L g2666 ( 
.A(n_2476),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2506),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2184),
.B(n_8),
.Y(n_2668)
);

CKINVDCx10_ASAP7_75t_R g2669 ( 
.A(n_2405),
.Y(n_2669)
);

AOI21xp5_ASAP7_75t_L g2670 ( 
.A1(n_2244),
.A2(n_1394),
.B(n_1200),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_SL g2671 ( 
.A(n_2342),
.B(n_1200),
.Y(n_2671)
);

AOI21xp5_ASAP7_75t_L g2672 ( 
.A1(n_2247),
.A2(n_1394),
.B(n_1200),
.Y(n_2672)
);

AOI21xp5_ASAP7_75t_L g2673 ( 
.A1(n_2253),
.A2(n_1394),
.B(n_1200),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2312),
.B(n_8),
.Y(n_2674)
);

CKINVDCx5p33_ASAP7_75t_R g2675 ( 
.A(n_2304),
.Y(n_2675)
);

AOI21xp5_ASAP7_75t_L g2676 ( 
.A1(n_2278),
.A2(n_1451),
.B(n_1441),
.Y(n_2676)
);

AOI21xp5_ASAP7_75t_L g2677 ( 
.A1(n_2308),
.A2(n_1451),
.B(n_1441),
.Y(n_2677)
);

BUFx12f_ASAP7_75t_L g2678 ( 
.A(n_2466),
.Y(n_2678)
);

AOI21xp5_ASAP7_75t_L g2679 ( 
.A1(n_2353),
.A2(n_1451),
.B(n_1441),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_SL g2680 ( 
.A(n_2342),
.B(n_1441),
.Y(n_2680)
);

BUFx2_ASAP7_75t_L g2681 ( 
.A(n_2456),
.Y(n_2681)
);

O2A1O1Ixp33_ASAP7_75t_L g2682 ( 
.A1(n_2372),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_2682)
);

AOI21xp5_ASAP7_75t_L g2683 ( 
.A1(n_2279),
.A2(n_1459),
.B(n_1451),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2377),
.B(n_9),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_SL g2685 ( 
.A(n_2458),
.B(n_1459),
.Y(n_2685)
);

O2A1O1Ixp5_ASAP7_75t_L g2686 ( 
.A1(n_2470),
.A2(n_1534),
.B(n_1459),
.C(n_12),
.Y(n_2686)
);

AOI21x1_ASAP7_75t_L g2687 ( 
.A1(n_2499),
.A2(n_1534),
.B(n_1459),
.Y(n_2687)
);

OAI21xp5_ASAP7_75t_L g2688 ( 
.A1(n_2517),
.A2(n_1534),
.B(n_10),
.Y(n_2688)
);

O2A1O1Ixp5_ASAP7_75t_L g2689 ( 
.A1(n_2314),
.A2(n_2321),
.B(n_2316),
.C(n_2396),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2431),
.B(n_10),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2225),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2240),
.Y(n_2692)
);

AOI21xp33_ASAP7_75t_L g2693 ( 
.A1(n_2270),
.A2(n_1534),
.B(n_11),
.Y(n_2693)
);

HB1xp67_ASAP7_75t_L g2694 ( 
.A(n_2381),
.Y(n_2694)
);

BUFx6f_ASAP7_75t_L g2695 ( 
.A(n_2458),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_SL g2696 ( 
.A(n_2458),
.B(n_12),
.Y(n_2696)
);

AOI22xp33_ASAP7_75t_L g2697 ( 
.A1(n_2339),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2697)
);

AOI21xp5_ASAP7_75t_L g2698 ( 
.A1(n_2230),
.A2(n_13),
.B(n_14),
.Y(n_2698)
);

BUFx3_ASAP7_75t_L g2699 ( 
.A(n_2264),
.Y(n_2699)
);

OR2x6_ASAP7_75t_L g2700 ( 
.A(n_2538),
.B(n_13),
.Y(n_2700)
);

INVx3_ASAP7_75t_L g2701 ( 
.A(n_2378),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2191),
.B(n_14),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2233),
.B(n_15),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2235),
.B(n_15),
.Y(n_2704)
);

OAI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2241),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2250),
.Y(n_2706)
);

AOI21xp5_ASAP7_75t_L g2707 ( 
.A1(n_2236),
.A2(n_17),
.B(n_18),
.Y(n_2707)
);

OAI21xp33_ASAP7_75t_L g2708 ( 
.A1(n_2183),
.A2(n_19),
.B(n_20),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2248),
.B(n_19),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2252),
.B(n_20),
.Y(n_2710)
);

O2A1O1Ixp33_ASAP7_75t_L g2711 ( 
.A1(n_2185),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2527),
.Y(n_2712)
);

AOI21x1_ASAP7_75t_L g2713 ( 
.A1(n_2460),
.A2(n_2397),
.B(n_2393),
.Y(n_2713)
);

INVx2_ASAP7_75t_SL g2714 ( 
.A(n_2385),
.Y(n_2714)
);

AND2x4_ASAP7_75t_L g2715 ( 
.A(n_2215),
.B(n_2433),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2282),
.Y(n_2716)
);

AOI21xp5_ASAP7_75t_L g2717 ( 
.A1(n_2257),
.A2(n_21),
.B(n_22),
.Y(n_2717)
);

AOI21xp5_ASAP7_75t_L g2718 ( 
.A1(n_2265),
.A2(n_21),
.B(n_22),
.Y(n_2718)
);

INVx3_ASAP7_75t_L g2719 ( 
.A(n_2511),
.Y(n_2719)
);

AOI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2269),
.A2(n_2271),
.B(n_2280),
.Y(n_2720)
);

AOI21xp5_ASAP7_75t_L g2721 ( 
.A1(n_2281),
.A2(n_23),
.B(n_24),
.Y(n_2721)
);

AOI21x1_ASAP7_75t_L g2722 ( 
.A1(n_2443),
.A2(n_23),
.B(n_24),
.Y(n_2722)
);

BUFx3_ASAP7_75t_L g2723 ( 
.A(n_2306),
.Y(n_2723)
);

AOI21xp5_ASAP7_75t_L g2724 ( 
.A1(n_2298),
.A2(n_25),
.B(n_26),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2254),
.B(n_25),
.Y(n_2725)
);

NAND2xp33_ASAP7_75t_L g2726 ( 
.A(n_2332),
.B(n_26),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2261),
.B(n_2263),
.Y(n_2727)
);

BUFx6f_ASAP7_75t_L g2728 ( 
.A(n_2242),
.Y(n_2728)
);

NOR2xp33_ASAP7_75t_SL g2729 ( 
.A(n_2385),
.B(n_2394),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2255),
.B(n_2273),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2287),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_SL g2732 ( 
.A(n_2347),
.B(n_27),
.Y(n_2732)
);

A2O1A1Ixp33_ASAP7_75t_L g2733 ( 
.A1(n_2349),
.A2(n_28),
.B(n_25),
.C(n_27),
.Y(n_2733)
);

AND2x4_ASAP7_75t_L g2734 ( 
.A(n_2474),
.B(n_27),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2290),
.B(n_28),
.Y(n_2735)
);

OAI321xp33_ASAP7_75t_L g2736 ( 
.A1(n_2386),
.A2(n_31),
.A3(n_33),
.B1(n_29),
.B2(n_30),
.C(n_32),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_SL g2737 ( 
.A(n_2259),
.B(n_2514),
.Y(n_2737)
);

AOI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2423),
.A2(n_29),
.B(n_30),
.Y(n_2738)
);

AOI22xp5_ASAP7_75t_L g2739 ( 
.A1(n_2332),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_2739)
);

NAND2xp33_ASAP7_75t_L g2740 ( 
.A(n_2332),
.B(n_34),
.Y(n_2740)
);

A2O1A1Ixp33_ASAP7_75t_L g2741 ( 
.A1(n_2267),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_2741)
);

OAI321xp33_ASAP7_75t_L g2742 ( 
.A1(n_2262),
.A2(n_36),
.A3(n_38),
.B1(n_33),
.B2(n_35),
.C(n_37),
.Y(n_2742)
);

INVx3_ASAP7_75t_L g2743 ( 
.A(n_2511),
.Y(n_2743)
);

AOI21xp5_ASAP7_75t_L g2744 ( 
.A1(n_2528),
.A2(n_35),
.B(n_38),
.Y(n_2744)
);

OAI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_2531),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_2745)
);

OAI21xp5_ASAP7_75t_L g2746 ( 
.A1(n_2532),
.A2(n_39),
.B(n_40),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_SL g2747 ( 
.A(n_2534),
.B(n_40),
.Y(n_2747)
);

OAI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2536),
.A2(n_2554),
.B(n_2545),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2291),
.B(n_39),
.Y(n_2749)
);

BUFx3_ASAP7_75t_L g2750 ( 
.A(n_2428),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2537),
.A2(n_41),
.B(n_42),
.Y(n_2751)
);

AOI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2332),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2752)
);

AO21x1_ASAP7_75t_L g2753 ( 
.A1(n_2301),
.A2(n_671),
.B(n_670),
.Y(n_2753)
);

A2O1A1Ixp33_ASAP7_75t_L g2754 ( 
.A1(n_2539),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2324),
.B(n_43),
.Y(n_2755)
);

BUFx6f_ASAP7_75t_L g2756 ( 
.A(n_2242),
.Y(n_2756)
);

AOI21xp5_ASAP7_75t_L g2757 ( 
.A1(n_2557),
.A2(n_44),
.B(n_45),
.Y(n_2757)
);

AOI21xp5_ASAP7_75t_L g2758 ( 
.A1(n_2242),
.A2(n_44),
.B(n_45),
.Y(n_2758)
);

OAI21xp5_ASAP7_75t_L g2759 ( 
.A1(n_2407),
.A2(n_46),
.B(n_47),
.Y(n_2759)
);

AOI21xp5_ASAP7_75t_L g2760 ( 
.A1(n_2525),
.A2(n_2533),
.B(n_2488),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2328),
.B(n_46),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2330),
.B(n_46),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2336),
.B(n_47),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2338),
.Y(n_2764)
);

HB1xp67_ASAP7_75t_L g2765 ( 
.A(n_2448),
.Y(n_2765)
);

AOI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2525),
.A2(n_47),
.B(n_48),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2346),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2360),
.Y(n_2768)
);

NAND2x1p5_ASAP7_75t_L g2769 ( 
.A(n_2448),
.B(n_48),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2374),
.B(n_48),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2390),
.B(n_49),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2399),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2406),
.B(n_49),
.Y(n_2773)
);

AOI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2525),
.A2(n_50),
.B(n_51),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2398),
.B(n_50),
.Y(n_2775)
);

INVx1_ASAP7_75t_SL g2776 ( 
.A(n_2268),
.Y(n_2776)
);

AOI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_2533),
.A2(n_51),
.B(n_52),
.Y(n_2777)
);

AOI21xp5_ASAP7_75t_L g2778 ( 
.A1(n_2533),
.A2(n_51),
.B(n_52),
.Y(n_2778)
);

AOI22xp33_ASAP7_75t_L g2779 ( 
.A1(n_2359),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_SL g2780 ( 
.A(n_2541),
.B(n_54),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2398),
.B(n_53),
.Y(n_2781)
);

CKINVDCx5p33_ASAP7_75t_R g2782 ( 
.A(n_2394),
.Y(n_2782)
);

INVx4_ASAP7_75t_L g2783 ( 
.A(n_2467),
.Y(n_2783)
);

AOI21xp5_ASAP7_75t_L g2784 ( 
.A1(n_2498),
.A2(n_53),
.B(n_55),
.Y(n_2784)
);

AOI21xp5_ASAP7_75t_L g2785 ( 
.A1(n_2501),
.A2(n_55),
.B(n_56),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2383),
.B(n_55),
.Y(n_2786)
);

BUFx4f_ASAP7_75t_L g2787 ( 
.A(n_2440),
.Y(n_2787)
);

NOR2xp33_ASAP7_75t_L g2788 ( 
.A(n_2320),
.B(n_2333),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2337),
.B(n_56),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2409),
.B(n_57),
.Y(n_2790)
);

A2O1A1Ixp33_ASAP7_75t_L g2791 ( 
.A1(n_2461),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2387),
.B(n_2425),
.Y(n_2792)
);

AOI33xp33_ASAP7_75t_L g2793 ( 
.A1(n_2441),
.A2(n_60),
.A3(n_62),
.B1(n_58),
.B2(n_59),
.B3(n_61),
.Y(n_2793)
);

OAI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2412),
.A2(n_60),
.B(n_61),
.Y(n_2794)
);

INVx3_ASAP7_75t_L g2795 ( 
.A(n_2369),
.Y(n_2795)
);

AOI21x1_ASAP7_75t_L g2796 ( 
.A1(n_2447),
.A2(n_61),
.B(n_62),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_L g2797 ( 
.A(n_2343),
.B(n_63),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2429),
.B(n_64),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2364),
.B(n_2421),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2414),
.B(n_64),
.Y(n_2800)
);

NOR2xp67_ASAP7_75t_L g2801 ( 
.A(n_2558),
.B(n_64),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2422),
.B(n_2420),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_SL g2803 ( 
.A(n_2522),
.B(n_66),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2323),
.B(n_2325),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2329),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2508),
.A2(n_65),
.B(n_66),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_SL g2807 ( 
.A(n_2535),
.B(n_66),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2227),
.B(n_65),
.Y(n_2808)
);

A2O1A1Ixp33_ASAP7_75t_L g2809 ( 
.A1(n_2462),
.A2(n_68),
.B(n_65),
.C(n_67),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2344),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_SL g2811 ( 
.A(n_2544),
.B(n_69),
.Y(n_2811)
);

AOI21xp5_ASAP7_75t_L g2812 ( 
.A1(n_2510),
.A2(n_68),
.B(n_69),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2542),
.B(n_68),
.Y(n_2813)
);

AOI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2512),
.A2(n_69),
.B(n_71),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2373),
.B(n_71),
.Y(n_2815)
);

BUFx12f_ASAP7_75t_L g2816 ( 
.A(n_2453),
.Y(n_2816)
);

AOI22xp33_ASAP7_75t_L g2817 ( 
.A1(n_2439),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_2817)
);

INVx1_ASAP7_75t_SL g2818 ( 
.A(n_2524),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2401),
.B(n_2408),
.Y(n_2819)
);

AOI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2480),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2424),
.B(n_73),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2418),
.B(n_75),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2549),
.B(n_76),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_L g2824 ( 
.A1(n_2516),
.A2(n_76),
.B(n_77),
.Y(n_2824)
);

AOI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2518),
.A2(n_77),
.B(n_78),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2559),
.B(n_78),
.Y(n_2826)
);

AOI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2526),
.A2(n_78),
.B(n_79),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2530),
.B(n_2543),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2487),
.Y(n_2829)
);

OAI21x1_ASAP7_75t_L g2830 ( 
.A1(n_2485),
.A2(n_671),
.B(n_670),
.Y(n_2830)
);

OAI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2463),
.A2(n_2300),
.B1(n_2299),
.B2(n_2192),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2358),
.B(n_79),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2548),
.B(n_2550),
.Y(n_2833)
);

AOI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2479),
.A2(n_79),
.B(n_80),
.Y(n_2834)
);

O2A1O1Ixp33_ASAP7_75t_L g2835 ( 
.A1(n_2395),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2402),
.B(n_81),
.Y(n_2836)
);

AND2x4_ASAP7_75t_L g2837 ( 
.A(n_2275),
.B(n_83),
.Y(n_2837)
);

OAI22xp5_ASAP7_75t_L g2838 ( 
.A1(n_2297),
.A2(n_2303),
.B1(n_2335),
.B2(n_2318),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2341),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2487),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2489),
.Y(n_2841)
);

AOI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2382),
.A2(n_2352),
.B(n_2351),
.Y(n_2842)
);

INVx4_ASAP7_75t_L g2843 ( 
.A(n_2348),
.Y(n_2843)
);

NAND2x1p5_ASAP7_75t_L g2844 ( 
.A(n_2362),
.B(n_83),
.Y(n_2844)
);

OAI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2366),
.A2(n_84),
.B(n_85),
.Y(n_2845)
);

OAI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2388),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_2846)
);

AOI21xp5_ASAP7_75t_L g2847 ( 
.A1(n_2392),
.A2(n_85),
.B(n_86),
.Y(n_2847)
);

AOI21xp5_ASAP7_75t_L g2848 ( 
.A1(n_2307),
.A2(n_87),
.B(n_88),
.Y(n_2848)
);

NOR2xp33_ASAP7_75t_SL g2849 ( 
.A(n_2334),
.B(n_2427),
.Y(n_2849)
);

OR2x6_ASAP7_75t_L g2850 ( 
.A(n_2504),
.B(n_88),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2432),
.B(n_89),
.Y(n_2851)
);

INVx3_ASAP7_75t_L g2852 ( 
.A(n_2369),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2417),
.Y(n_2853)
);

AOI21xp5_ASAP7_75t_L g2854 ( 
.A1(n_2379),
.A2(n_2198),
.B(n_2197),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2256),
.A2(n_89),
.B(n_90),
.Y(n_2855)
);

INVxp67_ASAP7_75t_L g2856 ( 
.A(n_2193),
.Y(n_2856)
);

OAI21xp5_ASAP7_75t_L g2857 ( 
.A1(n_2367),
.A2(n_89),
.B(n_90),
.Y(n_2857)
);

AOI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2493),
.A2(n_91),
.B(n_92),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2371),
.B(n_91),
.Y(n_2859)
);

OAI21xp33_ASAP7_75t_L g2860 ( 
.A1(n_2380),
.A2(n_91),
.B(n_92),
.Y(n_2860)
);

OAI21xp33_ASAP7_75t_L g2861 ( 
.A1(n_2444),
.A2(n_92),
.B(n_93),
.Y(n_2861)
);

NAND2x1_ASAP7_75t_L g2862 ( 
.A(n_2417),
.B(n_93),
.Y(n_2862)
);

O2A1O1Ixp33_ASAP7_75t_L g2863 ( 
.A1(n_2457),
.A2(n_2491),
.B(n_2400),
.C(n_2188),
.Y(n_2863)
);

AOI21xp5_ASAP7_75t_L g2864 ( 
.A1(n_2450),
.A2(n_94),
.B(n_95),
.Y(n_2864)
);

BUFx2_ASAP7_75t_L g2865 ( 
.A(n_2404),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_SL g2866 ( 
.A(n_2484),
.B(n_95),
.Y(n_2866)
);

CKINVDCx20_ASAP7_75t_R g2867 ( 
.A(n_2513),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_SL g2868 ( 
.A(n_2389),
.B(n_2435),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_L g2869 ( 
.A(n_2212),
.B(n_94),
.Y(n_2869)
);

AOI21xp5_ASAP7_75t_L g2870 ( 
.A1(n_2451),
.A2(n_94),
.B(n_96),
.Y(n_2870)
);

OAI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2413),
.A2(n_96),
.B(n_97),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2375),
.B(n_97),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2376),
.B(n_98),
.Y(n_2873)
);

AOI21xp5_ASAP7_75t_L g2874 ( 
.A1(n_2495),
.A2(n_2496),
.B(n_2490),
.Y(n_2874)
);

AOI22xp33_ASAP7_75t_L g2875 ( 
.A1(n_2449),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_2875)
);

A2O1A1Ixp33_ASAP7_75t_L g2876 ( 
.A1(n_2481),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2489),
.Y(n_2877)
);

AOI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2415),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_SL g2879 ( 
.A(n_2437),
.B(n_102),
.Y(n_2879)
);

AOI21xp5_ASAP7_75t_L g2880 ( 
.A1(n_2294),
.A2(n_101),
.B(n_102),
.Y(n_2880)
);

AOI21xp5_ASAP7_75t_L g2881 ( 
.A1(n_2482),
.A2(n_102),
.B(n_103),
.Y(n_2881)
);

AOI21xp5_ASAP7_75t_L g2882 ( 
.A1(n_2403),
.A2(n_103),
.B(n_104),
.Y(n_2882)
);

BUFx3_ASAP7_75t_L g2883 ( 
.A(n_2436),
.Y(n_2883)
);

AOI21xp5_ASAP7_75t_L g2884 ( 
.A1(n_2411),
.A2(n_103),
.B(n_104),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2331),
.B(n_2365),
.Y(n_2885)
);

AOI21xp5_ASAP7_75t_L g2886 ( 
.A1(n_2454),
.A2(n_104),
.B(n_105),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_SL g2887 ( 
.A(n_2434),
.B(n_106),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2445),
.B(n_105),
.Y(n_2888)
);

BUFx6f_ASAP7_75t_L g2889 ( 
.A(n_2363),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2502),
.B(n_2509),
.Y(n_2890)
);

OR2x2_ASAP7_75t_L g2891 ( 
.A(n_2515),
.B(n_106),
.Y(n_2891)
);

INVxp67_ASAP7_75t_L g2892 ( 
.A(n_2520),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2529),
.B(n_106),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2452),
.A2(n_2486),
.B(n_2203),
.Y(n_2894)
);

BUFx2_ASAP7_75t_L g2895 ( 
.A(n_2355),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_L g2896 ( 
.A1(n_2426),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_2896)
);

CKINVDCx5p33_ASAP7_75t_R g2897 ( 
.A(n_2410),
.Y(n_2897)
);

AOI21xp5_ASAP7_75t_L g2898 ( 
.A1(n_2201),
.A2(n_107),
.B(n_108),
.Y(n_2898)
);

OAI321xp33_ASAP7_75t_L g2899 ( 
.A1(n_2553),
.A2(n_110),
.A3(n_112),
.B1(n_107),
.B2(n_109),
.C(n_111),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2438),
.B(n_110),
.Y(n_2900)
);

INVx1_ASAP7_75t_SL g2901 ( 
.A(n_2319),
.Y(n_2901)
);

OAI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2340),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2494),
.Y(n_2903)
);

OAI321xp33_ASAP7_75t_L g2904 ( 
.A1(n_2350),
.A2(n_114),
.A3(n_116),
.B1(n_112),
.B2(n_113),
.C(n_115),
.Y(n_2904)
);

AOI21x1_ASAP7_75t_L g2905 ( 
.A1(n_2497),
.A2(n_113),
.B(n_115),
.Y(n_2905)
);

OR2x2_ASAP7_75t_L g2906 ( 
.A(n_2354),
.B(n_115),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2310),
.B(n_116),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2209),
.Y(n_2908)
);

BUFx10_ASAP7_75t_L g2909 ( 
.A(n_2315),
.Y(n_2909)
);

NOR2x1_ASAP7_75t_L g2910 ( 
.A(n_2229),
.B(n_116),
.Y(n_2910)
);

AOI21xp5_ASAP7_75t_L g2911 ( 
.A1(n_2234),
.A2(n_117),
.B(n_118),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2260),
.B(n_117),
.Y(n_2912)
);

OAI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2478),
.A2(n_117),
.B(n_118),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2492),
.A2(n_118),
.B(n_119),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2492),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2492),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_2492),
.B(n_120),
.Y(n_2917)
);

A2O1A1Ixp33_ASAP7_75t_L g2918 ( 
.A1(n_2492),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2208),
.B(n_120),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2468),
.A2(n_121),
.B(n_122),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2468),
.A2(n_121),
.B(n_122),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2468),
.Y(n_2922)
);

AOI21xp5_ASAP7_75t_L g2923 ( 
.A1(n_2468),
.A2(n_122),
.B(n_123),
.Y(n_2923)
);

A2O1A1Ixp33_ASAP7_75t_L g2924 ( 
.A1(n_2208),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_2924)
);

OAI21x1_ASAP7_75t_L g2925 ( 
.A1(n_2442),
.A2(n_674),
.B(n_673),
.Y(n_2925)
);

BUFx5_ASAP7_75t_L g2926 ( 
.A(n_2332),
.Y(n_2926)
);

NAND2x2_ASAP7_75t_L g2927 ( 
.A(n_2215),
.B(n_124),
.Y(n_2927)
);

NOR2xp67_ASAP7_75t_SL g2928 ( 
.A(n_2446),
.B(n_123),
.Y(n_2928)
);

AOI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2468),
.A2(n_125),
.B(n_126),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2468),
.Y(n_2930)
);

INVx2_ASAP7_75t_SL g2931 ( 
.A(n_2483),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2468),
.A2(n_125),
.B(n_126),
.Y(n_2932)
);

A2O1A1Ixp33_ASAP7_75t_L g2933 ( 
.A1(n_2208),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_2933)
);

BUFx4f_ASAP7_75t_L g2934 ( 
.A(n_2251),
.Y(n_2934)
);

AOI21xp5_ASAP7_75t_L g2935 ( 
.A1(n_2468),
.A2(n_127),
.B(n_128),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2208),
.B(n_127),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2208),
.B(n_129),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2208),
.B(n_129),
.Y(n_2938)
);

BUFx6f_ASAP7_75t_L g2939 ( 
.A(n_2313),
.Y(n_2939)
);

NOR2x1_ASAP7_75t_R g2940 ( 
.A(n_2189),
.B(n_130),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2208),
.B(n_130),
.Y(n_2941)
);

INVx5_ASAP7_75t_L g2942 ( 
.A(n_2313),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2468),
.Y(n_2943)
);

AO21x1_ASAP7_75t_L g2944 ( 
.A1(n_2357),
.A2(n_674),
.B(n_673),
.Y(n_2944)
);

AOI21xp5_ASAP7_75t_L g2945 ( 
.A1(n_2468),
.A2(n_131),
.B(n_132),
.Y(n_2945)
);

AOI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2468),
.A2(n_131),
.B(n_132),
.Y(n_2946)
);

AO21x1_ASAP7_75t_L g2947 ( 
.A1(n_2357),
.A2(n_676),
.B(n_675),
.Y(n_2947)
);

O2A1O1Ixp33_ASAP7_75t_L g2948 ( 
.A1(n_2245),
.A2(n_135),
.B(n_133),
.C(n_134),
.Y(n_2948)
);

INVx1_ASAP7_75t_SL g2949 ( 
.A(n_2507),
.Y(n_2949)
);

AOI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2468),
.A2(n_133),
.B(n_134),
.Y(n_2950)
);

AOI21xp5_ASAP7_75t_L g2951 ( 
.A1(n_2468),
.A2(n_133),
.B(n_134),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2249),
.Y(n_2952)
);

AOI22xp5_ASAP7_75t_L g2953 ( 
.A1(n_2288),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2208),
.B(n_135),
.Y(n_2954)
);

AOI21xp5_ASAP7_75t_L g2955 ( 
.A1(n_2468),
.A2(n_136),
.B(n_137),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2208),
.B(n_138),
.Y(n_2956)
);

NOR3xp33_ASAP7_75t_L g2957 ( 
.A(n_2277),
.B(n_140),
.C(n_139),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2208),
.B(n_138),
.Y(n_2958)
);

OAI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2208),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_SL g2960 ( 
.A(n_2507),
.B(n_141),
.Y(n_2960)
);

AOI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2468),
.A2(n_139),
.B(n_141),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2208),
.B(n_141),
.Y(n_2962)
);

INVxp67_ASAP7_75t_SL g2963 ( 
.A(n_2507),
.Y(n_2963)
);

INVxp67_ASAP7_75t_L g2964 ( 
.A(n_2507),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2208),
.B(n_142),
.Y(n_2965)
);

AOI21xp5_ASAP7_75t_L g2966 ( 
.A1(n_2468),
.A2(n_142),
.B(n_143),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2208),
.B(n_142),
.Y(n_2967)
);

INVx3_ASAP7_75t_L g2968 ( 
.A(n_2378),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2208),
.B(n_143),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2468),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2249),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2468),
.Y(n_2972)
);

NAND2xp33_ASAP7_75t_L g2973 ( 
.A(n_2313),
.B(n_144),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2208),
.B(n_143),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2208),
.B(n_144),
.Y(n_2975)
);

NOR3xp33_ASAP7_75t_L g2976 ( 
.A(n_2277),
.B(n_146),
.C(n_145),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_L g2977 ( 
.A(n_2288),
.B(n_144),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2249),
.Y(n_2978)
);

INVx3_ASAP7_75t_L g2979 ( 
.A(n_2378),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_SL g2980 ( 
.A(n_2507),
.B(n_146),
.Y(n_2980)
);

A2O1A1Ixp33_ASAP7_75t_L g2981 ( 
.A1(n_2208),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2208),
.B(n_145),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2208),
.B(n_147),
.Y(n_2983)
);

AOI21xp33_ASAP7_75t_L g2984 ( 
.A1(n_2305),
.A2(n_147),
.B(n_148),
.Y(n_2984)
);

INVxp67_ASAP7_75t_L g2985 ( 
.A(n_2507),
.Y(n_2985)
);

NOR2xp33_ASAP7_75t_L g2986 ( 
.A(n_2288),
.B(n_148),
.Y(n_2986)
);

OAI21x1_ASAP7_75t_L g2987 ( 
.A1(n_2442),
.A2(n_676),
.B(n_675),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2249),
.Y(n_2988)
);

A2O1A1Ixp33_ASAP7_75t_L g2989 ( 
.A1(n_2208),
.A2(n_150),
.B(n_148),
.C(n_149),
.Y(n_2989)
);

NOR3xp33_ASAP7_75t_L g2990 ( 
.A(n_2277),
.B(n_151),
.C(n_150),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2468),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2208),
.B(n_149),
.Y(n_2992)
);

BUFx6f_ASAP7_75t_L g2993 ( 
.A(n_2313),
.Y(n_2993)
);

OAI22xp5_ASAP7_75t_L g2994 ( 
.A1(n_2208),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2468),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2208),
.B(n_152),
.Y(n_2996)
);

AND2x4_ASAP7_75t_L g2997 ( 
.A(n_2208),
.B(n_152),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2208),
.B(n_152),
.Y(n_2998)
);

HB1xp67_ASAP7_75t_L g2999 ( 
.A(n_2507),
.Y(n_2999)
);

AO21x1_ASAP7_75t_L g3000 ( 
.A1(n_2357),
.A2(n_678),
.B(n_677),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2208),
.B(n_153),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2468),
.Y(n_3002)
);

AND2x2_ASAP7_75t_SL g3003 ( 
.A(n_2326),
.B(n_153),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_SL g3004 ( 
.A(n_2507),
.B(n_154),
.Y(n_3004)
);

NAND3xp33_ASAP7_75t_SL g3005 ( 
.A(n_2302),
.B(n_153),
.C(n_154),
.Y(n_3005)
);

OAI21xp33_ASAP7_75t_L g3006 ( 
.A1(n_2246),
.A2(n_154),
.B(n_155),
.Y(n_3006)
);

OR2x2_ASAP7_75t_L g3007 ( 
.A(n_2272),
.B(n_155),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2208),
.B(n_155),
.Y(n_3008)
);

AOI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_2468),
.A2(n_156),
.B(n_157),
.Y(n_3009)
);

INVx2_ASAP7_75t_SL g3010 ( 
.A(n_2483),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_SL g3011 ( 
.A(n_2507),
.B(n_157),
.Y(n_3011)
);

AOI21xp5_ASAP7_75t_L g3012 ( 
.A1(n_2468),
.A2(n_156),
.B(n_157),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2288),
.A2(n_159),
.B1(n_156),
.B2(n_158),
.Y(n_3013)
);

AOI21xp5_ASAP7_75t_L g3014 ( 
.A1(n_2468),
.A2(n_158),
.B(n_159),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_SL g3015 ( 
.A(n_2507),
.B(n_160),
.Y(n_3015)
);

BUFx3_ASAP7_75t_L g3016 ( 
.A(n_2274),
.Y(n_3016)
);

BUFx2_ASAP7_75t_L g3017 ( 
.A(n_2507),
.Y(n_3017)
);

AOI21xp5_ASAP7_75t_L g3018 ( 
.A1(n_2468),
.A2(n_158),
.B(n_160),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2288),
.B(n_160),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2208),
.B(n_161),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2468),
.A2(n_161),
.B(n_162),
.Y(n_3021)
);

INVx11_ASAP7_75t_L g3022 ( 
.A(n_2204),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2208),
.B(n_161),
.Y(n_3023)
);

OAI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2368),
.A2(n_162),
.B(n_163),
.Y(n_3024)
);

AOI21xp5_ASAP7_75t_L g3025 ( 
.A1(n_2468),
.A2(n_162),
.B(n_163),
.Y(n_3025)
);

NAND2xp33_ASAP7_75t_L g3026 ( 
.A(n_2313),
.B(n_164),
.Y(n_3026)
);

OAI21xp5_ASAP7_75t_L g3027 ( 
.A1(n_2368),
.A2(n_163),
.B(n_164),
.Y(n_3027)
);

O2A1O1Ixp33_ASAP7_75t_L g3028 ( 
.A1(n_2245),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_3028)
);

AO21x1_ASAP7_75t_L g3029 ( 
.A1(n_2357),
.A2(n_678),
.B(n_677),
.Y(n_3029)
);

AOI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2468),
.A2(n_165),
.B(n_166),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2468),
.Y(n_3031)
);

OAI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_2368),
.A2(n_167),
.B(n_168),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2208),
.B(n_167),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2208),
.B(n_167),
.Y(n_3034)
);

AOI21xp5_ASAP7_75t_L g3035 ( 
.A1(n_2468),
.A2(n_168),
.B(n_169),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2208),
.B(n_168),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_SL g3037 ( 
.A(n_2507),
.B(n_170),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_L g3038 ( 
.A(n_2288),
.B(n_169),
.Y(n_3038)
);

AOI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2322),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_3039)
);

O2A1O1Ixp33_ASAP7_75t_L g3040 ( 
.A1(n_2245),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2208),
.B(n_171),
.Y(n_3041)
);

BUFx8_ASAP7_75t_L g3042 ( 
.A(n_2204),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2208),
.B(n_172),
.Y(n_3043)
);

AOI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2468),
.A2(n_172),
.B(n_173),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2208),
.B(n_173),
.Y(n_3045)
);

AOI21xp33_ASAP7_75t_L g3046 ( 
.A1(n_2305),
.A2(n_174),
.B(n_175),
.Y(n_3046)
);

O2A1O1Ixp33_ASAP7_75t_SL g3047 ( 
.A1(n_2292),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2468),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2208),
.B(n_174),
.Y(n_3049)
);

AOI21xp33_ASAP7_75t_L g3050 ( 
.A1(n_2305),
.A2(n_175),
.B(n_176),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_SL g3051 ( 
.A(n_2507),
.B(n_177),
.Y(n_3051)
);

AO21x1_ASAP7_75t_L g3052 ( 
.A1(n_2357),
.A2(n_681),
.B(n_680),
.Y(n_3052)
);

AOI21xp5_ASAP7_75t_L g3053 ( 
.A1(n_2468),
.A2(n_176),
.B(n_177),
.Y(n_3053)
);

INVx3_ASAP7_75t_L g3054 ( 
.A(n_2378),
.Y(n_3054)
);

AOI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2468),
.A2(n_177),
.B(n_178),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2208),
.B(n_179),
.Y(n_3056)
);

CKINVDCx5p33_ASAP7_75t_R g3057 ( 
.A(n_2189),
.Y(n_3057)
);

OAI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_2368),
.A2(n_179),
.B(n_180),
.Y(n_3058)
);

NAND2x1p5_ASAP7_75t_L g3059 ( 
.A(n_2274),
.B(n_180),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2208),
.B(n_181),
.Y(n_3060)
);

NOR3xp33_ASAP7_75t_L g3061 ( 
.A(n_2277),
.B(n_183),
.C(n_182),
.Y(n_3061)
);

BUFx4f_ASAP7_75t_L g3062 ( 
.A(n_2251),
.Y(n_3062)
);

AOI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2468),
.A2(n_181),
.B(n_182),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2208),
.B(n_183),
.Y(n_3064)
);

O2A1O1Ixp33_ASAP7_75t_L g3065 ( 
.A1(n_2245),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_3065)
);

OAI22xp5_ASAP7_75t_L g3066 ( 
.A1(n_2208),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2208),
.B(n_184),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2208),
.B(n_185),
.Y(n_3068)
);

OAI21xp33_ASAP7_75t_L g3069 ( 
.A1(n_2246),
.A2(n_186),
.B(n_187),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2468),
.Y(n_3070)
);

AOI21x1_ASAP7_75t_L g3071 ( 
.A1(n_2468),
.A2(n_187),
.B(n_188),
.Y(n_3071)
);

A2O1A1Ixp33_ASAP7_75t_L g3072 ( 
.A1(n_2208),
.A2(n_189),
.B(n_187),
.C(n_188),
.Y(n_3072)
);

O2A1O1Ixp33_ASAP7_75t_L g3073 ( 
.A1(n_2245),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_3073)
);

AOI21xp5_ASAP7_75t_L g3074 ( 
.A1(n_2468),
.A2(n_189),
.B(n_190),
.Y(n_3074)
);

A2O1A1Ixp33_ASAP7_75t_L g3075 ( 
.A1(n_2208),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2468),
.A2(n_191),
.B(n_192),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_SL g3077 ( 
.A(n_2507),
.B(n_193),
.Y(n_3077)
);

AOI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2468),
.A2(n_192),
.B(n_193),
.Y(n_3078)
);

BUFx4f_ASAP7_75t_L g3079 ( 
.A(n_2251),
.Y(n_3079)
);

INVx3_ASAP7_75t_L g3080 ( 
.A(n_2378),
.Y(n_3080)
);

O2A1O1Ixp5_ASAP7_75t_L g3081 ( 
.A1(n_2292),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2208),
.B(n_194),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2468),
.A2(n_194),
.B(n_195),
.Y(n_3083)
);

BUFx6f_ASAP7_75t_L g3084 ( 
.A(n_2313),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2468),
.A2(n_196),
.B(n_197),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2208),
.B(n_196),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_L g3087 ( 
.A(n_2288),
.B(n_196),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2468),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2208),
.B(n_198),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_SL g3090 ( 
.A(n_2507),
.B(n_199),
.Y(n_3090)
);

BUFx6f_ASAP7_75t_L g3091 ( 
.A(n_2313),
.Y(n_3091)
);

AOI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2468),
.A2(n_198),
.B(n_199),
.Y(n_3092)
);

AND2x4_ASAP7_75t_L g3093 ( 
.A(n_2208),
.B(n_199),
.Y(n_3093)
);

OAI321xp33_ASAP7_75t_L g3094 ( 
.A1(n_2277),
.A2(n_202),
.A3(n_204),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_3094)
);

AOI21xp5_ASAP7_75t_L g3095 ( 
.A1(n_2468),
.A2(n_200),
.B(n_201),
.Y(n_3095)
);

AOI21x1_ASAP7_75t_L g3096 ( 
.A1(n_2468),
.A2(n_200),
.B(n_201),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2249),
.Y(n_3097)
);

BUFx6f_ASAP7_75t_L g3098 ( 
.A(n_2313),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_2468),
.A2(n_202),
.B(n_203),
.Y(n_3099)
);

AOI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2468),
.A2(n_202),
.B(n_204),
.Y(n_3100)
);

BUFx12f_ASAP7_75t_L g3101 ( 
.A(n_2189),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2208),
.B(n_204),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2208),
.B(n_205),
.Y(n_3103)
);

INVx4_ASAP7_75t_L g3104 ( 
.A(n_2251),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2208),
.B(n_205),
.Y(n_3105)
);

AOI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_2468),
.A2(n_205),
.B(n_206),
.Y(n_3106)
);

BUFx4f_ASAP7_75t_L g3107 ( 
.A(n_2251),
.Y(n_3107)
);

INVx2_ASAP7_75t_SL g3108 ( 
.A(n_2483),
.Y(n_3108)
);

OAI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2368),
.A2(n_206),
.B(n_207),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_SL g3110 ( 
.A(n_2507),
.B(n_208),
.Y(n_3110)
);

AOI21xp5_ASAP7_75t_L g3111 ( 
.A1(n_2468),
.A2(n_207),
.B(n_208),
.Y(n_3111)
);

AND2x2_ASAP7_75t_L g3112 ( 
.A(n_2208),
.B(n_208),
.Y(n_3112)
);

AOI21xp5_ASAP7_75t_L g3113 ( 
.A1(n_2468),
.A2(n_209),
.B(n_210),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2249),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2468),
.A2(n_209),
.B(n_210),
.Y(n_3115)
);

AOI21xp5_ASAP7_75t_L g3116 ( 
.A1(n_2468),
.A2(n_210),
.B(n_211),
.Y(n_3116)
);

INVx3_ASAP7_75t_L g3117 ( 
.A(n_2378),
.Y(n_3117)
);

AOI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2468),
.A2(n_211),
.B(n_212),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2208),
.B(n_211),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2468),
.Y(n_3120)
);

OAI22xp5_ASAP7_75t_L g3121 ( 
.A1(n_2208),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2208),
.B(n_212),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2208),
.B(n_213),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_2208),
.B(n_213),
.Y(n_3124)
);

OAI21xp33_ASAP7_75t_L g3125 ( 
.A1(n_2246),
.A2(n_214),
.B(n_215),
.Y(n_3125)
);

AOI21x1_ASAP7_75t_L g3126 ( 
.A1(n_2468),
.A2(n_214),
.B(n_215),
.Y(n_3126)
);

O2A1O1Ixp33_ASAP7_75t_L g3127 ( 
.A1(n_2245),
.A2(n_217),
.B(n_215),
.C(n_216),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2208),
.B(n_216),
.Y(n_3128)
);

HB1xp67_ASAP7_75t_L g3129 ( 
.A(n_2507),
.Y(n_3129)
);

OAI22xp33_ASAP7_75t_L g3130 ( 
.A1(n_2277),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_3130)
);

BUFx3_ASAP7_75t_L g3131 ( 
.A(n_2274),
.Y(n_3131)
);

BUFx6f_ASAP7_75t_L g3132 ( 
.A(n_2313),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2208),
.B(n_217),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2249),
.Y(n_3134)
);

AOI21xp5_ASAP7_75t_L g3135 ( 
.A1(n_2468),
.A2(n_218),
.B(n_219),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2322),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2208),
.B(n_219),
.Y(n_3137)
);

BUFx6f_ASAP7_75t_L g3138 ( 
.A(n_2313),
.Y(n_3138)
);

OAI22xp5_ASAP7_75t_L g3139 ( 
.A1(n_2208),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_2208),
.B(n_220),
.Y(n_3140)
);

OAI22xp5_ASAP7_75t_L g3141 ( 
.A1(n_2208),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_3141)
);

BUFx6f_ASAP7_75t_L g3142 ( 
.A(n_2313),
.Y(n_3142)
);

AOI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_2468),
.A2(n_224),
.B(n_225),
.Y(n_3143)
);

INVx8_ASAP7_75t_L g3144 ( 
.A(n_2251),
.Y(n_3144)
);

O2A1O1Ixp33_ASAP7_75t_L g3145 ( 
.A1(n_2245),
.A2(n_226),
.B(n_224),
.C(n_225),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2208),
.B(n_225),
.Y(n_3146)
);

AOI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_2322),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_3147)
);

AOI21xp5_ASAP7_75t_L g3148 ( 
.A1(n_2468),
.A2(n_226),
.B(n_227),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2249),
.Y(n_3149)
);

NOR2xp33_ASAP7_75t_L g3150 ( 
.A(n_2288),
.B(n_227),
.Y(n_3150)
);

A2O1A1Ixp33_ASAP7_75t_L g3151 ( 
.A1(n_2208),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2249),
.Y(n_3152)
);

NOR2xp33_ASAP7_75t_R g3153 ( 
.A(n_2189),
.B(n_229),
.Y(n_3153)
);

AOI21xp5_ASAP7_75t_L g3154 ( 
.A1(n_2468),
.A2(n_230),
.B(n_231),
.Y(n_3154)
);

BUFx6f_ASAP7_75t_L g3155 ( 
.A(n_2313),
.Y(n_3155)
);

A2O1A1Ixp33_ASAP7_75t_L g3156 ( 
.A1(n_2208),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_3156)
);

BUFx4f_ASAP7_75t_L g3157 ( 
.A(n_2251),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2468),
.A2(n_232),
.B(n_233),
.Y(n_3158)
);

AO21x1_ASAP7_75t_L g3159 ( 
.A1(n_2357),
.A2(n_681),
.B(n_680),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2249),
.Y(n_3160)
);

HB1xp67_ASAP7_75t_L g3161 ( 
.A(n_2507),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2208),
.B(n_232),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_SL g3163 ( 
.A(n_2507),
.B(n_234),
.Y(n_3163)
);

INVx3_ASAP7_75t_L g3164 ( 
.A(n_2378),
.Y(n_3164)
);

AOI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_2468),
.A2(n_233),
.B(n_234),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_L g3166 ( 
.A(n_2288),
.B(n_233),
.Y(n_3166)
);

NOR2xp33_ASAP7_75t_L g3167 ( 
.A(n_2288),
.B(n_235),
.Y(n_3167)
);

BUFx8_ASAP7_75t_L g3168 ( 
.A(n_2204),
.Y(n_3168)
);

AOI21xp5_ASAP7_75t_L g3169 ( 
.A1(n_2468),
.A2(n_235),
.B(n_236),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2249),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_2208),
.B(n_235),
.Y(n_3171)
);

OAI22xp5_ASAP7_75t_L g3172 ( 
.A1(n_2208),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_3172)
);

AND2x2_ASAP7_75t_L g3173 ( 
.A(n_2208),
.B(n_236),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2208),
.B(n_237),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2208),
.B(n_238),
.Y(n_3175)
);

AOI21xp5_ASAP7_75t_L g3176 ( 
.A1(n_2468),
.A2(n_239),
.B(n_240),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2249),
.Y(n_3177)
);

BUFx6f_ASAP7_75t_L g3178 ( 
.A(n_2313),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2208),
.B(n_239),
.Y(n_3179)
);

OAI22xp5_ASAP7_75t_L g3180 ( 
.A1(n_2208),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2208),
.B(n_240),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2208),
.B(n_241),
.Y(n_3182)
);

A2O1A1Ixp33_ASAP7_75t_L g3183 ( 
.A1(n_2208),
.A2(n_244),
.B(n_242),
.C(n_243),
.Y(n_3183)
);

AOI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_2468),
.A2(n_242),
.B(n_243),
.Y(n_3184)
);

NOR2xp33_ASAP7_75t_L g3185 ( 
.A(n_2288),
.B(n_242),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2468),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2208),
.B(n_243),
.Y(n_3187)
);

AOI21xp33_ASAP7_75t_L g3188 ( 
.A1(n_2305),
.A2(n_244),
.B(n_245),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2468),
.A2(n_244),
.B(n_245),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2208),
.B(n_246),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_2468),
.A2(n_246),
.B(n_247),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_2208),
.B(n_247),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_2468),
.A2(n_247),
.B(n_248),
.Y(n_3193)
);

AO22x1_ASAP7_75t_L g3194 ( 
.A1(n_2309),
.A2(n_250),
.B1(n_251),
.B2(n_249),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2468),
.Y(n_3195)
);

BUFx2_ASAP7_75t_L g3196 ( 
.A(n_2507),
.Y(n_3196)
);

OAI321xp33_ASAP7_75t_L g3197 ( 
.A1(n_2277),
.A2(n_250),
.A3(n_252),
.B1(n_248),
.B2(n_249),
.C(n_251),
.Y(n_3197)
);

AOI21xp5_ASAP7_75t_L g3198 ( 
.A1(n_2468),
.A2(n_249),
.B(n_250),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2996),
.Y(n_3199)
);

AOI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_2624),
.A2(n_251),
.B(n_252),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2571),
.B(n_252),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3020),
.Y(n_3202)
);

AOI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_2639),
.A2(n_253),
.B(n_254),
.Y(n_3203)
);

O2A1O1Ixp33_ASAP7_75t_L g3204 ( 
.A1(n_2627),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_3204)
);

CKINVDCx20_ASAP7_75t_R g3205 ( 
.A(n_3042),
.Y(n_3205)
);

BUFx12f_ASAP7_75t_L g3206 ( 
.A(n_3042),
.Y(n_3206)
);

AND2x2_ASAP7_75t_L g3207 ( 
.A(n_2952),
.B(n_2971),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3105),
.Y(n_3208)
);

A2O1A1Ixp33_ASAP7_75t_L g3209 ( 
.A1(n_2656),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_3209)
);

NAND3x1_ASAP7_75t_L g3210 ( 
.A(n_2957),
.B(n_255),
.C(n_256),
.Y(n_3210)
);

HB1xp67_ASAP7_75t_L g3211 ( 
.A(n_2949),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3112),
.Y(n_3212)
);

NOR2xp67_ASAP7_75t_L g3213 ( 
.A(n_2564),
.B(n_256),
.Y(n_3213)
);

INVx4_ASAP7_75t_L g3214 ( 
.A(n_3144),
.Y(n_3214)
);

AND2x4_ASAP7_75t_L g3215 ( 
.A(n_2978),
.B(n_256),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3124),
.Y(n_3216)
);

OR2x6_ASAP7_75t_L g3217 ( 
.A(n_3144),
.B(n_257),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2576),
.Y(n_3218)
);

INVxp67_ASAP7_75t_L g3219 ( 
.A(n_2999),
.Y(n_3219)
);

NOR3xp33_ASAP7_75t_SL g3220 ( 
.A(n_2897),
.B(n_257),
.C(n_258),
.Y(n_3220)
);

OR2x2_ASAP7_75t_L g3221 ( 
.A(n_2631),
.B(n_257),
.Y(n_3221)
);

OAI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_2720),
.A2(n_258),
.B(n_259),
.Y(n_3222)
);

OR2x6_ASAP7_75t_L g3223 ( 
.A(n_3144),
.B(n_258),
.Y(n_3223)
);

NOR2xp33_ASAP7_75t_L g3224 ( 
.A(n_2727),
.B(n_259),
.Y(n_3224)
);

O2A1O1Ixp33_ASAP7_75t_L g3225 ( 
.A1(n_2831),
.A2(n_262),
.B(n_259),
.C(n_261),
.Y(n_3225)
);

O2A1O1Ixp33_ASAP7_75t_L g3226 ( 
.A1(n_2984),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_3226)
);

CKINVDCx14_ASAP7_75t_R g3227 ( 
.A(n_3153),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2589),
.Y(n_3228)
);

AOI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_2874),
.A2(n_261),
.B(n_263),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_SL g3230 ( 
.A(n_2657),
.B(n_682),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2764),
.Y(n_3231)
);

AOI21xp5_ASAP7_75t_L g3232 ( 
.A1(n_2760),
.A2(n_263),
.B(n_264),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3133),
.Y(n_3233)
);

AND2x4_ASAP7_75t_L g3234 ( 
.A(n_2988),
.B(n_264),
.Y(n_3234)
);

NOR2xp33_ASAP7_75t_L g3235 ( 
.A(n_2560),
.B(n_265),
.Y(n_3235)
);

AOI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_2804),
.A2(n_265),
.B(n_266),
.Y(n_3236)
);

INVx1_ASAP7_75t_SL g3237 ( 
.A(n_3017),
.Y(n_3237)
);

O2A1O1Ixp5_ASAP7_75t_L g3238 ( 
.A1(n_2879),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2600),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_3097),
.B(n_267),
.Y(n_3240)
);

XOR2x2_ASAP7_75t_L g3241 ( 
.A(n_3003),
.B(n_267),
.Y(n_3241)
);

CKINVDCx20_ASAP7_75t_R g3242 ( 
.A(n_3168),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_2868),
.B(n_268),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3140),
.Y(n_3244)
);

AND2x4_ASAP7_75t_L g3245 ( 
.A(n_3114),
.B(n_268),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3171),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3173),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3134),
.B(n_269),
.Y(n_3248)
);

HB1xp67_ASAP7_75t_L g3249 ( 
.A(n_3196),
.Y(n_3249)
);

AOI21xp5_ASAP7_75t_L g3250 ( 
.A1(n_2828),
.A2(n_271),
.B(n_272),
.Y(n_3250)
);

INVx3_ASAP7_75t_L g3251 ( 
.A(n_2662),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3149),
.B(n_271),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3192),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_2610),
.A2(n_271),
.B(n_272),
.Y(n_3254)
);

O2A1O1Ixp33_ASAP7_75t_SL g3255 ( 
.A1(n_2862),
.A2(n_275),
.B(n_273),
.C(n_274),
.Y(n_3255)
);

AND2x2_ASAP7_75t_SL g3256 ( 
.A(n_2726),
.B(n_273),
.Y(n_3256)
);

AOI22xp5_ASAP7_75t_L g3257 ( 
.A1(n_2976),
.A2(n_276),
.B1(n_273),
.B2(n_275),
.Y(n_3257)
);

CKINVDCx5p33_ASAP7_75t_R g3258 ( 
.A(n_2669),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2574),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_3152),
.B(n_275),
.Y(n_3260)
);

AOI21xp5_ASAP7_75t_L g3261 ( 
.A1(n_2854),
.A2(n_276),
.B(n_277),
.Y(n_3261)
);

CKINVDCx6p67_ASAP7_75t_R g3262 ( 
.A(n_2669),
.Y(n_3262)
);

NOR2xp33_ASAP7_75t_L g3263 ( 
.A(n_2583),
.B(n_276),
.Y(n_3263)
);

AND2x2_ASAP7_75t_L g3264 ( 
.A(n_3160),
.B(n_277),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2585),
.Y(n_3265)
);

OAI22xp5_ASAP7_75t_L g3266 ( 
.A1(n_3170),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_SL g3267 ( 
.A(n_2818),
.B(n_686),
.Y(n_3267)
);

AOI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_2644),
.A2(n_2646),
.B(n_2645),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2598),
.Y(n_3269)
);

NOR2xp33_ASAP7_75t_SL g3270 ( 
.A(n_2662),
.B(n_278),
.Y(n_3270)
);

O2A1O1Ixp33_ASAP7_75t_L g3271 ( 
.A1(n_3188),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2716),
.Y(n_3272)
);

INVx3_ASAP7_75t_L g3273 ( 
.A(n_2934),
.Y(n_3273)
);

AOI21xp5_ASAP7_75t_L g3274 ( 
.A1(n_2649),
.A2(n_280),
.B(n_281),
.Y(n_3274)
);

AOI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_2651),
.A2(n_281),
.B(n_282),
.Y(n_3275)
);

AOI21xp5_ASAP7_75t_L g3276 ( 
.A1(n_2654),
.A2(n_282),
.B(n_283),
.Y(n_3276)
);

BUFx12f_ASAP7_75t_L g3277 ( 
.A(n_3168),
.Y(n_3277)
);

AOI22x1_ASAP7_75t_L g3278 ( 
.A1(n_2683),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_3278)
);

AOI22xp5_ASAP7_75t_L g3279 ( 
.A1(n_2990),
.A2(n_287),
.B1(n_284),
.B2(n_286),
.Y(n_3279)
);

OAI22xp5_ASAP7_75t_L g3280 ( 
.A1(n_3177),
.A2(n_287),
.B1(n_284),
.B2(n_286),
.Y(n_3280)
);

BUFx2_ASAP7_75t_SL g3281 ( 
.A(n_2606),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_2942),
.B(n_686),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_2643),
.A2(n_286),
.B(n_287),
.Y(n_3283)
);

O2A1O1Ixp33_ASAP7_75t_L g3284 ( 
.A1(n_3046),
.A2(n_290),
.B(n_288),
.C(n_289),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2731),
.Y(n_3285)
);

NOR2xp33_ASAP7_75t_SL g3286 ( 
.A(n_2934),
.B(n_3062),
.Y(n_3286)
);

AND2x4_ASAP7_75t_L g3287 ( 
.A(n_2805),
.B(n_288),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_2842),
.A2(n_288),
.B(n_290),
.Y(n_3288)
);

BUFx2_ASAP7_75t_L g3289 ( 
.A(n_2700),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2810),
.B(n_290),
.Y(n_3290)
);

AOI21xp5_ASAP7_75t_L g3291 ( 
.A1(n_2730),
.A2(n_291),
.B(n_292),
.Y(n_3291)
);

AOI21x1_ASAP7_75t_L g3292 ( 
.A1(n_2687),
.A2(n_2713),
.B(n_2677),
.Y(n_3292)
);

AOI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_3061),
.A2(n_294),
.B1(n_291),
.B2(n_293),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_2599),
.A2(n_291),
.B(n_293),
.Y(n_3294)
);

BUFx6f_ASAP7_75t_L g3295 ( 
.A(n_2728),
.Y(n_3295)
);

INVxp67_ASAP7_75t_L g3296 ( 
.A(n_3129),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2767),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_SL g3298 ( 
.A(n_2942),
.B(n_687),
.Y(n_3298)
);

BUFx12f_ASAP7_75t_L g3299 ( 
.A(n_3101),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_2922),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2768),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_2603),
.A2(n_2620),
.B(n_2605),
.Y(n_3302)
);

NOR2xp33_ASAP7_75t_L g3303 ( 
.A(n_2583),
.B(n_2737),
.Y(n_3303)
);

AOI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_2626),
.A2(n_293),
.B(n_294),
.Y(n_3304)
);

O2A1O1Ixp33_ASAP7_75t_L g3305 ( 
.A1(n_3050),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_2930),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_2612),
.B(n_295),
.Y(n_3307)
);

NOR2xp33_ASAP7_75t_L g3308 ( 
.A(n_2666),
.B(n_295),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_2943),
.Y(n_3309)
);

INVxp67_ASAP7_75t_L g3310 ( 
.A(n_3161),
.Y(n_3310)
);

NOR2x1_ASAP7_75t_L g3311 ( 
.A(n_2700),
.B(n_296),
.Y(n_3311)
);

OR2x6_ASAP7_75t_L g3312 ( 
.A(n_2700),
.B(n_297),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_2625),
.B(n_297),
.Y(n_3313)
);

NAND2x1p5_ASAP7_75t_L g3314 ( 
.A(n_3062),
.B(n_298),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_SL g3315 ( 
.A(n_2942),
.B(n_687),
.Y(n_3315)
);

OAI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_2997),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_3316)
);

NOR3xp33_ASAP7_75t_L g3317 ( 
.A(n_3005),
.B(n_299),
.C(n_300),
.Y(n_3317)
);

CKINVDCx20_ASAP7_75t_R g3318 ( 
.A(n_2867),
.Y(n_3318)
);

NOR2xp33_ASAP7_75t_SL g3319 ( 
.A(n_3079),
.B(n_299),
.Y(n_3319)
);

AND2x4_ASAP7_75t_L g3320 ( 
.A(n_2564),
.B(n_300),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2819),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_2640),
.B(n_301),
.Y(n_3322)
);

NOR2xp33_ASAP7_75t_L g3323 ( 
.A(n_2833),
.B(n_302),
.Y(n_3323)
);

A2O1A1Ixp33_ASAP7_75t_L g3324 ( 
.A1(n_2871),
.A2(n_304),
.B(n_302),
.C(n_303),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_SL g3325 ( 
.A(n_2849),
.B(n_688),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_2619),
.Y(n_3326)
);

OAI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_2792),
.A2(n_302),
.B(n_303),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_2652),
.Y(n_3328)
);

OAI21xp33_ASAP7_75t_L g3329 ( 
.A1(n_2595),
.A2(n_304),
.B(n_306),
.Y(n_3329)
);

OAI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_2997),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_3330)
);

A2O1A1Ixp33_ASAP7_75t_L g3331 ( 
.A1(n_2721),
.A2(n_308),
.B(n_306),
.C(n_307),
.Y(n_3331)
);

BUFx6f_ASAP7_75t_L g3332 ( 
.A(n_2728),
.Y(n_3332)
);

AOI21xp5_ASAP7_75t_L g3333 ( 
.A1(n_2826),
.A2(n_308),
.B(n_309),
.Y(n_3333)
);

INVxp67_ASAP7_75t_L g3334 ( 
.A(n_3093),
.Y(n_3334)
);

A2O1A1Ixp33_ASAP7_75t_L g3335 ( 
.A1(n_2724),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2691),
.Y(n_3336)
);

A2O1A1Ixp33_ASAP7_75t_SL g3337 ( 
.A1(n_2607),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_2602),
.B(n_310),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_L g3339 ( 
.A(n_2856),
.B(n_2776),
.Y(n_3339)
);

INVx3_ASAP7_75t_L g3340 ( 
.A(n_3079),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_2602),
.B(n_312),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_2813),
.B(n_312),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_3093),
.B(n_688),
.Y(n_3343)
);

A2O1A1Ixp33_ASAP7_75t_L g3344 ( 
.A1(n_2784),
.A2(n_2785),
.B(n_2812),
.C(n_2806),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2692),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_2885),
.B(n_312),
.Y(n_3346)
);

AOI22xp5_ASAP7_75t_L g3347 ( 
.A1(n_2579),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_3347)
);

NOR2xp33_ASAP7_75t_L g3348 ( 
.A(n_2892),
.B(n_313),
.Y(n_3348)
);

O2A1O1Ixp33_ASAP7_75t_L g3349 ( 
.A1(n_2803),
.A2(n_316),
.B(n_313),
.C(n_314),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_2970),
.Y(n_3350)
);

OA22x2_ASAP7_75t_L g3351 ( 
.A1(n_2850),
.A2(n_317),
.B1(n_314),
.B2(n_316),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_2823),
.B(n_316),
.Y(n_3352)
);

CKINVDCx20_ASAP7_75t_R g3353 ( 
.A(n_3057),
.Y(n_3353)
);

BUFx12f_ASAP7_75t_L g3354 ( 
.A(n_2931),
.Y(n_3354)
);

A2O1A1Ixp33_ASAP7_75t_L g3355 ( 
.A1(n_2814),
.A2(n_319),
.B(n_317),
.C(n_318),
.Y(n_3355)
);

O2A1O1Ixp33_ASAP7_75t_L g3356 ( 
.A1(n_2807),
.A2(n_319),
.B(n_317),
.C(n_318),
.Y(n_3356)
);

HB1xp67_ASAP7_75t_L g3357 ( 
.A(n_2681),
.Y(n_3357)
);

O2A1O1Ixp5_ASAP7_75t_SL g3358 ( 
.A1(n_2693),
.A2(n_690),
.B(n_691),
.C(n_689),
.Y(n_3358)
);

AOI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_2740),
.A2(n_318),
.B(n_319),
.Y(n_3359)
);

INVx2_ASAP7_75t_SL g3360 ( 
.A(n_3107),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_2706),
.Y(n_3361)
);

INVx4_ASAP7_75t_L g3362 ( 
.A(n_2616),
.Y(n_3362)
);

AOI21xp5_ASAP7_75t_L g3363 ( 
.A1(n_2679),
.A2(n_321),
.B(n_322),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_2869),
.B(n_321),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2772),
.Y(n_3365)
);

BUFx8_ASAP7_75t_SL g3366 ( 
.A(n_2678),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_2637),
.B(n_321),
.Y(n_3367)
);

INVx3_ASAP7_75t_L g3368 ( 
.A(n_3107),
.Y(n_3368)
);

OAI21x1_ASAP7_75t_L g3369 ( 
.A1(n_2670),
.A2(n_322),
.B(n_323),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_2702),
.B(n_323),
.Y(n_3370)
);

AOI21x1_ASAP7_75t_L g3371 ( 
.A1(n_3071),
.A2(n_323),
.B(n_324),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_2964),
.B(n_324),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_2972),
.Y(n_3373)
);

O2A1O1Ixp33_ASAP7_75t_L g3374 ( 
.A1(n_2811),
.A2(n_3130),
.B(n_2876),
.C(n_2780),
.Y(n_3374)
);

AOI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_2689),
.A2(n_324),
.B(n_325),
.Y(n_3375)
);

BUFx12f_ASAP7_75t_L g3376 ( 
.A(n_3010),
.Y(n_3376)
);

OAI22xp5_ASAP7_75t_L g3377 ( 
.A1(n_2739),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_3377)
);

AOI22xp5_ASAP7_75t_L g3378 ( 
.A1(n_2789),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_3378)
);

CKINVDCx16_ASAP7_75t_R g3379 ( 
.A(n_2729),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_2919),
.Y(n_3380)
);

BUFx6f_ASAP7_75t_L g3381 ( 
.A(n_2728),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_2668),
.B(n_326),
.Y(n_3382)
);

INVx1_ASAP7_75t_SL g3383 ( 
.A(n_2584),
.Y(n_3383)
);

A2O1A1Ixp33_ASAP7_75t_L g3384 ( 
.A1(n_2824),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_3384)
);

NOR2xp33_ASAP7_75t_R g3385 ( 
.A(n_2782),
.B(n_329),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_2617),
.B(n_329),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2936),
.Y(n_3387)
);

NOR2x1_ASAP7_75t_SL g3388 ( 
.A(n_2850),
.B(n_330),
.Y(n_3388)
);

BUFx6f_ASAP7_75t_L g3389 ( 
.A(n_2756),
.Y(n_3389)
);

OAI21xp33_ASAP7_75t_SL g3390 ( 
.A1(n_2739),
.A2(n_330),
.B(n_331),
.Y(n_3390)
);

OAI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_2636),
.A2(n_330),
.B(n_331),
.Y(n_3391)
);

NOR2xp33_ASAP7_75t_SL g3392 ( 
.A(n_3157),
.B(n_332),
.Y(n_3392)
);

O2A1O1Ixp33_ASAP7_75t_L g3393 ( 
.A1(n_2747),
.A2(n_334),
.B(n_332),
.C(n_333),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_2594),
.B(n_332),
.Y(n_3394)
);

BUFx3_ASAP7_75t_L g3395 ( 
.A(n_3016),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_2594),
.B(n_334),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_2797),
.B(n_335),
.Y(n_3397)
);

AOI22xp5_ASAP7_75t_L g3398 ( 
.A1(n_2788),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_3398)
);

OR2x6_ASAP7_75t_L g3399 ( 
.A(n_3108),
.B(n_335),
.Y(n_3399)
);

AOI22xp33_ASAP7_75t_L g3400 ( 
.A1(n_2850),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_3400)
);

NOR2xp67_ASAP7_75t_L g3401 ( 
.A(n_3104),
.B(n_336),
.Y(n_3401)
);

O2A1O1Ixp5_ASAP7_75t_L g3402 ( 
.A1(n_2887),
.A2(n_340),
.B(n_338),
.C(n_339),
.Y(n_3402)
);

A2O1A1Ixp33_ASAP7_75t_L g3403 ( 
.A1(n_2825),
.A2(n_340),
.B(n_338),
.C(n_339),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_2991),
.Y(n_3404)
);

AOI21xp5_ASAP7_75t_L g3405 ( 
.A1(n_2748),
.A2(n_340),
.B(n_341),
.Y(n_3405)
);

AND2x4_ASAP7_75t_L g3406 ( 
.A(n_3104),
.B(n_341),
.Y(n_3406)
);

AND2x2_ASAP7_75t_L g3407 ( 
.A(n_3007),
.B(n_2963),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_SL g3408 ( 
.A(n_2926),
.B(n_689),
.Y(n_3408)
);

OAI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_2752),
.A2(n_344),
.B1(n_341),
.B2(n_342),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_2985),
.B(n_342),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_2937),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_2799),
.B(n_342),
.Y(n_3412)
);

AOI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_2703),
.A2(n_344),
.B(n_345),
.Y(n_3413)
);

O2A1O1Ixp5_ASAP7_75t_SL g3414 ( 
.A1(n_2917),
.A2(n_2732),
.B(n_2696),
.C(n_2688),
.Y(n_3414)
);

AND2x2_ASAP7_75t_L g3415 ( 
.A(n_3059),
.B(n_344),
.Y(n_3415)
);

AOI21xp5_ASAP7_75t_L g3416 ( 
.A1(n_2704),
.A2(n_345),
.B(n_346),
.Y(n_3416)
);

OAI22xp5_ASAP7_75t_L g3417 ( 
.A1(n_2752),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_3417)
);

AOI21xp5_ASAP7_75t_L g3418 ( 
.A1(n_2709),
.A2(n_346),
.B(n_347),
.Y(n_3418)
);

AOI21xp5_ASAP7_75t_L g3419 ( 
.A1(n_2710),
.A2(n_347),
.B(n_348),
.Y(n_3419)
);

OAI22xp5_ASAP7_75t_L g3420 ( 
.A1(n_3039),
.A2(n_3147),
.B1(n_2618),
.B2(n_2820),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_2995),
.Y(n_3421)
);

AOI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_2615),
.A2(n_348),
.B(n_349),
.Y(n_3422)
);

HB1xp67_ASAP7_75t_L g3423 ( 
.A(n_3131),
.Y(n_3423)
);

NOR2xp33_ASAP7_75t_L g3424 ( 
.A(n_2621),
.B(n_349),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_2938),
.Y(n_3425)
);

OAI22x1_ASAP7_75t_L g3426 ( 
.A1(n_3039),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_2903),
.B(n_350),
.Y(n_3427)
);

AND2x4_ASAP7_75t_L g3428 ( 
.A(n_2865),
.B(n_350),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2941),
.Y(n_3429)
);

AND2x4_ASAP7_75t_L g3430 ( 
.A(n_2908),
.B(n_351),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_2808),
.B(n_351),
.Y(n_3431)
);

INVx2_ASAP7_75t_L g3432 ( 
.A(n_3002),
.Y(n_3432)
);

AOI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_2838),
.A2(n_352),
.B(n_353),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_2672),
.A2(n_354),
.B(n_355),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_2829),
.B(n_354),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_2840),
.B(n_354),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_2841),
.B(n_355),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_2673),
.A2(n_355),
.B(n_356),
.Y(n_3438)
);

HB1xp67_ASAP7_75t_L g3439 ( 
.A(n_2660),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_2877),
.B(n_356),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_2836),
.B(n_356),
.Y(n_3441)
);

OR2x2_ASAP7_75t_L g3442 ( 
.A(n_2609),
.B(n_2570),
.Y(n_3442)
);

INVx3_ASAP7_75t_L g3443 ( 
.A(n_3157),
.Y(n_3443)
);

AOI22x1_ASAP7_75t_L g3444 ( 
.A1(n_2855),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_3444)
);

INVx4_ASAP7_75t_L g3445 ( 
.A(n_3022),
.Y(n_3445)
);

INVx2_ASAP7_75t_SL g3446 ( 
.A(n_2659),
.Y(n_3446)
);

AOI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_2676),
.A2(n_357),
.B(n_358),
.Y(n_3447)
);

OAI21x1_ASAP7_75t_L g3448 ( 
.A1(n_2925),
.A2(n_357),
.B(n_358),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_2926),
.B(n_690),
.Y(n_3449)
);

OAI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_2567),
.A2(n_360),
.B(n_361),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3031),
.Y(n_3451)
);

OAI22xp5_ASAP7_75t_L g3452 ( 
.A1(n_3147),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_3452)
);

AOI21xp33_ASAP7_75t_L g3453 ( 
.A1(n_2863),
.A2(n_361),
.B(n_362),
.Y(n_3453)
);

A2O1A1Ixp33_ASAP7_75t_L g3454 ( 
.A1(n_2827),
.A2(n_364),
.B(n_362),
.C(n_363),
.Y(n_3454)
);

AND2x2_ASAP7_75t_L g3455 ( 
.A(n_2634),
.B(n_363),
.Y(n_3455)
);

NOR3xp33_ASAP7_75t_SL g3456 ( 
.A(n_2675),
.B(n_363),
.C(n_364),
.Y(n_3456)
);

AOI22xp33_ASAP7_75t_L g3457 ( 
.A1(n_2837),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_3457)
);

BUFx2_ASAP7_75t_L g3458 ( 
.A(n_2609),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_L g3459 ( 
.A(n_2566),
.B(n_365),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_2674),
.A2(n_365),
.B(n_366),
.Y(n_3460)
);

NAND2xp33_ASAP7_75t_L g3461 ( 
.A(n_2926),
.B(n_366),
.Y(n_3461)
);

NOR2xp33_ASAP7_75t_L g3462 ( 
.A(n_2569),
.B(n_367),
.Y(n_3462)
);

A2O1A1Ixp33_ASAP7_75t_L g3463 ( 
.A1(n_3006),
.A2(n_369),
.B(n_367),
.C(n_368),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_2954),
.B(n_368),
.Y(n_3464)
);

INVx4_ASAP7_75t_L g3465 ( 
.A(n_2609),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_2956),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_2684),
.A2(n_369),
.B(n_370),
.Y(n_3467)
);

OAI22xp5_ASAP7_75t_SL g3468 ( 
.A1(n_2844),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_3468)
);

A2O1A1Ixp33_ASAP7_75t_SL g3469 ( 
.A1(n_2928),
.A2(n_372),
.B(n_370),
.C(n_371),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_2613),
.A2(n_2614),
.B(n_2771),
.Y(n_3470)
);

AOI221xp5_ASAP7_75t_L g3471 ( 
.A1(n_2977),
.A2(n_374),
.B1(n_371),
.B2(n_373),
.C(n_375),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3048),
.Y(n_3472)
);

O2A1O1Ixp33_ASAP7_75t_L g3473 ( 
.A1(n_2948),
.A2(n_375),
.B(n_373),
.C(n_374),
.Y(n_3473)
);

OAI22xp5_ASAP7_75t_SL g3474 ( 
.A1(n_2697),
.A2(n_376),
.B1(n_373),
.B2(n_375),
.Y(n_3474)
);

BUFx6f_ASAP7_75t_L g3475 ( 
.A(n_2756),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_2958),
.B(n_376),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3070),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_2962),
.B(n_3187),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_2965),
.B(n_377),
.Y(n_3479)
);

A2O1A1Ixp33_ASAP7_75t_L g3480 ( 
.A1(n_3069),
.A2(n_379),
.B(n_377),
.C(n_378),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_2967),
.B(n_377),
.Y(n_3481)
);

AOI21xp5_ASAP7_75t_L g3482 ( 
.A1(n_2773),
.A2(n_378),
.B(n_379),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_L g3483 ( 
.A(n_2694),
.B(n_380),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_2969),
.B(n_380),
.Y(n_3484)
);

NOR2xp33_ASAP7_75t_L g3485 ( 
.A(n_2563),
.B(n_380),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_2974),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_2975),
.Y(n_3487)
);

AOI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_2786),
.A2(n_381),
.B(n_382),
.Y(n_3488)
);

OR2x6_ASAP7_75t_L g3489 ( 
.A(n_2565),
.B(n_381),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_2982),
.Y(n_3490)
);

AOI21xp5_ASAP7_75t_L g3491 ( 
.A1(n_2790),
.A2(n_381),
.B(n_382),
.Y(n_3491)
);

A2O1A1Ixp33_ASAP7_75t_SL g3492 ( 
.A1(n_2857),
.A2(n_385),
.B(n_383),
.C(n_384),
.Y(n_3492)
);

CKINVDCx8_ASAP7_75t_R g3493 ( 
.A(n_2659),
.Y(n_3493)
);

INVx3_ASAP7_75t_SL g3494 ( 
.A(n_2714),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_2983),
.Y(n_3495)
);

CKINVDCx5p33_ASAP7_75t_R g3496 ( 
.A(n_2816),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_2992),
.B(n_2998),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3088),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3001),
.B(n_383),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3008),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3023),
.B(n_384),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3033),
.B(n_384),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_2815),
.A2(n_385),
.B(n_386),
.Y(n_3503)
);

AOI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_2894),
.A2(n_386),
.B(n_387),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_3120),
.Y(n_3505)
);

INVx1_ASAP7_75t_SL g3506 ( 
.A(n_2699),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3034),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_SL g3508 ( 
.A(n_2926),
.B(n_2618),
.Y(n_3508)
);

AOI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_2986),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_SL g3510 ( 
.A(n_2926),
.B(n_691),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3036),
.B(n_387),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_3186),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_SL g3513 ( 
.A(n_2575),
.B(n_692),
.Y(n_3513)
);

AOI21x1_ASAP7_75t_L g3514 ( 
.A1(n_3096),
.A2(n_388),
.B(n_389),
.Y(n_3514)
);

OAI21x1_ASAP7_75t_L g3515 ( 
.A1(n_2987),
.A2(n_388),
.B(n_389),
.Y(n_3515)
);

OAI21xp33_ASAP7_75t_L g3516 ( 
.A1(n_2861),
.A2(n_389),
.B(n_390),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3041),
.B(n_390),
.Y(n_3517)
);

OR2x6_ASAP7_75t_L g3518 ( 
.A(n_3194),
.B(n_390),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3043),
.Y(n_3519)
);

HB1xp67_ASAP7_75t_L g3520 ( 
.A(n_2769),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_SL g3521 ( 
.A(n_2575),
.B(n_692),
.Y(n_3521)
);

CKINVDCx5p33_ASAP7_75t_R g3522 ( 
.A(n_2783),
.Y(n_3522)
);

NAND3xp33_ASAP7_75t_SL g3523 ( 
.A(n_2793),
.B(n_2820),
.C(n_2682),
.Y(n_3523)
);

INVxp67_ASAP7_75t_L g3524 ( 
.A(n_2940),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3045),
.B(n_391),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_SL g3526 ( 
.A(n_2575),
.B(n_2577),
.Y(n_3526)
);

NAND3x1_ASAP7_75t_L g3527 ( 
.A(n_2888),
.B(n_391),
.C(n_392),
.Y(n_3527)
);

INVx1_ASAP7_75t_SL g3528 ( 
.A(n_2765),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_2591),
.B(n_391),
.Y(n_3529)
);

OAI22xp33_ASAP7_75t_SL g3530 ( 
.A1(n_2927),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_3530)
);

BUFx6f_ASAP7_75t_L g3531 ( 
.A(n_2756),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3049),
.B(n_392),
.Y(n_3532)
);

AND2x2_ASAP7_75t_L g3533 ( 
.A(n_2591),
.B(n_393),
.Y(n_3533)
);

BUFx6f_ASAP7_75t_L g3534 ( 
.A(n_2577),
.Y(n_3534)
);

O2A1O1Ixp5_ASAP7_75t_L g3535 ( 
.A1(n_2686),
.A2(n_395),
.B(n_393),
.C(n_394),
.Y(n_3535)
);

AND2x2_ASAP7_75t_L g3536 ( 
.A(n_3019),
.B(n_395),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3056),
.B(n_396),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3060),
.Y(n_3538)
);

BUFx2_ASAP7_75t_L g3539 ( 
.A(n_2783),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_SL g3540 ( 
.A(n_2577),
.B(n_693),
.Y(n_3540)
);

NOR3xp33_ASAP7_75t_SL g3541 ( 
.A(n_3094),
.B(n_396),
.C(n_397),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_SL g3542 ( 
.A(n_2588),
.B(n_693),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_R g3543 ( 
.A(n_2787),
.B(n_396),
.Y(n_3543)
);

INVx1_ASAP7_75t_SL g3544 ( 
.A(n_2665),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3064),
.B(n_397),
.Y(n_3545)
);

AOI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3038),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_3546)
);

OR2x6_ASAP7_75t_L g3547 ( 
.A(n_2665),
.B(n_398),
.Y(n_3547)
);

AOI21xp5_ASAP7_75t_L g3548 ( 
.A1(n_2562),
.A2(n_398),
.B(n_399),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_3195),
.Y(n_3549)
);

NOR2x1_ASAP7_75t_L g3550 ( 
.A(n_2843),
.B(n_399),
.Y(n_3550)
);

OAI21x1_ASAP7_75t_L g3551 ( 
.A1(n_2830),
.A2(n_400),
.B(n_401),
.Y(n_3551)
);

OAI22xp5_ASAP7_75t_L g3552 ( 
.A1(n_3067),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3068),
.B(n_401),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_2630),
.Y(n_3554)
);

OR2x6_ASAP7_75t_L g3555 ( 
.A(n_2734),
.B(n_2843),
.Y(n_3555)
);

AND2x4_ASAP7_75t_L g3556 ( 
.A(n_2623),
.B(n_402),
.Y(n_3556)
);

AOI22xp5_ASAP7_75t_L g3557 ( 
.A1(n_3087),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_3557)
);

NOR2xp33_ASAP7_75t_L g3558 ( 
.A(n_2890),
.B(n_403),
.Y(n_3558)
);

OR2x6_ASAP7_75t_L g3559 ( 
.A(n_2734),
.B(n_404),
.Y(n_3559)
);

NOR2xp67_ASAP7_75t_SL g3560 ( 
.A(n_3197),
.B(n_404),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3150),
.B(n_405),
.Y(n_3561)
);

NOR3xp33_ASAP7_75t_SL g3562 ( 
.A(n_2904),
.B(n_406),
.C(n_407),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3082),
.B(n_406),
.Y(n_3563)
);

BUFx2_ASAP7_75t_L g3564 ( 
.A(n_2940),
.Y(n_3564)
);

AOI22x1_ASAP7_75t_L g3565 ( 
.A1(n_2628),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3086),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3089),
.Y(n_3567)
);

BUFx3_ASAP7_75t_L g3568 ( 
.A(n_2723),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3102),
.B(n_408),
.Y(n_3569)
);

HB1xp67_ASAP7_75t_L g3570 ( 
.A(n_2837),
.Y(n_3570)
);

INVx1_ASAP7_75t_SL g3571 ( 
.A(n_2750),
.Y(n_3571)
);

INVx1_ASAP7_75t_SL g3572 ( 
.A(n_2715),
.Y(n_3572)
);

AOI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_2802),
.A2(n_408),
.B(n_409),
.Y(n_3573)
);

AND2x4_ASAP7_75t_L g3574 ( 
.A(n_2623),
.B(n_409),
.Y(n_3574)
);

OAI22xp5_ASAP7_75t_L g3575 ( 
.A1(n_3103),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3119),
.B(n_410),
.Y(n_3576)
);

NOR2xp67_ASAP7_75t_L g3577 ( 
.A(n_3166),
.B(n_410),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3122),
.B(n_411),
.Y(n_3578)
);

NOR2xp67_ASAP7_75t_L g3579 ( 
.A(n_3167),
.B(n_411),
.Y(n_3579)
);

BUFx2_ASAP7_75t_L g3580 ( 
.A(n_2787),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_3185),
.B(n_412),
.Y(n_3581)
);

A2O1A1Ixp33_ASAP7_75t_L g3582 ( 
.A1(n_3125),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_3582)
);

OAI21xp5_ASAP7_75t_L g3583 ( 
.A1(n_2568),
.A2(n_412),
.B(n_413),
.Y(n_3583)
);

NAND3xp33_ASAP7_75t_L g3584 ( 
.A(n_2601),
.B(n_3081),
.C(n_2741),
.Y(n_3584)
);

AOI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_2866),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_3585)
);

AO32x1_ASAP7_75t_L g3586 ( 
.A1(n_2902),
.A2(n_416),
.A3(n_414),
.B1(n_415),
.B2(n_417),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3123),
.Y(n_3587)
);

AO22x1_ASAP7_75t_L g3588 ( 
.A1(n_2794),
.A2(n_418),
.B1(n_416),
.B2(n_417),
.Y(n_3588)
);

OAI21x1_ASAP7_75t_L g3589 ( 
.A1(n_2915),
.A2(n_418),
.B(n_419),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_2633),
.B(n_2572),
.Y(n_3590)
);

AOI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_2638),
.A2(n_418),
.B(n_419),
.Y(n_3591)
);

BUFx3_ASAP7_75t_L g3592 ( 
.A(n_2715),
.Y(n_3592)
);

A2O1A1Ixp33_ASAP7_75t_L g3593 ( 
.A1(n_2711),
.A2(n_421),
.B(n_419),
.C(n_420),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_2635),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_2642),
.A2(n_420),
.B(n_421),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_SL g3596 ( 
.A(n_2588),
.B(n_694),
.Y(n_3596)
);

NOR2xp33_ASAP7_75t_SL g3597 ( 
.A(n_2588),
.B(n_420),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3128),
.B(n_421),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3137),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3146),
.Y(n_3600)
);

CKINVDCx8_ASAP7_75t_R g3601 ( 
.A(n_2895),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3162),
.B(n_3190),
.Y(n_3602)
);

HB1xp67_ASAP7_75t_L g3603 ( 
.A(n_2650),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_2695),
.B(n_2939),
.Y(n_3604)
);

OAI21x1_ASAP7_75t_L g3605 ( 
.A1(n_2916),
.A2(n_422),
.B(n_423),
.Y(n_3605)
);

AOI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_2690),
.A2(n_422),
.B(n_423),
.Y(n_3606)
);

OAI22xp5_ASAP7_75t_L g3607 ( 
.A1(n_3174),
.A2(n_425),
.B1(n_422),
.B2(n_424),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3175),
.Y(n_3608)
);

NAND2x1p5_ASAP7_75t_L g3609 ( 
.A(n_2695),
.B(n_424),
.Y(n_3609)
);

INVxp67_ASAP7_75t_L g3610 ( 
.A(n_2832),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_2851),
.A2(n_424),
.B(n_425),
.Y(n_3611)
);

BUFx6f_ASAP7_75t_L g3612 ( 
.A(n_2695),
.Y(n_3612)
);

AND2x2_ASAP7_75t_L g3613 ( 
.A(n_2633),
.B(n_425),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_2653),
.Y(n_3614)
);

A2O1A1Ixp33_ASAP7_75t_SL g3615 ( 
.A1(n_2907),
.A2(n_428),
.B(n_426),
.C(n_427),
.Y(n_3615)
);

NAND2x1p5_ASAP7_75t_L g3616 ( 
.A(n_2939),
.B(n_426),
.Y(n_3616)
);

BUFx3_ASAP7_75t_L g3617 ( 
.A(n_2883),
.Y(n_3617)
);

OAI21x1_ASAP7_75t_L g3618 ( 
.A1(n_3126),
.A2(n_426),
.B(n_427),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_2953),
.B(n_427),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_2661),
.Y(n_3620)
);

NOR2xp33_ASAP7_75t_L g3621 ( 
.A(n_2901),
.B(n_428),
.Y(n_3621)
);

INVx3_ASAP7_75t_L g3622 ( 
.A(n_2909),
.Y(n_3622)
);

INVx4_ASAP7_75t_L g3623 ( 
.A(n_2939),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3179),
.B(n_428),
.Y(n_3624)
);

BUFx2_ASAP7_75t_L g3625 ( 
.A(n_2993),
.Y(n_3625)
);

OAI21xp33_ASAP7_75t_SL g3626 ( 
.A1(n_2746),
.A2(n_429),
.B(n_430),
.Y(n_3626)
);

AOI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_2658),
.A2(n_430),
.B(n_431),
.Y(n_3627)
);

INVx3_ASAP7_75t_SL g3628 ( 
.A(n_2906),
.Y(n_3628)
);

OAI22xp5_ASAP7_75t_L g3629 ( 
.A1(n_3181),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_3629)
);

INVx1_ASAP7_75t_SL g3630 ( 
.A(n_2891),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3182),
.Y(n_3631)
);

AOI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_2592),
.A2(n_2561),
.B(n_2798),
.Y(n_3632)
);

BUFx6f_ASAP7_75t_L g3633 ( 
.A(n_2993),
.Y(n_3633)
);

BUFx3_ASAP7_75t_L g3634 ( 
.A(n_2993),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_3013),
.B(n_431),
.Y(n_3635)
);

AOI22xp5_ASAP7_75t_L g3636 ( 
.A1(n_2960),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_3636)
);

AOI21x1_ASAP7_75t_L g3637 ( 
.A1(n_2722),
.A2(n_433),
.B(n_434),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_2663),
.Y(n_3638)
);

NOR2xp33_ASAP7_75t_SL g3639 ( 
.A(n_3084),
.B(n_433),
.Y(n_3639)
);

NOR2xp33_ASAP7_75t_L g3640 ( 
.A(n_2582),
.B(n_435),
.Y(n_3640)
);

OAI21x1_ASAP7_75t_L g3641 ( 
.A1(n_2671),
.A2(n_436),
.B(n_437),
.Y(n_3641)
);

AOI21xp5_ASAP7_75t_L g3642 ( 
.A1(n_2800),
.A2(n_436),
.B(n_437),
.Y(n_3642)
);

AND2x2_ASAP7_75t_L g3643 ( 
.A(n_3136),
.B(n_436),
.Y(n_3643)
);

OAI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_2878),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_3644)
);

AND2x4_ASAP7_75t_L g3645 ( 
.A(n_2701),
.B(n_438),
.Y(n_3645)
);

AOI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_2597),
.A2(n_438),
.B(n_439),
.Y(n_3646)
);

AND2x4_ASAP7_75t_L g3647 ( 
.A(n_2701),
.B(n_440),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_2664),
.Y(n_3648)
);

AOI22xp5_ASAP7_75t_L g3649 ( 
.A1(n_2980),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_3649)
);

A2O1A1Ixp33_ASAP7_75t_L g3650 ( 
.A1(n_2835),
.A2(n_443),
.B(n_441),
.C(n_442),
.Y(n_3650)
);

A2O1A1Ixp33_ASAP7_75t_SL g3651 ( 
.A1(n_3024),
.A2(n_443),
.B(n_441),
.C(n_442),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_SL g3652 ( 
.A(n_3084),
.B(n_3091),
.Y(n_3652)
);

BUFx6f_ASAP7_75t_L g3653 ( 
.A(n_3084),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_2632),
.B(n_445),
.Y(n_3654)
);

AOI21xp5_ASAP7_75t_L g3655 ( 
.A1(n_2973),
.A2(n_446),
.B(n_447),
.Y(n_3655)
);

A2O1A1Ixp33_ASAP7_75t_L g3656 ( 
.A1(n_2698),
.A2(n_448),
.B(n_446),
.C(n_447),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_2775),
.B(n_448),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_2641),
.B(n_448),
.Y(n_3658)
);

AOI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3004),
.A2(n_3011),
.B1(n_3037),
.B2(n_3015),
.Y(n_3659)
);

BUFx6f_ASAP7_75t_L g3660 ( 
.A(n_3091),
.Y(n_3660)
);

AOI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_3026),
.A2(n_449),
.B(n_450),
.Y(n_3661)
);

O2A1O1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_3028),
.A2(n_451),
.B(n_449),
.C(n_450),
.Y(n_3662)
);

AO32x2_ASAP7_75t_L g3663 ( 
.A1(n_2959),
.A2(n_3066),
.A3(n_3139),
.B1(n_3121),
.B2(n_2994),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_2622),
.B(n_449),
.Y(n_3664)
);

NOR2x1_ASAP7_75t_SL g3665 ( 
.A(n_3091),
.B(n_3098),
.Y(n_3665)
);

INVx3_ASAP7_75t_L g3666 ( 
.A(n_2909),
.Y(n_3666)
);

OAI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_2580),
.A2(n_450),
.B(n_452),
.Y(n_3667)
);

AOI22xp5_ASAP7_75t_L g3668 ( 
.A1(n_3051),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_3668)
);

AOI22xp5_ASAP7_75t_L g3669 ( 
.A1(n_3077),
.A2(n_3090),
.B1(n_3163),
.B2(n_3110),
.Y(n_3669)
);

AO21x1_ASAP7_75t_L g3670 ( 
.A1(n_2845),
.A2(n_696),
.B(n_694),
.Y(n_3670)
);

NOR3xp33_ASAP7_75t_L g3671 ( 
.A(n_3040),
.B(n_452),
.C(n_453),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_2735),
.Y(n_3672)
);

AOI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_2587),
.A2(n_453),
.B(n_454),
.Y(n_3673)
);

INVxp67_ASAP7_75t_L g3674 ( 
.A(n_2781),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_2573),
.B(n_454),
.Y(n_3675)
);

NAND3xp33_ASAP7_75t_SL g3676 ( 
.A(n_3065),
.B(n_455),
.C(n_456),
.Y(n_3676)
);

O2A1O1Ixp33_ASAP7_75t_L g3677 ( 
.A1(n_3073),
.A2(n_458),
.B(n_455),
.C(n_457),
.Y(n_3677)
);

INVx1_ASAP7_75t_SL g3678 ( 
.A(n_2893),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_2749),
.Y(n_3679)
);

BUFx6f_ASAP7_75t_L g3680 ( 
.A(n_3098),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_2590),
.B(n_457),
.Y(n_3681)
);

CKINVDCx5p33_ASAP7_75t_R g3682 ( 
.A(n_2896),
.Y(n_3682)
);

CKINVDCx20_ASAP7_75t_R g3683 ( 
.A(n_3098),
.Y(n_3683)
);

OAI22xp5_ASAP7_75t_L g3684 ( 
.A1(n_2875),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_3684)
);

AOI222xp33_ASAP7_75t_L g3685 ( 
.A1(n_3141),
.A2(n_461),
.B1(n_463),
.B2(n_458),
.C1(n_459),
.C2(n_462),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_2593),
.B(n_461),
.Y(n_3686)
);

O2A1O1Ixp33_ASAP7_75t_L g3687 ( 
.A1(n_3127),
.A2(n_3145),
.B(n_2809),
.C(n_2791),
.Y(n_3687)
);

INVx3_ASAP7_75t_L g3688 ( 
.A(n_2968),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_2755),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_2596),
.B(n_461),
.Y(n_3690)
);

AOI21xp5_ASAP7_75t_L g3691 ( 
.A1(n_2629),
.A2(n_462),
.B(n_463),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_2761),
.Y(n_3692)
);

OAI22xp5_ASAP7_75t_L g3693 ( 
.A1(n_2762),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_SL g3694 ( 
.A(n_3132),
.B(n_697),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_SL g3695 ( 
.A(n_3132),
.B(n_698),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_SL g3696 ( 
.A(n_3132),
.B(n_464),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_2667),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_2725),
.B(n_464),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_2763),
.B(n_465),
.Y(n_3699)
);

AND2x6_ASAP7_75t_SL g3700 ( 
.A(n_2859),
.B(n_466),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3047),
.A2(n_2712),
.B(n_2839),
.Y(n_3701)
);

CKINVDCx5p33_ASAP7_75t_R g3702 ( 
.A(n_3172),
.Y(n_3702)
);

NAND2x1p5_ASAP7_75t_L g3703 ( 
.A(n_3138),
.B(n_466),
.Y(n_3703)
);

BUFx2_ASAP7_75t_L g3704 ( 
.A(n_3138),
.Y(n_3704)
);

NOR2xp33_ASAP7_75t_R g3705 ( 
.A(n_3138),
.B(n_3142),
.Y(n_3705)
);

A2O1A1Ixp33_ASAP7_75t_L g3706 ( 
.A1(n_2707),
.A2(n_468),
.B(n_466),
.C(n_467),
.Y(n_3706)
);

OAI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_2770),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_2821),
.A2(n_467),
.B(n_468),
.Y(n_3708)
);

NOR2xp33_ASAP7_75t_L g3709 ( 
.A(n_2578),
.B(n_469),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_2796),
.Y(n_3710)
);

NAND3xp33_ASAP7_75t_SL g3711 ( 
.A(n_2733),
.B(n_2779),
.C(n_2881),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_2905),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_SL g3713 ( 
.A(n_3142),
.B(n_698),
.Y(n_3713)
);

O2A1O1Ixp33_ASAP7_75t_L g3714 ( 
.A1(n_2924),
.A2(n_471),
.B(n_469),
.C(n_470),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_2581),
.B(n_471),
.Y(n_3715)
);

OAI22x1_ASAP7_75t_L g3716 ( 
.A1(n_2910),
.A2(n_2736),
.B1(n_2899),
.B2(n_2742),
.Y(n_3716)
);

INVx3_ASAP7_75t_L g3717 ( 
.A(n_2968),
.Y(n_3717)
);

OAI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_2817),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.Y(n_3718)
);

A2O1A1Ixp33_ASAP7_75t_L g3719 ( 
.A1(n_2717),
.A2(n_475),
.B(n_472),
.C(n_474),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_2872),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_2873),
.B(n_472),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_SL g3722 ( 
.A(n_3142),
.B(n_699),
.Y(n_3722)
);

OAI22xp5_ASAP7_75t_L g3723 ( 
.A1(n_2801),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_2822),
.Y(n_3724)
);

BUFx6f_ASAP7_75t_L g3725 ( 
.A(n_3155),
.Y(n_3725)
);

O2A1O1Ixp33_ASAP7_75t_L g3726 ( 
.A1(n_2933),
.A2(n_479),
.B(n_477),
.C(n_478),
.Y(n_3726)
);

OR2x6_ASAP7_75t_L g3727 ( 
.A(n_2884),
.B(n_478),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_2900),
.B(n_478),
.Y(n_3728)
);

INVxp67_ASAP7_75t_SL g3729 ( 
.A(n_3155),
.Y(n_3729)
);

NOR2xp33_ASAP7_75t_L g3730 ( 
.A(n_2912),
.B(n_479),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3180),
.Y(n_3731)
);

BUFx6f_ASAP7_75t_L g3732 ( 
.A(n_3155),
.Y(n_3732)
);

BUFx3_ASAP7_75t_L g3733 ( 
.A(n_3178),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3178),
.Y(n_3734)
);

BUFx2_ASAP7_75t_L g3735 ( 
.A(n_3178),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3207),
.Y(n_3736)
);

INVx3_ASAP7_75t_SL g3737 ( 
.A(n_3205),
.Y(n_3737)
);

AO31x2_ASAP7_75t_L g3738 ( 
.A1(n_3710),
.A2(n_2753),
.A3(n_2947),
.B(n_2944),
.Y(n_3738)
);

INVxp67_ASAP7_75t_L g3739 ( 
.A(n_3211),
.Y(n_3739)
);

NOR2xp33_ASAP7_75t_L g3740 ( 
.A(n_3628),
.B(n_2647),
.Y(n_3740)
);

OAI21x1_ASAP7_75t_L g3741 ( 
.A1(n_3292),
.A2(n_2685),
.B(n_2680),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3231),
.Y(n_3742)
);

AO31x2_ASAP7_75t_L g3743 ( 
.A1(n_3712),
.A2(n_3029),
.A3(n_3052),
.B(n_3000),
.Y(n_3743)
);

AOI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_3461),
.A2(n_2611),
.B(n_2655),
.Y(n_3744)
);

INVx2_ASAP7_75t_SL g3745 ( 
.A(n_3206),
.Y(n_3745)
);

OAI21x1_ASAP7_75t_L g3746 ( 
.A1(n_3268),
.A2(n_2766),
.B(n_2758),
.Y(n_3746)
);

BUFx3_ASAP7_75t_L g3747 ( 
.A(n_3277),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_3321),
.B(n_2718),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3346),
.B(n_2738),
.Y(n_3749)
);

CKINVDCx20_ASAP7_75t_R g3750 ( 
.A(n_3242),
.Y(n_3750)
);

O2A1O1Ixp33_ASAP7_75t_SL g3751 ( 
.A1(n_3230),
.A2(n_2918),
.B(n_2989),
.C(n_2981),
.Y(n_3751)
);

CKINVDCx5p33_ASAP7_75t_R g3752 ( 
.A(n_3262),
.Y(n_3752)
);

AOI21xp5_ASAP7_75t_L g3753 ( 
.A1(n_3632),
.A2(n_2611),
.B(n_2708),
.Y(n_3753)
);

AOI21xp5_ASAP7_75t_L g3754 ( 
.A1(n_3470),
.A2(n_3032),
.B(n_3027),
.Y(n_3754)
);

OAI21x1_ASAP7_75t_L g3755 ( 
.A1(n_3701),
.A2(n_2777),
.B(n_2774),
.Y(n_3755)
);

HB1xp67_ASAP7_75t_L g3756 ( 
.A(n_3439),
.Y(n_3756)
);

O2A1O1Ixp33_ASAP7_75t_L g3757 ( 
.A1(n_3530),
.A2(n_3072),
.B(n_3151),
.C(n_3075),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3303),
.B(n_2759),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3259),
.Y(n_3759)
);

INVx3_ASAP7_75t_SL g3760 ( 
.A(n_3362),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3265),
.Y(n_3761)
);

OAI21x1_ASAP7_75t_L g3762 ( 
.A1(n_3526),
.A2(n_2778),
.B(n_2979),
.Y(n_3762)
);

OAI21x1_ASAP7_75t_L g3763 ( 
.A1(n_3604),
.A2(n_3054),
.B(n_2979),
.Y(n_3763)
);

OA21x2_ASAP7_75t_L g3764 ( 
.A1(n_3448),
.A2(n_2913),
.B(n_2848),
.Y(n_3764)
);

NAND3xp33_ASAP7_75t_L g3765 ( 
.A(n_3456),
.B(n_3183),
.C(n_3156),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_3344),
.A2(n_3109),
.B(n_3058),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3300),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3306),
.Y(n_3768)
);

OAI21xp5_ASAP7_75t_L g3769 ( 
.A1(n_3414),
.A2(n_2870),
.B(n_2864),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3309),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3529),
.B(n_2882),
.Y(n_3771)
);

NAND2x1p5_ASAP7_75t_L g3772 ( 
.A(n_3214),
.B(n_3054),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3508),
.A2(n_2860),
.B(n_2914),
.Y(n_3773)
);

AND2x4_ASAP7_75t_L g3774 ( 
.A(n_3214),
.B(n_2719),
.Y(n_3774)
);

NOR2xp33_ASAP7_75t_L g3775 ( 
.A(n_3289),
.B(n_2648),
.Y(n_3775)
);

AOI22xp5_ASAP7_75t_L g3776 ( 
.A1(n_3420),
.A2(n_2801),
.B1(n_2705),
.B2(n_2745),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3533),
.B(n_2886),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3407),
.B(n_2586),
.Y(n_3778)
);

OAI21x1_ASAP7_75t_L g3779 ( 
.A1(n_3652),
.A2(n_3117),
.B(n_3080),
.Y(n_3779)
);

AO21x2_ASAP7_75t_L g3780 ( 
.A1(n_3222),
.A2(n_3159),
.B(n_2751),
.Y(n_3780)
);

BUFx6f_ASAP7_75t_L g3781 ( 
.A(n_3395),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_L g3782 ( 
.A(n_3224),
.B(n_2604),
.Y(n_3782)
);

AOI21xp5_ASAP7_75t_L g3783 ( 
.A1(n_3302),
.A2(n_2757),
.B(n_2744),
.Y(n_3783)
);

OR2x2_ASAP7_75t_L g3784 ( 
.A(n_3428),
.B(n_2846),
.Y(n_3784)
);

OA21x2_ASAP7_75t_L g3785 ( 
.A1(n_3515),
.A2(n_2847),
.B(n_2920),
.Y(n_3785)
);

NOR4xp25_ASAP7_75t_L g3786 ( 
.A(n_3527),
.B(n_2754),
.C(n_2853),
.D(n_2852),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3269),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3312),
.B(n_479),
.Y(n_3788)
);

AOI21xp5_ASAP7_75t_SL g3789 ( 
.A1(n_3312),
.A2(n_2923),
.B(n_2921),
.Y(n_3789)
);

NOR2xp33_ASAP7_75t_L g3790 ( 
.A(n_3610),
.B(n_2880),
.Y(n_3790)
);

AOI221xp5_ASAP7_75t_SL g3791 ( 
.A1(n_3400),
.A2(n_2911),
.B1(n_2898),
.B2(n_2834),
.C(n_2858),
.Y(n_3791)
);

OA21x2_ASAP7_75t_L g3792 ( 
.A1(n_3551),
.A2(n_2932),
.B(n_2929),
.Y(n_3792)
);

AOI22xp33_ASAP7_75t_L g3793 ( 
.A1(n_3523),
.A2(n_3135),
.B1(n_3143),
.B2(n_3118),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3323),
.B(n_2608),
.Y(n_3794)
);

INVx3_ASAP7_75t_SL g3795 ( 
.A(n_3362),
.Y(n_3795)
);

AOI21x1_ASAP7_75t_L g3796 ( 
.A1(n_3637),
.A2(n_2945),
.B(n_2935),
.Y(n_3796)
);

NAND3xp33_ASAP7_75t_L g3797 ( 
.A(n_3358),
.B(n_3169),
.C(n_3165),
.Y(n_3797)
);

AOI22xp5_ASAP7_75t_L g3798 ( 
.A1(n_3256),
.A2(n_2950),
.B1(n_2951),
.B2(n_2946),
.Y(n_3798)
);

OAI21x1_ASAP7_75t_L g3799 ( 
.A1(n_3734),
.A2(n_3117),
.B(n_3080),
.Y(n_3799)
);

AOI21xp5_ASAP7_75t_L g3800 ( 
.A1(n_3478),
.A2(n_3602),
.B(n_3497),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3428),
.B(n_2795),
.Y(n_3801)
);

AND2x2_ASAP7_75t_L g3802 ( 
.A(n_3518),
.B(n_3455),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3272),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_SL g3804 ( 
.A(n_3597),
.B(n_3164),
.Y(n_3804)
);

AOI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_3307),
.A2(n_3198),
.B(n_3193),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3350),
.Y(n_3806)
);

OAI21x1_ASAP7_75t_L g3807 ( 
.A1(n_3618),
.A2(n_3164),
.B(n_2852),
.Y(n_3807)
);

AO32x2_ASAP7_75t_L g3808 ( 
.A1(n_3468),
.A2(n_2966),
.A3(n_3009),
.B1(n_2961),
.B2(n_2955),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3373),
.Y(n_3809)
);

BUFx10_ASAP7_75t_L g3810 ( 
.A(n_3258),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3285),
.Y(n_3811)
);

AOI21xp5_ASAP7_75t_L g3812 ( 
.A1(n_3584),
.A2(n_3115),
.B(n_3113),
.Y(n_3812)
);

OAI21x1_ASAP7_75t_L g3813 ( 
.A1(n_3371),
.A2(n_2795),
.B(n_3012),
.Y(n_3813)
);

OAI21xp5_ASAP7_75t_L g3814 ( 
.A1(n_3374),
.A2(n_3535),
.B(n_3687),
.Y(n_3814)
);

BUFx10_ASAP7_75t_L g3815 ( 
.A(n_3496),
.Y(n_3815)
);

BUFx6f_ASAP7_75t_L g3816 ( 
.A(n_3568),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3297),
.Y(n_3817)
);

OAI21x1_ASAP7_75t_L g3818 ( 
.A1(n_3514),
.A2(n_3018),
.B(n_3014),
.Y(n_3818)
);

INVxp67_ASAP7_75t_SL g3819 ( 
.A(n_3603),
.Y(n_3819)
);

A2O1A1Ixp33_ASAP7_75t_L g3820 ( 
.A1(n_3225),
.A2(n_3025),
.B(n_3030),
.C(n_3021),
.Y(n_3820)
);

AOI21xp5_ASAP7_75t_L g3821 ( 
.A1(n_3639),
.A2(n_3191),
.B(n_3044),
.Y(n_3821)
);

INVx2_ASAP7_75t_L g3822 ( 
.A(n_3404),
.Y(n_3822)
);

AOI22xp5_ASAP7_75t_L g3823 ( 
.A1(n_3702),
.A2(n_3053),
.B1(n_3055),
.B2(n_3035),
.Y(n_3823)
);

O2A1O1Ixp33_ASAP7_75t_L g3824 ( 
.A1(n_3615),
.A2(n_3074),
.B(n_3076),
.C(n_3063),
.Y(n_3824)
);

OAI21x1_ASAP7_75t_L g3825 ( 
.A1(n_3589),
.A2(n_3083),
.B(n_3078),
.Y(n_3825)
);

NOR2xp33_ASAP7_75t_L g3826 ( 
.A(n_3465),
.B(n_2719),
.Y(n_3826)
);

INVx3_ASAP7_75t_L g3827 ( 
.A(n_3445),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3696),
.A2(n_3154),
.B(n_3148),
.Y(n_3828)
);

BUFx3_ASAP7_75t_L g3829 ( 
.A(n_3683),
.Y(n_3829)
);

AOI21xp5_ASAP7_75t_L g3830 ( 
.A1(n_3711),
.A2(n_3724),
.B(n_3651),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3301),
.Y(n_3831)
);

OAI21x1_ASAP7_75t_L g3832 ( 
.A1(n_3605),
.A2(n_3092),
.B(n_3085),
.Y(n_3832)
);

OAI21x1_ASAP7_75t_L g3833 ( 
.A1(n_3229),
.A2(n_3099),
.B(n_3095),
.Y(n_3833)
);

A2O1A1Ixp33_ASAP7_75t_L g3834 ( 
.A1(n_3359),
.A2(n_3626),
.B(n_3390),
.C(n_3473),
.Y(n_3834)
);

OR2x6_ASAP7_75t_L g3835 ( 
.A(n_3445),
.B(n_3100),
.Y(n_3835)
);

AOI21xp33_ASAP7_75t_L g3836 ( 
.A1(n_3492),
.A2(n_2743),
.B(n_2889),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3630),
.B(n_3106),
.Y(n_3837)
);

AOI22xp33_ASAP7_75t_L g3838 ( 
.A1(n_3559),
.A2(n_3111),
.B1(n_3158),
.B2(n_3116),
.Y(n_3838)
);

O2A1O1Ixp33_ASAP7_75t_SL g3839 ( 
.A1(n_3324),
.A2(n_3176),
.B(n_3189),
.C(n_3184),
.Y(n_3839)
);

BUFx12f_ASAP7_75t_L g3840 ( 
.A(n_3299),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3235),
.B(n_2743),
.Y(n_3841)
);

AO31x2_ASAP7_75t_L g3842 ( 
.A1(n_3670),
.A2(n_3716),
.A3(n_3209),
.B(n_3665),
.Y(n_3842)
);

OR2x2_ASAP7_75t_L g3843 ( 
.A(n_3547),
.B(n_480),
.Y(n_3843)
);

BUFx2_ASAP7_75t_L g3844 ( 
.A(n_3617),
.Y(n_3844)
);

INVx4_ASAP7_75t_L g3845 ( 
.A(n_3217),
.Y(n_3845)
);

NAND3x1_ASAP7_75t_L g3846 ( 
.A(n_3311),
.B(n_481),
.C(n_482),
.Y(n_3846)
);

OAI22xp5_ASAP7_75t_L g3847 ( 
.A1(n_3559),
.A2(n_2889),
.B1(n_483),
.B2(n_481),
.Y(n_3847)
);

O2A1O1Ixp33_ASAP7_75t_SL g3848 ( 
.A1(n_3469),
.A2(n_483),
.B(n_481),
.C(n_482),
.Y(n_3848)
);

OAI221xp5_ASAP7_75t_L g3849 ( 
.A1(n_3674),
.A2(n_2889),
.B1(n_485),
.B2(n_482),
.C(n_484),
.Y(n_3849)
);

AOI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_3380),
.A2(n_484),
.B(n_485),
.Y(n_3850)
);

BUFx6f_ASAP7_75t_L g3851 ( 
.A(n_3494),
.Y(n_3851)
);

A2O1A1Ixp33_ASAP7_75t_L g3852 ( 
.A1(n_3662),
.A2(n_486),
.B(n_484),
.C(n_485),
.Y(n_3852)
);

AO31x2_ASAP7_75t_L g3853 ( 
.A1(n_3463),
.A2(n_488),
.A3(n_486),
.B(n_487),
.Y(n_3853)
);

NAND2x1_ASAP7_75t_L g3854 ( 
.A(n_3623),
.B(n_487),
.Y(n_3854)
);

OAI21x1_ASAP7_75t_L g3855 ( 
.A1(n_3369),
.A2(n_489),
.B(n_488),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3682),
.B(n_487),
.Y(n_3856)
);

OAI22xp33_ASAP7_75t_L g3857 ( 
.A1(n_3518),
.A2(n_490),
.B1(n_488),
.B2(n_489),
.Y(n_3857)
);

AO32x2_ASAP7_75t_L g3858 ( 
.A1(n_3452),
.A2(n_491),
.A3(n_489),
.B1(n_490),
.B2(n_492),
.Y(n_3858)
);

OAI21x1_ASAP7_75t_L g3859 ( 
.A1(n_3729),
.A2(n_495),
.B(n_494),
.Y(n_3859)
);

A2O1A1Ixp33_ASAP7_75t_L g3860 ( 
.A1(n_3677),
.A2(n_495),
.B(n_493),
.C(n_494),
.Y(n_3860)
);

AO32x2_ASAP7_75t_L g3861 ( 
.A1(n_3723),
.A2(n_495),
.A3(n_493),
.B1(n_494),
.B2(n_496),
.Y(n_3861)
);

AO31x2_ASAP7_75t_L g3862 ( 
.A1(n_3480),
.A2(n_497),
.A3(n_493),
.B(n_496),
.Y(n_3862)
);

OAI21x1_ASAP7_75t_L g3863 ( 
.A1(n_3641),
.A2(n_498),
.B(n_497),
.Y(n_3863)
);

OA21x2_ASAP7_75t_L g3864 ( 
.A1(n_3516),
.A2(n_496),
.B(n_497),
.Y(n_3864)
);

INVx1_ASAP7_75t_SL g3865 ( 
.A(n_3383),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3199),
.B(n_498),
.Y(n_3866)
);

NOR2xp33_ASAP7_75t_SL g3867 ( 
.A(n_3493),
.B(n_498),
.Y(n_3867)
);

INVxp67_ASAP7_75t_SL g3868 ( 
.A(n_3334),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3202),
.B(n_499),
.Y(n_3869)
);

AOI21xp33_ASAP7_75t_L g3870 ( 
.A1(n_3731),
.A2(n_499),
.B(n_500),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_3387),
.A2(n_3425),
.B(n_3411),
.Y(n_3871)
);

OAI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3402),
.A2(n_499),
.B(n_501),
.Y(n_3872)
);

NOR2xp33_ASAP7_75t_L g3873 ( 
.A(n_3465),
.B(n_3544),
.Y(n_3873)
);

AOI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3429),
.A2(n_501),
.B(n_502),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_SL g3875 ( 
.A(n_3601),
.B(n_502),
.Y(n_3875)
);

AOI221xp5_ASAP7_75t_L g3876 ( 
.A1(n_3308),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.C(n_505),
.Y(n_3876)
);

AOI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_3466),
.A2(n_3487),
.B(n_3486),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3388),
.B(n_503),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_SL g3879 ( 
.A1(n_3547),
.A2(n_503),
.B(n_504),
.Y(n_3879)
);

INVx2_ASAP7_75t_SL g3880 ( 
.A(n_3251),
.Y(n_3880)
);

OAI21x1_ASAP7_75t_L g3881 ( 
.A1(n_3203),
.A2(n_3200),
.B(n_3276),
.Y(n_3881)
);

NOR2xp67_ASAP7_75t_L g3882 ( 
.A(n_3524),
.B(n_3273),
.Y(n_3882)
);

OAI22xp5_ASAP7_75t_L g3883 ( 
.A1(n_3555),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3490),
.A2(n_505),
.B(n_506),
.Y(n_3884)
);

OAI21x1_ASAP7_75t_SL g3885 ( 
.A1(n_3327),
.A2(n_507),
.B(n_508),
.Y(n_3885)
);

AO31x2_ASAP7_75t_L g3886 ( 
.A1(n_3582),
.A2(n_510),
.A3(n_507),
.B(n_509),
.Y(n_3886)
);

CKINVDCx11_ASAP7_75t_R g3887 ( 
.A(n_3353),
.Y(n_3887)
);

AOI21xp5_ASAP7_75t_L g3888 ( 
.A1(n_3495),
.A2(n_510),
.B(n_511),
.Y(n_3888)
);

BUFx3_ASAP7_75t_L g3889 ( 
.A(n_3354),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3326),
.Y(n_3890)
);

AOI21xp33_ASAP7_75t_SL g3891 ( 
.A1(n_3379),
.A2(n_510),
.B(n_511),
.Y(n_3891)
);

BUFx6f_ASAP7_75t_L g3892 ( 
.A(n_3376),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3208),
.B(n_3212),
.Y(n_3893)
);

OAI21x1_ASAP7_75t_L g3894 ( 
.A1(n_3375),
.A2(n_513),
.B(n_512),
.Y(n_3894)
);

AND2x4_ASAP7_75t_L g3895 ( 
.A(n_3360),
.B(n_511),
.Y(n_3895)
);

O2A1O1Ixp33_ASAP7_75t_SL g3896 ( 
.A1(n_3593),
.A2(n_514),
.B(n_512),
.C(n_513),
.Y(n_3896)
);

BUFx2_ASAP7_75t_L g3897 ( 
.A(n_3217),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3216),
.B(n_512),
.Y(n_3898)
);

AO31x2_ASAP7_75t_L g3899 ( 
.A1(n_3426),
.A2(n_3650),
.A3(n_3261),
.B(n_3405),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3328),
.Y(n_3900)
);

CKINVDCx5p33_ASAP7_75t_R g3901 ( 
.A(n_3366),
.Y(n_3901)
);

CKINVDCx14_ASAP7_75t_R g3902 ( 
.A(n_3227),
.Y(n_3902)
);

OAI21x1_ASAP7_75t_L g3903 ( 
.A1(n_3232),
.A2(n_516),
.B(n_515),
.Y(n_3903)
);

INVx2_ASAP7_75t_SL g3904 ( 
.A(n_3340),
.Y(n_3904)
);

A2O1A1Ixp33_ASAP7_75t_L g3905 ( 
.A1(n_3714),
.A2(n_516),
.B(n_513),
.C(n_515),
.Y(n_3905)
);

OAI21x1_ASAP7_75t_L g3906 ( 
.A1(n_3609),
.A2(n_517),
.B(n_516),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3500),
.A2(n_515),
.B(n_517),
.Y(n_3907)
);

AOI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_3507),
.A2(n_517),
.B(n_518),
.Y(n_3908)
);

INVx3_ASAP7_75t_L g3909 ( 
.A(n_3368),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_3233),
.B(n_518),
.Y(n_3910)
);

OAI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3555),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.Y(n_3911)
);

CKINVDCx5p33_ASAP7_75t_R g3912 ( 
.A(n_3446),
.Y(n_3912)
);

A2O1A1Ixp33_ASAP7_75t_L g3913 ( 
.A1(n_3726),
.A2(n_521),
.B(n_519),
.C(n_520),
.Y(n_3913)
);

NAND2x1p5_ASAP7_75t_L g3914 ( 
.A(n_3443),
.B(n_3580),
.Y(n_3914)
);

OAI21xp5_ASAP7_75t_L g3915 ( 
.A1(n_3238),
.A2(n_519),
.B(n_520),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3336),
.Y(n_3916)
);

O2A1O1Ixp33_ASAP7_75t_L g3917 ( 
.A1(n_3343),
.A2(n_523),
.B(n_521),
.C(n_522),
.Y(n_3917)
);

INVx2_ASAP7_75t_L g3918 ( 
.A(n_3421),
.Y(n_3918)
);

AOI21x1_ASAP7_75t_L g3919 ( 
.A1(n_3588),
.A2(n_701),
.B(n_700),
.Y(n_3919)
);

AOI22xp5_ASAP7_75t_L g3920 ( 
.A1(n_3270),
.A2(n_524),
.B1(n_522),
.B2(n_523),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3244),
.B(n_524),
.Y(n_3921)
);

AOI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_3519),
.A2(n_524),
.B(n_525),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3246),
.B(n_3247),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3432),
.Y(n_3924)
);

AOI21xp5_ASAP7_75t_L g3925 ( 
.A1(n_3538),
.A2(n_525),
.B(n_526),
.Y(n_3925)
);

INVx5_ASAP7_75t_L g3926 ( 
.A(n_3223),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3345),
.Y(n_3927)
);

OAI22x1_ASAP7_75t_L g3928 ( 
.A1(n_3564),
.A2(n_527),
.B1(n_525),
.B2(n_526),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3451),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3253),
.B(n_527),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_3566),
.A2(n_528),
.B(n_529),
.Y(n_3931)
);

AOI22xp33_ASAP7_75t_L g3932 ( 
.A1(n_3671),
.A2(n_530),
.B1(n_528),
.B2(n_529),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3590),
.B(n_529),
.Y(n_3933)
);

AND2x4_ASAP7_75t_L g3934 ( 
.A(n_3223),
.B(n_531),
.Y(n_3934)
);

OAI21xp5_ASAP7_75t_L g3935 ( 
.A1(n_3709),
.A2(n_531),
.B(n_532),
.Y(n_3935)
);

AO31x2_ASAP7_75t_L g3936 ( 
.A1(n_3623),
.A2(n_533),
.A3(n_531),
.B(n_532),
.Y(n_3936)
);

O2A1O1Ixp33_ASAP7_75t_L g3937 ( 
.A1(n_3317),
.A2(n_3364),
.B(n_3397),
.C(n_3676),
.Y(n_3937)
);

AO31x2_ASAP7_75t_L g3938 ( 
.A1(n_3377),
.A2(n_535),
.A3(n_533),
.B(n_534),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3472),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3567),
.B(n_533),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3477),
.Y(n_3941)
);

AOI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_3587),
.A2(n_534),
.B(n_535),
.Y(n_3942)
);

BUFx12f_ASAP7_75t_L g3943 ( 
.A(n_3489),
.Y(n_3943)
);

AO31x2_ASAP7_75t_L g3944 ( 
.A1(n_3409),
.A2(n_538),
.A3(n_536),
.B(n_537),
.Y(n_3944)
);

O2A1O1Ixp33_ASAP7_75t_L g3945 ( 
.A1(n_3386),
.A2(n_3367),
.B(n_3384),
.C(n_3355),
.Y(n_3945)
);

BUFx2_ASAP7_75t_L g3946 ( 
.A(n_3539),
.Y(n_3946)
);

BUFx3_ASAP7_75t_L g3947 ( 
.A(n_3423),
.Y(n_3947)
);

BUFx4f_ASAP7_75t_L g3948 ( 
.A(n_3489),
.Y(n_3948)
);

A2O1A1Ixp33_ASAP7_75t_L g3949 ( 
.A1(n_3329),
.A2(n_540),
.B(n_537),
.C(n_539),
.Y(n_3949)
);

AOI21xp5_ASAP7_75t_SL g3950 ( 
.A1(n_3215),
.A2(n_537),
.B(n_539),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3361),
.Y(n_3951)
);

OAI21x1_ASAP7_75t_L g3952 ( 
.A1(n_3616),
.A2(n_3703),
.B(n_3278),
.Y(n_3952)
);

AO21x2_ASAP7_75t_L g3953 ( 
.A1(n_3453),
.A2(n_539),
.B(n_541),
.Y(n_3953)
);

AND2x2_ASAP7_75t_L g3954 ( 
.A(n_3215),
.B(n_3234),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3365),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3599),
.B(n_3600),
.Y(n_3956)
);

CKINVDCx20_ASAP7_75t_R g3957 ( 
.A(n_3318),
.Y(n_3957)
);

OAI21x1_ASAP7_75t_L g3958 ( 
.A1(n_3444),
.A2(n_543),
.B(n_542),
.Y(n_3958)
);

OAI21x1_ASAP7_75t_L g3959 ( 
.A1(n_3408),
.A2(n_543),
.B(n_542),
.Y(n_3959)
);

OAI21x1_ASAP7_75t_L g3960 ( 
.A1(n_3449),
.A2(n_544),
.B(n_542),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3608),
.B(n_541),
.Y(n_3961)
);

AOI21xp5_ASAP7_75t_L g3962 ( 
.A1(n_3631),
.A2(n_3679),
.B(n_3672),
.Y(n_3962)
);

AOI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3689),
.A2(n_541),
.B(n_544),
.Y(n_3963)
);

OAI21x1_ASAP7_75t_L g3964 ( 
.A1(n_3510),
.A2(n_546),
.B(n_545),
.Y(n_3964)
);

INVx4_ASAP7_75t_L g3965 ( 
.A(n_3399),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3263),
.B(n_544),
.Y(n_3966)
);

AOI31xp67_ASAP7_75t_L g3967 ( 
.A1(n_3513),
.A2(n_547),
.A3(n_545),
.B(n_546),
.Y(n_3967)
);

OAI21x1_ASAP7_75t_L g3968 ( 
.A1(n_3565),
.A2(n_548),
.B(n_547),
.Y(n_3968)
);

AOI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3692),
.A2(n_546),
.B(n_547),
.Y(n_3969)
);

OAI21x1_ASAP7_75t_L g3970 ( 
.A1(n_3274),
.A2(n_550),
.B(n_549),
.Y(n_3970)
);

AOI21xp5_ASAP7_75t_L g3971 ( 
.A1(n_3720),
.A2(n_548),
.B(n_549),
.Y(n_3971)
);

AOI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_3464),
.A2(n_549),
.B(n_550),
.Y(n_3972)
);

NOR2xp33_ASAP7_75t_L g3973 ( 
.A(n_3520),
.B(n_551),
.Y(n_3973)
);

AOI21xp33_ASAP7_75t_L g3974 ( 
.A1(n_3476),
.A2(n_552),
.B(n_553),
.Y(n_3974)
);

OAI22xp5_ASAP7_75t_L g3975 ( 
.A1(n_3234),
.A2(n_3245),
.B1(n_3287),
.B2(n_3457),
.Y(n_3975)
);

NOR2xp67_ASAP7_75t_L g3976 ( 
.A(n_3622),
.B(n_552),
.Y(n_3976)
);

AOI22xp5_ASAP7_75t_L g3977 ( 
.A1(n_3319),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3264),
.B(n_553),
.Y(n_3978)
);

NOR2xp33_ASAP7_75t_L g3979 ( 
.A(n_3572),
.B(n_3458),
.Y(n_3979)
);

BUFx8_ASAP7_75t_L g3980 ( 
.A(n_3320),
.Y(n_3980)
);

INVx2_ASAP7_75t_L g3981 ( 
.A(n_3498),
.Y(n_3981)
);

AOI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3479),
.A2(n_554),
.B(n_556),
.Y(n_3982)
);

AND2x4_ASAP7_75t_L g3983 ( 
.A(n_3506),
.B(n_3571),
.Y(n_3983)
);

OAI21x1_ASAP7_75t_L g3984 ( 
.A1(n_3275),
.A2(n_558),
.B(n_557),
.Y(n_3984)
);

AOI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3481),
.A2(n_556),
.B(n_557),
.Y(n_3985)
);

AO22x2_ASAP7_75t_L g3986 ( 
.A1(n_3417),
.A2(n_559),
.B1(n_556),
.B2(n_558),
.Y(n_3986)
);

AOI21xp5_ASAP7_75t_L g3987 ( 
.A1(n_3484),
.A2(n_559),
.B(n_560),
.Y(n_3987)
);

OAI21x1_ASAP7_75t_L g3988 ( 
.A1(n_3688),
.A2(n_3717),
.B(n_3288),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_3505),
.Y(n_3989)
);

A2O1A1Ixp33_ASAP7_75t_L g3990 ( 
.A1(n_3204),
.A2(n_561),
.B(n_559),
.C(n_560),
.Y(n_3990)
);

OAI21x1_ASAP7_75t_L g3991 ( 
.A1(n_3283),
.A2(n_562),
.B(n_561),
.Y(n_3991)
);

AOI21x1_ASAP7_75t_L g3992 ( 
.A1(n_3625),
.A2(n_702),
.B(n_701),
.Y(n_3992)
);

OAI21xp5_ASAP7_75t_SL g3993 ( 
.A1(n_3314),
.A2(n_569),
.B(n_560),
.Y(n_3993)
);

AO22x2_ASAP7_75t_L g3994 ( 
.A1(n_3316),
.A2(n_563),
.B1(n_561),
.B2(n_562),
.Y(n_3994)
);

OAI21xp5_ASAP7_75t_L g3995 ( 
.A1(n_3577),
.A2(n_3579),
.B(n_3583),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3339),
.B(n_562),
.Y(n_3996)
);

AOI221x1_ASAP7_75t_L g3997 ( 
.A1(n_3330),
.A2(n_566),
.B1(n_564),
.B2(n_565),
.C(n_568),
.Y(n_3997)
);

BUFx3_ASAP7_75t_L g3998 ( 
.A(n_3592),
.Y(n_3998)
);

AOI221x1_ASAP7_75t_L g3999 ( 
.A1(n_3673),
.A2(n_568),
.B1(n_564),
.B2(n_565),
.C(n_569),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3512),
.Y(n_4000)
);

AO31x2_ASAP7_75t_L g4001 ( 
.A1(n_3403),
.A2(n_571),
.A3(n_569),
.B(n_570),
.Y(n_4001)
);

OAI22xp5_ASAP7_75t_L g4002 ( 
.A1(n_3245),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_4002)
);

NAND2x1p5_ASAP7_75t_L g4003 ( 
.A(n_3320),
.B(n_571),
.Y(n_4003)
);

AOI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3499),
.A2(n_572),
.B(n_573),
.Y(n_4004)
);

AOI21xp5_ASAP7_75t_L g4005 ( 
.A1(n_3501),
.A2(n_573),
.B(n_574),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3502),
.A2(n_573),
.B(n_574),
.Y(n_4006)
);

AOI21x1_ASAP7_75t_L g4007 ( 
.A1(n_3704),
.A2(n_704),
.B(n_702),
.Y(n_4007)
);

OAI22x1_ASAP7_75t_L g4008 ( 
.A1(n_3406),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_4008)
);

AOI221xp5_ASAP7_75t_SL g4009 ( 
.A1(n_3474),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.C(n_578),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3549),
.Y(n_4010)
);

INVx2_ASAP7_75t_SL g4011 ( 
.A(n_3522),
.Y(n_4011)
);

NOR2xp67_ASAP7_75t_L g4012 ( 
.A(n_3666),
.B(n_575),
.Y(n_4012)
);

AND2x2_ASAP7_75t_L g4013 ( 
.A(n_3613),
.B(n_576),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3619),
.B(n_578),
.Y(n_4014)
);

AOI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_3511),
.A2(n_579),
.B(n_580),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3517),
.A2(n_579),
.B(n_580),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3239),
.Y(n_4017)
);

A2O1A1Ixp33_ASAP7_75t_L g4018 ( 
.A1(n_3450),
.A2(n_582),
.B(n_580),
.C(n_581),
.Y(n_4018)
);

OR2x2_ASAP7_75t_L g4019 ( 
.A(n_3221),
.B(n_3528),
.Y(n_4019)
);

AOI21xp5_ASAP7_75t_L g4020 ( 
.A1(n_3525),
.A2(n_581),
.B(n_582),
.Y(n_4020)
);

AOI221x1_ASAP7_75t_L g4021 ( 
.A1(n_3548),
.A2(n_584),
.B1(n_581),
.B2(n_583),
.C(n_585),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3287),
.Y(n_4022)
);

OAI21x1_ASAP7_75t_L g4023 ( 
.A1(n_3391),
.A2(n_583),
.B(n_584),
.Y(n_4023)
);

AOI21xp5_ASAP7_75t_L g4024 ( 
.A1(n_3532),
.A2(n_583),
.B(n_584),
.Y(n_4024)
);

O2A1O1Ixp5_ASAP7_75t_L g4025 ( 
.A1(n_3325),
.A2(n_587),
.B(n_585),
.C(n_586),
.Y(n_4025)
);

OAI21x1_ASAP7_75t_L g4026 ( 
.A1(n_3521),
.A2(n_585),
.B(n_586),
.Y(n_4026)
);

AO21x2_ASAP7_75t_L g4027 ( 
.A1(n_3540),
.A2(n_586),
.B(n_587),
.Y(n_4027)
);

AO21x1_ASAP7_75t_L g4028 ( 
.A1(n_3392),
.A2(n_588),
.B(n_589),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3218),
.Y(n_4029)
);

AOI221xp5_ASAP7_75t_L g4030 ( 
.A1(n_3412),
.A2(n_590),
.B1(n_588),
.B2(n_589),
.C(n_591),
.Y(n_4030)
);

INVx2_ASAP7_75t_L g4031 ( 
.A(n_3228),
.Y(n_4031)
);

OR2x2_ASAP7_75t_L g4032 ( 
.A(n_3237),
.B(n_590),
.Y(n_4032)
);

INVx2_ASAP7_75t_L g4033 ( 
.A(n_3554),
.Y(n_4033)
);

OAI21xp5_ASAP7_75t_L g4034 ( 
.A1(n_3250),
.A2(n_591),
.B(n_592),
.Y(n_4034)
);

A2O1A1Ixp33_ASAP7_75t_L g4035 ( 
.A1(n_3667),
.A2(n_3356),
.B(n_3349),
.C(n_3655),
.Y(n_4035)
);

OAI21xp5_ASAP7_75t_L g4036 ( 
.A1(n_3243),
.A2(n_3669),
.B(n_3659),
.Y(n_4036)
);

INVx6_ASAP7_75t_L g4037 ( 
.A(n_3399),
.Y(n_4037)
);

AO21x2_ASAP7_75t_L g4038 ( 
.A1(n_3542),
.A2(n_591),
.B(n_592),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_SL g4039 ( 
.A(n_3556),
.B(n_593),
.Y(n_4039)
);

AND2x4_ASAP7_75t_L g4040 ( 
.A(n_3406),
.B(n_593),
.Y(n_4040)
);

AOI221xp5_ASAP7_75t_SL g4041 ( 
.A1(n_3611),
.A2(n_595),
.B1(n_593),
.B2(n_594),
.C(n_596),
.Y(n_4041)
);

OAI21x1_ASAP7_75t_L g4042 ( 
.A1(n_3596),
.A2(n_594),
.B(n_595),
.Y(n_4042)
);

NAND3x1_ASAP7_75t_L g4043 ( 
.A(n_3550),
.B(n_594),
.C(n_595),
.Y(n_4043)
);

OAI21x1_ASAP7_75t_L g4044 ( 
.A1(n_3694),
.A2(n_596),
.B(n_597),
.Y(n_4044)
);

OAI21x1_ASAP7_75t_L g4045 ( 
.A1(n_3695),
.A2(n_598),
.B(n_599),
.Y(n_4045)
);

NAND2xp33_ASAP7_75t_SL g4046 ( 
.A(n_3543),
.B(n_598),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3201),
.Y(n_4047)
);

AOI21xp5_ASAP7_75t_L g4048 ( 
.A1(n_3537),
.A2(n_599),
.B(n_600),
.Y(n_4048)
);

NAND2x1p5_ASAP7_75t_L g4049 ( 
.A(n_3556),
.B(n_599),
.Y(n_4049)
);

NOR2xp67_ASAP7_75t_L g4050 ( 
.A(n_3219),
.B(n_600),
.Y(n_4050)
);

OAI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_3291),
.A2(n_600),
.B(n_601),
.Y(n_4051)
);

INVx3_ASAP7_75t_SL g4052 ( 
.A(n_3241),
.Y(n_4052)
);

O2A1O1Ixp33_ASAP7_75t_L g4053 ( 
.A1(n_3454),
.A2(n_3331),
.B(n_3656),
.C(n_3335),
.Y(n_4053)
);

OAI21x1_ASAP7_75t_L g4054 ( 
.A1(n_3713),
.A2(n_601),
.B(n_602),
.Y(n_4054)
);

AOI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_3545),
.A2(n_602),
.B(n_603),
.Y(n_4055)
);

CKINVDCx5p33_ASAP7_75t_R g4056 ( 
.A(n_3385),
.Y(n_4056)
);

AOI21xp5_ASAP7_75t_L g4057 ( 
.A1(n_3553),
.A2(n_603),
.B(n_604),
.Y(n_4057)
);

AOI21xp5_ASAP7_75t_L g4058 ( 
.A1(n_3563),
.A2(n_603),
.B(n_604),
.Y(n_4058)
);

AND2x4_ASAP7_75t_L g4059 ( 
.A(n_3357),
.B(n_604),
.Y(n_4059)
);

OAI21xp5_ASAP7_75t_L g4060 ( 
.A1(n_3681),
.A2(n_605),
.B(n_606),
.Y(n_4060)
);

AOI21xp5_ASAP7_75t_L g4061 ( 
.A1(n_3569),
.A2(n_605),
.B(n_606),
.Y(n_4061)
);

AO31x2_ASAP7_75t_L g4062 ( 
.A1(n_3706),
.A2(n_608),
.A3(n_605),
.B(n_607),
.Y(n_4062)
);

CKINVDCx5p33_ASAP7_75t_R g4063 ( 
.A(n_3281),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3240),
.Y(n_4064)
);

BUFx3_ASAP7_75t_L g4065 ( 
.A(n_3249),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_4013),
.B(n_3351),
.Y(n_4066)
);

INVx4_ASAP7_75t_L g4067 ( 
.A(n_3760),
.Y(n_4067)
);

BUFx3_ASAP7_75t_L g4068 ( 
.A(n_3851),
.Y(n_4068)
);

AOI22xp5_ASAP7_75t_SL g4069 ( 
.A1(n_3750),
.A2(n_3415),
.B1(n_3570),
.B2(n_3574),
.Y(n_4069)
);

BUFx6f_ASAP7_75t_L g4070 ( 
.A(n_3851),
.Y(n_4070)
);

OAI21xp5_ASAP7_75t_L g4071 ( 
.A1(n_3830),
.A2(n_3210),
.B(n_3661),
.Y(n_4071)
);

INVx6_ASAP7_75t_L g4072 ( 
.A(n_3840),
.Y(n_4072)
);

OAI22xp5_ASAP7_75t_L g4073 ( 
.A1(n_3948),
.A2(n_3257),
.B1(n_3293),
.B2(n_3279),
.Y(n_4073)
);

INVx4_ASAP7_75t_L g4074 ( 
.A(n_3795),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3761),
.Y(n_4075)
);

NAND2x1p5_ASAP7_75t_L g4076 ( 
.A(n_3926),
.B(n_3574),
.Y(n_4076)
);

INVx2_ASAP7_75t_SL g4077 ( 
.A(n_4063),
.Y(n_4077)
);

OAI22xp5_ASAP7_75t_SL g4078 ( 
.A1(n_3943),
.A2(n_3442),
.B1(n_3424),
.B2(n_3483),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_4046),
.A2(n_3643),
.B1(n_3635),
.B2(n_3685),
.Y(n_4079)
);

INVx6_ASAP7_75t_L g4080 ( 
.A(n_3980),
.Y(n_4080)
);

BUFx4f_ASAP7_75t_SL g4081 ( 
.A(n_3747),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3736),
.B(n_3430),
.Y(n_4082)
);

AOI22xp5_ASAP7_75t_L g4083 ( 
.A1(n_3975),
.A2(n_3485),
.B1(n_3462),
.B2(n_3558),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3787),
.Y(n_4084)
);

BUFx12f_ASAP7_75t_L g4085 ( 
.A(n_3887),
.Y(n_4085)
);

AOI22xp33_ASAP7_75t_L g4086 ( 
.A1(n_3765),
.A2(n_3644),
.B1(n_3647),
.B2(n_3645),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3803),
.Y(n_4087)
);

INVx8_ASAP7_75t_L g4088 ( 
.A(n_3926),
.Y(n_4088)
);

HB1xp67_ASAP7_75t_L g4089 ( 
.A(n_3819),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3811),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_3742),
.Y(n_4091)
);

AOI22xp33_ASAP7_75t_L g4092 ( 
.A1(n_3758),
.A2(n_3647),
.B1(n_3645),
.B2(n_3727),
.Y(n_4092)
);

BUFx3_ASAP7_75t_L g4093 ( 
.A(n_3781),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3788),
.B(n_3954),
.Y(n_4094)
);

AOI22xp33_ASAP7_75t_SL g4095 ( 
.A1(n_4037),
.A2(n_3430),
.B1(n_3286),
.B2(n_3280),
.Y(n_4095)
);

OAI22xp33_ASAP7_75t_L g4096 ( 
.A1(n_3993),
.A2(n_3401),
.B1(n_3213),
.B2(n_3347),
.Y(n_4096)
);

AOI22xp33_ASAP7_75t_L g4097 ( 
.A1(n_3847),
.A2(n_3727),
.B1(n_3684),
.B2(n_3471),
.Y(n_4097)
);

AOI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3934),
.A2(n_3348),
.B1(n_3621),
.B2(n_3730),
.Y(n_4098)
);

AOI22xp33_ASAP7_75t_L g4099 ( 
.A1(n_4036),
.A2(n_3560),
.B1(n_3561),
.B2(n_3536),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3800),
.B(n_3956),
.Y(n_4100)
);

OAI22xp33_ASAP7_75t_L g4101 ( 
.A1(n_3845),
.A2(n_4052),
.B1(n_4003),
.B2(n_3843),
.Y(n_4101)
);

CKINVDCx11_ASAP7_75t_R g4102 ( 
.A(n_3737),
.Y(n_4102)
);

INVx2_ASAP7_75t_L g4103 ( 
.A(n_3759),
.Y(n_4103)
);

AOI22xp33_ASAP7_75t_L g4104 ( 
.A1(n_3790),
.A2(n_3581),
.B1(n_3640),
.B2(n_3459),
.Y(n_4104)
);

OAI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_4049),
.A2(n_3541),
.B1(n_3378),
.B2(n_3562),
.Y(n_4105)
);

AOI22xp33_ASAP7_75t_SL g4106 ( 
.A1(n_4037),
.A2(n_3266),
.B1(n_3707),
.B2(n_3693),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_3767),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_L g4108 ( 
.A1(n_3986),
.A2(n_3267),
.B1(n_3718),
.B2(n_3575),
.Y(n_4108)
);

CKINVDCx20_ASAP7_75t_R g4109 ( 
.A(n_3957),
.Y(n_4109)
);

INVx2_ASAP7_75t_L g4110 ( 
.A(n_3768),
.Y(n_4110)
);

OAI22xp5_ASAP7_75t_L g4111 ( 
.A1(n_3897),
.A2(n_3398),
.B1(n_3546),
.B2(n_3509),
.Y(n_4111)
);

BUFx12f_ASAP7_75t_L g4112 ( 
.A(n_3815),
.Y(n_4112)
);

BUFx6f_ASAP7_75t_L g4113 ( 
.A(n_3781),
.Y(n_4113)
);

BUFx4f_ASAP7_75t_L g4114 ( 
.A(n_3892),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_3817),
.Y(n_4115)
);

AOI22xp33_ASAP7_75t_L g4116 ( 
.A1(n_3986),
.A2(n_3552),
.B1(n_3629),
.B2(n_3607),
.Y(n_4116)
);

INVx11_ASAP7_75t_L g4117 ( 
.A(n_3902),
.Y(n_4117)
);

OAI22xp5_ASAP7_75t_L g4118 ( 
.A1(n_3776),
.A2(n_3557),
.B1(n_3649),
.B2(n_3636),
.Y(n_4118)
);

OAI22xp33_ASAP7_75t_SL g4119 ( 
.A1(n_3867),
.A2(n_3341),
.B1(n_3338),
.B2(n_3298),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3770),
.Y(n_4120)
);

INVx2_ASAP7_75t_L g4121 ( 
.A(n_3806),
.Y(n_4121)
);

OAI22xp5_ASAP7_75t_L g4122 ( 
.A1(n_3965),
.A2(n_3668),
.B1(n_3585),
.B2(n_3370),
.Y(n_4122)
);

OAI22xp33_ASAP7_75t_SL g4123 ( 
.A1(n_3946),
.A2(n_3315),
.B1(n_3282),
.B2(n_3394),
.Y(n_4123)
);

BUFx4f_ASAP7_75t_SL g4124 ( 
.A(n_3745),
.Y(n_4124)
);

BUFx2_ASAP7_75t_L g4125 ( 
.A(n_3947),
.Y(n_4125)
);

BUFx12f_ASAP7_75t_L g4126 ( 
.A(n_3901),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3871),
.B(n_3342),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3809),
.Y(n_4128)
);

INVx6_ASAP7_75t_L g4129 ( 
.A(n_3816),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_3822),
.Y(n_4130)
);

CKINVDCx5p33_ASAP7_75t_R g4131 ( 
.A(n_3752),
.Y(n_4131)
);

OAI22xp5_ASAP7_75t_L g4132 ( 
.A1(n_3950),
.A2(n_3352),
.B1(n_3396),
.B2(n_3719),
.Y(n_4132)
);

HB1xp67_ASAP7_75t_L g4133 ( 
.A(n_3756),
.Y(n_4133)
);

AOI22xp33_ASAP7_75t_SL g4134 ( 
.A1(n_3802),
.A2(n_3410),
.B1(n_3372),
.B2(n_3678),
.Y(n_4134)
);

BUFx6f_ASAP7_75t_L g4135 ( 
.A(n_3816),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3831),
.Y(n_4136)
);

AOI22xp33_ASAP7_75t_L g4137 ( 
.A1(n_3849),
.A2(n_3675),
.B1(n_3657),
.B2(n_3382),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3890),
.Y(n_4138)
);

INVx1_ASAP7_75t_SL g4139 ( 
.A(n_3844),
.Y(n_4139)
);

INVxp67_ASAP7_75t_SL g4140 ( 
.A(n_3739),
.Y(n_4140)
);

AND2x2_ASAP7_75t_L g4141 ( 
.A(n_4040),
.B(n_3594),
.Y(n_4141)
);

AOI22xp33_ASAP7_75t_SL g4142 ( 
.A1(n_3995),
.A2(n_3431),
.B1(n_3441),
.B2(n_3735),
.Y(n_4142)
);

BUFx4f_ASAP7_75t_SL g4143 ( 
.A(n_3889),
.Y(n_4143)
);

OAI22xp5_ASAP7_75t_L g4144 ( 
.A1(n_4050),
.A2(n_3220),
.B1(n_3310),
.B2(n_3296),
.Y(n_4144)
);

AOI22xp33_ASAP7_75t_L g4145 ( 
.A1(n_3994),
.A2(n_3254),
.B1(n_3236),
.B2(n_3708),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3900),
.Y(n_4146)
);

INVx1_ASAP7_75t_SL g4147 ( 
.A(n_3829),
.Y(n_4147)
);

OAI22xp5_ASAP7_75t_L g4148 ( 
.A1(n_3846),
.A2(n_3690),
.B1(n_3686),
.B2(n_3578),
.Y(n_4148)
);

AOI22xp33_ASAP7_75t_L g4149 ( 
.A1(n_3994),
.A2(n_3333),
.B1(n_3491),
.B2(n_3488),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3916),
.Y(n_4150)
);

CKINVDCx6p67_ASAP7_75t_R g4151 ( 
.A(n_3892),
.Y(n_4151)
);

NAND2xp33_ASAP7_75t_SL g4152 ( 
.A(n_4008),
.B(n_3705),
.Y(n_4152)
);

BUFx2_ASAP7_75t_SL g4153 ( 
.A(n_3827),
.Y(n_4153)
);

INVx6_ASAP7_75t_L g4154 ( 
.A(n_3983),
.Y(n_4154)
);

INVx4_ASAP7_75t_L g4155 ( 
.A(n_3914),
.Y(n_4155)
);

INVx3_ASAP7_75t_L g4156 ( 
.A(n_3774),
.Y(n_4156)
);

AOI22xp33_ASAP7_75t_SL g4157 ( 
.A1(n_3878),
.A2(n_3700),
.B1(n_3248),
.B2(n_3260),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_3918),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3927),
.Y(n_4159)
);

INVx2_ASAP7_75t_SL g4160 ( 
.A(n_4065),
.Y(n_4160)
);

AOI22xp33_ASAP7_75t_L g4161 ( 
.A1(n_4030),
.A2(n_3606),
.B1(n_3627),
.B2(n_3413),
.Y(n_4161)
);

BUFx6f_ASAP7_75t_L g4162 ( 
.A(n_3998),
.Y(n_4162)
);

AOI22xp33_ASAP7_75t_L g4163 ( 
.A1(n_3935),
.A2(n_3416),
.B1(n_3419),
.B2(n_3418),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3951),
.Y(n_4164)
);

BUFx4_ASAP7_75t_R g4165 ( 
.A(n_3810),
.Y(n_4165)
);

AND2x4_ASAP7_75t_L g4166 ( 
.A(n_3865),
.B(n_3634),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3955),
.Y(n_4167)
);

OAI22xp5_ASAP7_75t_L g4168 ( 
.A1(n_3834),
.A2(n_3598),
.B1(n_3624),
.B2(n_3576),
.Y(n_4168)
);

HB1xp67_ASAP7_75t_L g4169 ( 
.A(n_4019),
.Y(n_4169)
);

OAI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_3784),
.A2(n_3252),
.B1(n_3699),
.B2(n_3698),
.Y(n_4170)
);

BUFx10_ASAP7_75t_L g4171 ( 
.A(n_4056),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3989),
.Y(n_4172)
);

INVx3_ASAP7_75t_L g4173 ( 
.A(n_3772),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4000),
.Y(n_4174)
);

INVx4_ASAP7_75t_SL g4175 ( 
.A(n_3895),
.Y(n_4175)
);

OAI22xp5_ASAP7_75t_L g4176 ( 
.A1(n_3879),
.A2(n_3290),
.B1(n_3728),
.B2(n_3721),
.Y(n_4176)
);

INVx6_ASAP7_75t_L g4177 ( 
.A(n_3801),
.Y(n_4177)
);

BUFx8_ASAP7_75t_L g4178 ( 
.A(n_4011),
.Y(n_4178)
);

AOI22xp5_ASAP7_75t_L g4179 ( 
.A1(n_3857),
.A2(n_3715),
.B1(n_3664),
.B2(n_3427),
.Y(n_4179)
);

AOI22xp33_ASAP7_75t_L g4180 ( 
.A1(n_3749),
.A2(n_3460),
.B1(n_3467),
.B2(n_3482),
.Y(n_4180)
);

AOI22xp33_ASAP7_75t_L g4181 ( 
.A1(n_3782),
.A2(n_3911),
.B1(n_3883),
.B2(n_3777),
.Y(n_4181)
);

AOI22xp33_ASAP7_75t_L g4182 ( 
.A1(n_3771),
.A2(n_3503),
.B1(n_3642),
.B2(n_3595),
.Y(n_4182)
);

AOI22xp33_ASAP7_75t_L g4183 ( 
.A1(n_3932),
.A2(n_3591),
.B1(n_3422),
.B2(n_3573),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3877),
.B(n_3697),
.Y(n_4184)
);

INVx11_ASAP7_75t_L g4185 ( 
.A(n_3912),
.Y(n_4185)
);

INVx2_ASAP7_75t_L g4186 ( 
.A(n_3924),
.Y(n_4186)
);

AOI22xp33_ASAP7_75t_L g4187 ( 
.A1(n_3794),
.A2(n_3433),
.B1(n_3658),
.B2(n_3654),
.Y(n_4187)
);

INVx6_ASAP7_75t_L g4188 ( 
.A(n_3835),
.Y(n_4188)
);

AOI22xp33_ASAP7_75t_L g4189 ( 
.A1(n_3966),
.A2(n_3504),
.B1(n_3322),
.B2(n_3313),
.Y(n_4189)
);

BUFx3_ASAP7_75t_L g4190 ( 
.A(n_3909),
.Y(n_4190)
);

OAI22xp5_ASAP7_75t_L g4191 ( 
.A1(n_3920),
.A2(n_3722),
.B1(n_3393),
.B2(n_3271),
.Y(n_4191)
);

OAI22xp5_ASAP7_75t_L g4192 ( 
.A1(n_3977),
.A2(n_3284),
.B1(n_3305),
.B2(n_3226),
.Y(n_4192)
);

BUFx3_ASAP7_75t_L g4193 ( 
.A(n_3880),
.Y(n_4193)
);

INVx5_ASAP7_75t_L g4194 ( 
.A(n_3835),
.Y(n_4194)
);

AOI22xp33_ASAP7_75t_L g4195 ( 
.A1(n_4028),
.A2(n_3363),
.B1(n_3646),
.B2(n_3294),
.Y(n_4195)
);

BUFx6f_ASAP7_75t_L g4196 ( 
.A(n_3904),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3962),
.B(n_3614),
.Y(n_4197)
);

INVx5_ASAP7_75t_L g4198 ( 
.A(n_4059),
.Y(n_4198)
);

AOI22xp5_ASAP7_75t_L g4199 ( 
.A1(n_4009),
.A2(n_3435),
.B1(n_3437),
.B2(n_3436),
.Y(n_4199)
);

AOI22xp33_ASAP7_75t_SL g4200 ( 
.A1(n_3885),
.A2(n_3733),
.B1(n_3295),
.B2(n_3381),
.Y(n_4200)
);

BUFx10_ASAP7_75t_L g4201 ( 
.A(n_3973),
.Y(n_4201)
);

INVx2_ASAP7_75t_L g4202 ( 
.A(n_3929),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4010),
.Y(n_4203)
);

INVx1_ASAP7_75t_SL g4204 ( 
.A(n_4032),
.Y(n_4204)
);

OAI21xp5_ASAP7_75t_SL g4205 ( 
.A1(n_3891),
.A2(n_4002),
.B(n_3997),
.Y(n_4205)
);

AOI22xp33_ASAP7_75t_L g4206 ( 
.A1(n_3838),
.A2(n_4039),
.B1(n_4022),
.B2(n_3876),
.Y(n_4206)
);

AOI22xp33_ASAP7_75t_L g4207 ( 
.A1(n_4034),
.A2(n_3304),
.B1(n_3691),
.B2(n_3440),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_3893),
.Y(n_4208)
);

INVx6_ASAP7_75t_L g4209 ( 
.A(n_3882),
.Y(n_4209)
);

AOI22xp33_ASAP7_75t_L g4210 ( 
.A1(n_3778),
.A2(n_3438),
.B1(n_3447),
.B2(n_3434),
.Y(n_4210)
);

AOI22xp33_ASAP7_75t_SL g4211 ( 
.A1(n_3873),
.A2(n_3295),
.B1(n_3381),
.B2(n_3332),
.Y(n_4211)
);

AOI22xp33_ASAP7_75t_L g4212 ( 
.A1(n_4047),
.A2(n_3638),
.B1(n_3648),
.B2(n_3620),
.Y(n_4212)
);

CKINVDCx12_ASAP7_75t_R g4213 ( 
.A(n_3939),
.Y(n_4213)
);

OAI22xp33_ASAP7_75t_L g4214 ( 
.A1(n_3976),
.A2(n_4012),
.B1(n_3856),
.B2(n_3928),
.Y(n_4214)
);

CKINVDCx20_ASAP7_75t_R g4215 ( 
.A(n_3875),
.Y(n_4215)
);

INVxp67_ASAP7_75t_SL g4216 ( 
.A(n_3804),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_3923),
.Y(n_4217)
);

OAI21xp33_ASAP7_75t_L g4218 ( 
.A1(n_3786),
.A2(n_3586),
.B(n_3255),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4017),
.Y(n_4219)
);

BUFx10_ASAP7_75t_L g4220 ( 
.A(n_3979),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3941),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_3981),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_4029),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4031),
.Y(n_4224)
);

AOI22xp33_ASAP7_75t_L g4225 ( 
.A1(n_4064),
.A2(n_3332),
.B1(n_3381),
.B2(n_3295),
.Y(n_4225)
);

INVx2_ASAP7_75t_L g4226 ( 
.A(n_4033),
.Y(n_4226)
);

BUFx2_ASAP7_75t_L g4227 ( 
.A(n_3868),
.Y(n_4227)
);

BUFx10_ASAP7_75t_L g4228 ( 
.A(n_3826),
.Y(n_4228)
);

AOI22xp33_ASAP7_75t_L g4229 ( 
.A1(n_4051),
.A2(n_3814),
.B1(n_3870),
.B2(n_3974),
.Y(n_4229)
);

CKINVDCx5p33_ASAP7_75t_R g4230 ( 
.A(n_3740),
.Y(n_4230)
);

BUFx6f_ASAP7_75t_L g4231 ( 
.A(n_3854),
.Y(n_4231)
);

BUFx2_ASAP7_75t_L g4232 ( 
.A(n_3799),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_4014),
.B(n_607),
.Y(n_4233)
);

CKINVDCx6p67_ASAP7_75t_R g4234 ( 
.A(n_3933),
.Y(n_4234)
);

BUFx4f_ASAP7_75t_SL g4235 ( 
.A(n_4043),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_3936),
.Y(n_4236)
);

AOI22xp33_ASAP7_75t_SL g4237 ( 
.A1(n_4060),
.A2(n_3389),
.B1(n_3475),
.B2(n_3332),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3936),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_3940),
.Y(n_4239)
);

INVx6_ASAP7_75t_L g4240 ( 
.A(n_3789),
.Y(n_4240)
);

CKINVDCx5p33_ASAP7_75t_R g4241 ( 
.A(n_3996),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_3961),
.Y(n_4242)
);

BUFx6f_ASAP7_75t_L g4243 ( 
.A(n_3906),
.Y(n_4243)
);

CKINVDCx5p33_ASAP7_75t_R g4244 ( 
.A(n_3866),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3869),
.Y(n_4245)
);

INVx3_ASAP7_75t_L g4246 ( 
.A(n_3992),
.Y(n_4246)
);

AOI22xp33_ASAP7_75t_L g4247 ( 
.A1(n_3823),
.A2(n_3389),
.B1(n_3531),
.B2(n_3475),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_3898),
.Y(n_4248)
);

INVx4_ASAP7_75t_L g4249 ( 
.A(n_4027),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_3855),
.Y(n_4250)
);

INVx4_ASAP7_75t_L g4251 ( 
.A(n_4038),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_3910),
.Y(n_4252)
);

INVx2_ASAP7_75t_SL g4253 ( 
.A(n_3978),
.Y(n_4253)
);

INVx6_ASAP7_75t_L g4254 ( 
.A(n_3775),
.Y(n_4254)
);

INVx1_ASAP7_75t_SL g4255 ( 
.A(n_3921),
.Y(n_4255)
);

CKINVDCx16_ASAP7_75t_R g4256 ( 
.A(n_3872),
.Y(n_4256)
);

CKINVDCx5p33_ASAP7_75t_R g4257 ( 
.A(n_3930),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_3938),
.Y(n_4258)
);

AOI22xp33_ASAP7_75t_L g4259 ( 
.A1(n_3837),
.A2(n_3389),
.B1(n_3531),
.B2(n_3475),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_3748),
.B(n_4041),
.Y(n_4260)
);

CKINVDCx20_ASAP7_75t_R g4261 ( 
.A(n_3841),
.Y(n_4261)
);

OR2x2_ASAP7_75t_L g4262 ( 
.A(n_3938),
.B(n_607),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_3937),
.B(n_608),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3944),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_3859),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_3958),
.Y(n_4266)
);

AOI22xp33_ASAP7_75t_L g4267 ( 
.A1(n_3793),
.A2(n_3798),
.B1(n_3982),
.B2(n_3972),
.Y(n_4267)
);

CKINVDCx5p33_ASAP7_75t_R g4268 ( 
.A(n_3985),
.Y(n_4268)
);

INVx2_ASAP7_75t_SL g4269 ( 
.A(n_3944),
.Y(n_4269)
);

BUFx6f_ASAP7_75t_L g4270 ( 
.A(n_3763),
.Y(n_4270)
);

BUFx3_ASAP7_75t_L g4271 ( 
.A(n_3779),
.Y(n_4271)
);

AOI22xp33_ASAP7_75t_L g4272 ( 
.A1(n_3987),
.A2(n_3531),
.B1(n_3612),
.B2(n_3534),
.Y(n_4272)
);

BUFx6f_ASAP7_75t_L g4273 ( 
.A(n_3762),
.Y(n_4273)
);

BUFx10_ASAP7_75t_L g4274 ( 
.A(n_3858),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_4094),
.B(n_3858),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4089),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_L g4277 ( 
.A(n_4169),
.B(n_3766),
.Y(n_4277)
);

BUFx2_ASAP7_75t_L g4278 ( 
.A(n_4188),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4091),
.Y(n_4279)
);

AND2x4_ASAP7_75t_L g4280 ( 
.A(n_4194),
.B(n_3988),
.Y(n_4280)
);

INVx2_ASAP7_75t_SL g4281 ( 
.A(n_4129),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4075),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4084),
.Y(n_4283)
);

BUFx2_ASAP7_75t_L g4284 ( 
.A(n_4188),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4087),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_4103),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_4107),
.Y(n_4287)
);

AND2x2_ASAP7_75t_L g4288 ( 
.A(n_4125),
.B(n_3861),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4090),
.Y(n_4289)
);

INVx2_ASAP7_75t_L g4290 ( 
.A(n_4110),
.Y(n_4290)
);

HB1xp67_ASAP7_75t_L g4291 ( 
.A(n_4227),
.Y(n_4291)
);

OAI21xp5_ASAP7_75t_L g4292 ( 
.A1(n_4148),
.A2(n_3949),
.B(n_4018),
.Y(n_4292)
);

BUFx2_ASAP7_75t_L g4293 ( 
.A(n_4194),
.Y(n_4293)
);

OR2x6_ASAP7_75t_L g4294 ( 
.A(n_4088),
.B(n_4007),
.Y(n_4294)
);

OAI21x1_ASAP7_75t_L g4295 ( 
.A1(n_4246),
.A2(n_3952),
.B(n_3741),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4115),
.Y(n_4296)
);

AOI221xp5_ASAP7_75t_L g4297 ( 
.A1(n_4170),
.A2(n_4214),
.B1(n_4263),
.B2(n_4111),
.C(n_4168),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4136),
.Y(n_4298)
);

OAI21x1_ASAP7_75t_L g4299 ( 
.A1(n_4266),
.A2(n_3753),
.B(n_3746),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4138),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4146),
.Y(n_4301)
);

INVx2_ASAP7_75t_L g4302 ( 
.A(n_4120),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4150),
.Y(n_4303)
);

AND2x2_ASAP7_75t_L g4304 ( 
.A(n_4208),
.B(n_3861),
.Y(n_4304)
);

INVx2_ASAP7_75t_SL g4305 ( 
.A(n_4129),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4159),
.Y(n_4306)
);

INVx3_ASAP7_75t_L g4307 ( 
.A(n_4067),
.Y(n_4307)
);

INVxp67_ASAP7_75t_L g4308 ( 
.A(n_4153),
.Y(n_4308)
);

OR2x2_ASAP7_75t_L g4309 ( 
.A(n_4133),
.B(n_4139),
.Y(n_4309)
);

BUFx3_ASAP7_75t_L g4310 ( 
.A(n_4143),
.Y(n_4310)
);

INVx2_ASAP7_75t_L g4311 ( 
.A(n_4121),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4164),
.Y(n_4312)
);

BUFx2_ASAP7_75t_L g4313 ( 
.A(n_4232),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_4128),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4167),
.Y(n_4315)
);

INVx3_ASAP7_75t_L g4316 ( 
.A(n_4074),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_4130),
.Y(n_4317)
);

OAI21xp5_ASAP7_75t_L g4318 ( 
.A1(n_4157),
.A2(n_4025),
.B(n_4058),
.Y(n_4318)
);

CKINVDCx20_ASAP7_75t_R g4319 ( 
.A(n_4081),
.Y(n_4319)
);

INVx3_ASAP7_75t_L g4320 ( 
.A(n_4155),
.Y(n_4320)
);

INVx3_ASAP7_75t_L g4321 ( 
.A(n_4124),
.Y(n_4321)
);

HB1xp67_ASAP7_75t_L g4322 ( 
.A(n_4213),
.Y(n_4322)
);

BUFx6f_ASAP7_75t_L g4323 ( 
.A(n_4162),
.Y(n_4323)
);

AOI22xp33_ASAP7_75t_L g4324 ( 
.A1(n_4073),
.A2(n_3953),
.B1(n_3915),
.B2(n_3780),
.Y(n_4324)
);

AOI22xp33_ASAP7_75t_L g4325 ( 
.A1(n_4235),
.A2(n_3836),
.B1(n_3754),
.B2(n_3797),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4172),
.Y(n_4326)
);

BUFx3_ASAP7_75t_L g4327 ( 
.A(n_4114),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4174),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4203),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4217),
.B(n_3853),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_4158),
.Y(n_4331)
);

CKINVDCx5p33_ASAP7_75t_R g4332 ( 
.A(n_4185),
.Y(n_4332)
);

HB1xp67_ASAP7_75t_L g4333 ( 
.A(n_4160),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4219),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4140),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4221),
.Y(n_4336)
);

INVx3_ASAP7_75t_L g4337 ( 
.A(n_4209),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4222),
.Y(n_4338)
);

BUFx6f_ASAP7_75t_L g4339 ( 
.A(n_4162),
.Y(n_4339)
);

INVx2_ASAP7_75t_L g4340 ( 
.A(n_4186),
.Y(n_4340)
);

OAI21x1_ASAP7_75t_L g4341 ( 
.A1(n_4265),
.A2(n_3755),
.B(n_3807),
.Y(n_4341)
);

BUFx6f_ASAP7_75t_L g4342 ( 
.A(n_4113),
.Y(n_4342)
);

BUFx12f_ASAP7_75t_L g4343 ( 
.A(n_4102),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4224),
.Y(n_4344)
);

HB1xp67_ASAP7_75t_L g4345 ( 
.A(n_4100),
.Y(n_4345)
);

INVx3_ASAP7_75t_L g4346 ( 
.A(n_4209),
.Y(n_4346)
);

HB1xp67_ASAP7_75t_L g4347 ( 
.A(n_4202),
.Y(n_4347)
);

INVx5_ASAP7_75t_L g4348 ( 
.A(n_4088),
.Y(n_4348)
);

OAI22xp5_ASAP7_75t_L g4349 ( 
.A1(n_4256),
.A2(n_3852),
.B1(n_3860),
.B2(n_3905),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4223),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4226),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4141),
.B(n_3853),
.Y(n_4352)
);

INVx2_ASAP7_75t_L g4353 ( 
.A(n_4269),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_4236),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_L g4355 ( 
.A(n_4239),
.B(n_4242),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_4238),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4274),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4258),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4264),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4082),
.Y(n_4360)
);

OA21x2_ASAP7_75t_L g4361 ( 
.A1(n_4247),
.A2(n_3999),
.B(n_3773),
.Y(n_4361)
);

BUFx12f_ASAP7_75t_L g4362 ( 
.A(n_4080),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4184),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4197),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4250),
.Y(n_4365)
);

INVx3_ASAP7_75t_L g4366 ( 
.A(n_4231),
.Y(n_4366)
);

AOI22xp5_ASAP7_75t_L g4367 ( 
.A1(n_4105),
.A2(n_3850),
.B1(n_3884),
.B2(n_3874),
.Y(n_4367)
);

HB1xp67_ASAP7_75t_L g4368 ( 
.A(n_4166),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4245),
.Y(n_4369)
);

INVx2_ASAP7_75t_L g4370 ( 
.A(n_4262),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4248),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4252),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_4249),
.Y(n_4373)
);

O2A1O1Ixp33_ASAP7_75t_L g4374 ( 
.A1(n_4144),
.A2(n_3913),
.B(n_3990),
.C(n_3945),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4216),
.Y(n_4375)
);

HB1xp67_ASAP7_75t_L g4376 ( 
.A(n_4154),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4251),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4154),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4228),
.Y(n_4379)
);

INVx3_ASAP7_75t_L g4380 ( 
.A(n_4231),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4204),
.B(n_4001),
.Y(n_4381)
);

AND2x2_ASAP7_75t_L g4382 ( 
.A(n_4066),
.B(n_3862),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_4177),
.Y(n_4383)
);

INVx3_ASAP7_75t_L g4384 ( 
.A(n_4240),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_4177),
.Y(n_4385)
);

HB1xp67_ASAP7_75t_L g4386 ( 
.A(n_4175),
.Y(n_4386)
);

AOI22xp33_ASAP7_75t_L g4387 ( 
.A1(n_4096),
.A2(n_4048),
.B1(n_4055),
.B2(n_4024),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_4255),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4254),
.Y(n_4389)
);

OA21x2_ASAP7_75t_L g4390 ( 
.A1(n_4218),
.A2(n_3769),
.B(n_4021),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4254),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4127),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4243),
.Y(n_4393)
);

AO31x2_ASAP7_75t_L g4394 ( 
.A1(n_4260),
.A2(n_3744),
.A3(n_3812),
.B(n_4035),
.Y(n_4394)
);

INVx8_ASAP7_75t_L g4395 ( 
.A(n_4112),
.Y(n_4395)
);

OR2x2_ASAP7_75t_L g4396 ( 
.A(n_4253),
.B(n_4001),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4220),
.Y(n_4397)
);

INVx2_ASAP7_75t_L g4398 ( 
.A(n_4243),
.Y(n_4398)
);

OAI21x1_ASAP7_75t_L g4399 ( 
.A1(n_4259),
.A2(n_3813),
.B(n_3783),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4198),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4198),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_4069),
.B(n_4062),
.Y(n_4402)
);

BUFx6f_ASAP7_75t_L g4403 ( 
.A(n_4113),
.Y(n_4403)
);

BUFx2_ASAP7_75t_L g4404 ( 
.A(n_4271),
.Y(n_4404)
);

OAI21x1_ASAP7_75t_L g4405 ( 
.A1(n_4272),
.A2(n_3968),
.B(n_3881),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4175),
.Y(n_4406)
);

INVx2_ASAP7_75t_L g4407 ( 
.A(n_4273),
.Y(n_4407)
);

BUFx2_ASAP7_75t_L g4408 ( 
.A(n_4240),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4193),
.Y(n_4409)
);

AO21x2_ASAP7_75t_L g4410 ( 
.A1(n_4071),
.A2(n_3919),
.B(n_3848),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4212),
.Y(n_4411)
);

INVx2_ASAP7_75t_L g4412 ( 
.A(n_4273),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4196),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4196),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4076),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4190),
.Y(n_4416)
);

AND2x2_ASAP7_75t_L g4417 ( 
.A(n_4261),
.B(n_3862),
.Y(n_4417)
);

OA21x2_ASAP7_75t_L g4418 ( 
.A1(n_4357),
.A2(n_4267),
.B(n_4205),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4282),
.Y(n_4419)
);

A2O1A1Ixp33_ASAP7_75t_L g4420 ( 
.A1(n_4297),
.A2(n_4152),
.B(n_4095),
.C(n_4173),
.Y(n_4420)
);

AOI22xp33_ASAP7_75t_L g4421 ( 
.A1(n_4349),
.A2(n_4417),
.B1(n_4292),
.B2(n_4382),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4275),
.B(n_4181),
.Y(n_4422)
);

AND2x2_ASAP7_75t_L g4423 ( 
.A(n_4291),
.B(n_4234),
.Y(n_4423)
);

INVx6_ASAP7_75t_L g4424 ( 
.A(n_4348),
.Y(n_4424)
);

OA21x2_ASAP7_75t_L g4425 ( 
.A1(n_4402),
.A2(n_4277),
.B(n_4373),
.Y(n_4425)
);

AO21x1_ASAP7_75t_L g4426 ( 
.A1(n_4276),
.A2(n_4101),
.B(n_4123),
.Y(n_4426)
);

INVx2_ASAP7_75t_SL g4427 ( 
.A(n_4348),
.Y(n_4427)
);

AO21x1_ASAP7_75t_L g4428 ( 
.A1(n_4335),
.A2(n_4119),
.B(n_4176),
.Y(n_4428)
);

BUFx6f_ASAP7_75t_L g4429 ( 
.A(n_4323),
.Y(n_4429)
);

OR2x2_ASAP7_75t_L g4430 ( 
.A(n_4345),
.B(n_4147),
.Y(n_4430)
);

AND2x4_ASAP7_75t_L g4431 ( 
.A(n_4348),
.B(n_4068),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4383),
.B(n_4093),
.Y(n_4432)
);

OR2x2_ASAP7_75t_L g4433 ( 
.A(n_4347),
.B(n_4135),
.Y(n_4433)
);

INVx2_ASAP7_75t_SL g4434 ( 
.A(n_4323),
.Y(n_4434)
);

OA21x2_ASAP7_75t_L g4435 ( 
.A1(n_4377),
.A2(n_4099),
.B(n_4225),
.Y(n_4435)
);

NOR3xp33_ASAP7_75t_SL g4436 ( 
.A(n_4332),
.B(n_4131),
.C(n_4268),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4385),
.B(n_4135),
.Y(n_4437)
);

INVxp67_ASAP7_75t_SL g4438 ( 
.A(n_4309),
.Y(n_4438)
);

NOR2x1_ASAP7_75t_SL g4439 ( 
.A(n_4294),
.B(n_4362),
.Y(n_4439)
);

OAI22xp5_ASAP7_75t_L g4440 ( 
.A1(n_4308),
.A2(n_4092),
.B1(n_4142),
.B2(n_4086),
.Y(n_4440)
);

NAND2x1_ASAP7_75t_L g4441 ( 
.A(n_4293),
.B(n_4080),
.Y(n_4441)
);

O2A1O1Ixp33_ASAP7_75t_SL g4442 ( 
.A1(n_4386),
.A2(n_4215),
.B(n_4077),
.C(n_4165),
.Y(n_4442)
);

OAI22xp5_ASAP7_75t_L g4443 ( 
.A1(n_4294),
.A2(n_4237),
.B1(n_4079),
.B2(n_4134),
.Y(n_4443)
);

AND2x2_ASAP7_75t_L g4444 ( 
.A(n_4389),
.B(n_4070),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4283),
.Y(n_4445)
);

OR2x6_ASAP7_75t_L g4446 ( 
.A(n_4395),
.B(n_4072),
.Y(n_4446)
);

OAI21xp5_ASAP7_75t_L g4447 ( 
.A1(n_4318),
.A2(n_4098),
.B(n_4083),
.Y(n_4447)
);

AND2x2_ASAP7_75t_L g4448 ( 
.A(n_4391),
.B(n_4070),
.Y(n_4448)
);

A2O1A1Ixp33_ASAP7_75t_L g4449 ( 
.A1(n_4320),
.A2(n_3917),
.B(n_4156),
.C(n_4230),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_4285),
.Y(n_4450)
);

A2O1A1Ixp33_ASAP7_75t_L g4451 ( 
.A1(n_4374),
.A2(n_4106),
.B(n_4257),
.C(n_4244),
.Y(n_4451)
);

AND2x2_ASAP7_75t_L g4452 ( 
.A(n_4368),
.B(n_4333),
.Y(n_4452)
);

OAI22xp5_ASAP7_75t_L g4453 ( 
.A1(n_4387),
.A2(n_4104),
.B1(n_4229),
.B2(n_4137),
.Y(n_4453)
);

AND2x4_ASAP7_75t_L g4454 ( 
.A(n_4278),
.B(n_4270),
.Y(n_4454)
);

AND2x2_ASAP7_75t_L g4455 ( 
.A(n_4388),
.B(n_4241),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_4360),
.B(n_4201),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4289),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4352),
.B(n_4211),
.Y(n_4458)
);

AOI221xp5_ASAP7_75t_L g4459 ( 
.A1(n_4392),
.A2(n_4233),
.B1(n_4132),
.B2(n_4118),
.C(n_4122),
.Y(n_4459)
);

BUFx12f_ASAP7_75t_L g4460 ( 
.A(n_4343),
.Y(n_4460)
);

AND2x2_ASAP7_75t_L g4461 ( 
.A(n_4369),
.B(n_4270),
.Y(n_4461)
);

AND2x2_ASAP7_75t_L g4462 ( 
.A(n_4371),
.B(n_4200),
.Y(n_4462)
);

AND2x6_ASAP7_75t_L g4463 ( 
.A(n_4280),
.B(n_4117),
.Y(n_4463)
);

OA21x2_ASAP7_75t_L g4464 ( 
.A1(n_4293),
.A2(n_4206),
.B(n_3818),
.Y(n_4464)
);

AND2x2_ASAP7_75t_L g4465 ( 
.A(n_4372),
.B(n_4413),
.Y(n_4465)
);

AOI22xp5_ASAP7_75t_L g4466 ( 
.A1(n_4411),
.A2(n_4078),
.B1(n_4097),
.B2(n_4108),
.Y(n_4466)
);

AOI221xp5_ASAP7_75t_L g4467 ( 
.A1(n_4381),
.A2(n_4006),
.B1(n_4015),
.B2(n_4005),
.C(n_4004),
.Y(n_4467)
);

OAI21xp5_ASAP7_75t_L g4468 ( 
.A1(n_4325),
.A2(n_4020),
.B(n_4016),
.Y(n_4468)
);

AND2x4_ASAP7_75t_L g4469 ( 
.A(n_4278),
.B(n_4109),
.Y(n_4469)
);

OR2x2_ASAP7_75t_L g4470 ( 
.A(n_4296),
.B(n_4151),
.Y(n_4470)
);

OA21x2_ASAP7_75t_L g4471 ( 
.A1(n_4295),
.A2(n_4145),
.B(n_4023),
.Y(n_4471)
);

OA21x2_ASAP7_75t_L g4472 ( 
.A1(n_4404),
.A2(n_4149),
.B(n_3894),
.Y(n_4472)
);

OAI211xp5_ASAP7_75t_L g4473 ( 
.A1(n_4367),
.A2(n_4324),
.B(n_4379),
.C(n_4376),
.Y(n_4473)
);

AND2x4_ASAP7_75t_L g4474 ( 
.A(n_4284),
.B(n_4323),
.Y(n_4474)
);

CKINVDCx20_ASAP7_75t_R g4475 ( 
.A(n_4319),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4414),
.B(n_4298),
.Y(n_4476)
);

AND2x2_ASAP7_75t_L g4477 ( 
.A(n_4300),
.B(n_4301),
.Y(n_4477)
);

AND2x4_ASAP7_75t_SL g4478 ( 
.A(n_4307),
.B(n_4171),
.Y(n_4478)
);

INVxp67_ASAP7_75t_L g4479 ( 
.A(n_4397),
.Y(n_4479)
);

AND2x4_ASAP7_75t_L g4480 ( 
.A(n_4284),
.B(n_3842),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_L g4481 ( 
.A(n_4288),
.B(n_4179),
.Y(n_4481)
);

AOI21xp5_ASAP7_75t_L g4482 ( 
.A1(n_4280),
.A2(n_4410),
.B(n_4408),
.Y(n_4482)
);

BUFx6f_ASAP7_75t_L g4483 ( 
.A(n_4339),
.Y(n_4483)
);

AND2x4_ASAP7_75t_L g4484 ( 
.A(n_4339),
.B(n_3842),
.Y(n_4484)
);

AND2x2_ASAP7_75t_L g4485 ( 
.A(n_4303),
.B(n_3886),
.Y(n_4485)
);

OAI21xp5_ASAP7_75t_L g4486 ( 
.A1(n_4316),
.A2(n_4061),
.B(n_4057),
.Y(n_4486)
);

INVxp67_ASAP7_75t_L g4487 ( 
.A(n_4339),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4306),
.B(n_3886),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_4304),
.B(n_4116),
.Y(n_4489)
);

BUFx5_ASAP7_75t_L g4490 ( 
.A(n_4415),
.Y(n_4490)
);

OAI221xp5_ASAP7_75t_L g4491 ( 
.A1(n_4400),
.A2(n_4189),
.B1(n_4163),
.B2(n_4180),
.C(n_4161),
.Y(n_4491)
);

BUFx2_ASAP7_75t_L g4492 ( 
.A(n_4342),
.Y(n_4492)
);

A2O1A1Ixp33_ASAP7_75t_L g4493 ( 
.A1(n_4406),
.A2(n_3757),
.B(n_3907),
.C(n_3888),
.Y(n_4493)
);

AND2x4_ASAP7_75t_L g4494 ( 
.A(n_4378),
.B(n_4062),
.Y(n_4494)
);

AND2x2_ASAP7_75t_L g4495 ( 
.A(n_4312),
.B(n_3743),
.Y(n_4495)
);

OAI21xp5_ASAP7_75t_L g4496 ( 
.A1(n_4396),
.A2(n_3922),
.B(n_3908),
.Y(n_4496)
);

AND2x4_ASAP7_75t_L g4497 ( 
.A(n_4366),
.B(n_3534),
.Y(n_4497)
);

NOR2x1_ASAP7_75t_SL g4498 ( 
.A(n_4310),
.B(n_4085),
.Y(n_4498)
);

NOR2x1_ASAP7_75t_SL g4499 ( 
.A(n_4401),
.B(n_4126),
.Y(n_4499)
);

OR2x2_ASAP7_75t_L g4500 ( 
.A(n_4315),
.B(n_3743),
.Y(n_4500)
);

AND2x4_ASAP7_75t_L g4501 ( 
.A(n_4366),
.B(n_3534),
.Y(n_4501)
);

AOI221xp5_ASAP7_75t_L g4502 ( 
.A1(n_4370),
.A2(n_4192),
.B1(n_4191),
.B2(n_3896),
.C(n_3925),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4326),
.B(n_3738),
.Y(n_4503)
);

AOI22xp5_ASAP7_75t_L g4504 ( 
.A1(n_4330),
.A2(n_4182),
.B1(n_4199),
.B2(n_4187),
.Y(n_4504)
);

OAI22xp5_ASAP7_75t_SL g4505 ( 
.A1(n_4321),
.A2(n_4072),
.B1(n_4178),
.B2(n_3864),
.Y(n_4505)
);

OR2x2_ASAP7_75t_L g4506 ( 
.A(n_4438),
.B(n_4375),
.Y(n_4506)
);

AND2x2_ASAP7_75t_L g4507 ( 
.A(n_4452),
.B(n_4458),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4423),
.B(n_4409),
.Y(n_4508)
);

INVx2_ASAP7_75t_L g4509 ( 
.A(n_4430),
.Y(n_4509)
);

INVx3_ASAP7_75t_L g4510 ( 
.A(n_4463),
.Y(n_4510)
);

OR2x2_ASAP7_75t_L g4511 ( 
.A(n_4489),
.B(n_4363),
.Y(n_4511)
);

BUFx6f_ASAP7_75t_L g4512 ( 
.A(n_4429),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_4432),
.B(n_4416),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4419),
.Y(n_4514)
);

AND2x2_ASAP7_75t_L g4515 ( 
.A(n_4476),
.B(n_4322),
.Y(n_4515)
);

AND2x2_ASAP7_75t_L g4516 ( 
.A(n_4425),
.B(n_4364),
.Y(n_4516)
);

INVx2_ASAP7_75t_SL g4517 ( 
.A(n_4446),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4445),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4495),
.B(n_4328),
.Y(n_4519)
);

BUFx2_ASAP7_75t_L g4520 ( 
.A(n_4463),
.Y(n_4520)
);

HB1xp67_ASAP7_75t_L g4521 ( 
.A(n_4433),
.Y(n_4521)
);

AND2x2_ASAP7_75t_SL g4522 ( 
.A(n_4431),
.B(n_4408),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4450),
.Y(n_4523)
);

INVx2_ASAP7_75t_L g4524 ( 
.A(n_4490),
.Y(n_4524)
);

AND2x4_ASAP7_75t_L g4525 ( 
.A(n_4480),
.B(n_4454),
.Y(n_4525)
);

INVx2_ASAP7_75t_L g4526 ( 
.A(n_4490),
.Y(n_4526)
);

AND2x2_ASAP7_75t_L g4527 ( 
.A(n_4437),
.B(n_4337),
.Y(n_4527)
);

AND2x2_ASAP7_75t_L g4528 ( 
.A(n_4465),
.B(n_4337),
.Y(n_4528)
);

NOR2xp33_ASAP7_75t_L g4529 ( 
.A(n_4479),
.B(n_4346),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4457),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_4503),
.B(n_4329),
.Y(n_4531)
);

NAND2xp5_ASAP7_75t_L g4532 ( 
.A(n_4422),
.B(n_4334),
.Y(n_4532)
);

INVx2_ASAP7_75t_SL g4533 ( 
.A(n_4446),
.Y(n_4533)
);

INVx2_ASAP7_75t_L g4534 ( 
.A(n_4490),
.Y(n_4534)
);

AND2x4_ASAP7_75t_L g4535 ( 
.A(n_4461),
.B(n_4353),
.Y(n_4535)
);

INVxp67_ASAP7_75t_L g4536 ( 
.A(n_4418),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4477),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_4500),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_SL g4539 ( 
.A(n_4426),
.B(n_4342),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4485),
.Y(n_4540)
);

INVx2_ASAP7_75t_L g4541 ( 
.A(n_4492),
.Y(n_4541)
);

AOI221xp5_ASAP7_75t_L g4542 ( 
.A1(n_4447),
.A2(n_4355),
.B1(n_4338),
.B2(n_4344),
.C(n_4336),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_4488),
.B(n_4350),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4481),
.Y(n_4544)
);

INVxp67_ASAP7_75t_SL g4545 ( 
.A(n_4428),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4444),
.B(n_4448),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4462),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4456),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4470),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4455),
.B(n_4346),
.Y(n_4550)
);

INVxp67_ASAP7_75t_L g4551 ( 
.A(n_4435),
.Y(n_4551)
);

BUFx2_ASAP7_75t_L g4552 ( 
.A(n_4463),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4469),
.B(n_4404),
.Y(n_4553)
);

INVx2_ASAP7_75t_L g4554 ( 
.A(n_4474),
.Y(n_4554)
);

OAI22xp5_ASAP7_75t_L g4555 ( 
.A1(n_4421),
.A2(n_4384),
.B1(n_4351),
.B2(n_4380),
.Y(n_4555)
);

OR2x2_ASAP7_75t_L g4556 ( 
.A(n_4487),
.B(n_4354),
.Y(n_4556)
);

NAND2xp5_ASAP7_75t_L g4557 ( 
.A(n_4494),
.B(n_4358),
.Y(n_4557)
);

AND2x2_ASAP7_75t_L g4558 ( 
.A(n_4434),
.B(n_4393),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4504),
.B(n_4359),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4441),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4484),
.B(n_4398),
.Y(n_4561)
);

INVx3_ASAP7_75t_L g4562 ( 
.A(n_4424),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4482),
.B(n_4313),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4439),
.B(n_4313),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4473),
.Y(n_4565)
);

HB1xp67_ASAP7_75t_L g4566 ( 
.A(n_4472),
.Y(n_4566)
);

HB1xp67_ASAP7_75t_L g4567 ( 
.A(n_4471),
.Y(n_4567)
);

AND2x2_ASAP7_75t_L g4568 ( 
.A(n_4429),
.B(n_4279),
.Y(n_4568)
);

INVx2_ASAP7_75t_L g4569 ( 
.A(n_4483),
.Y(n_4569)
);

AND2x2_ASAP7_75t_L g4570 ( 
.A(n_4483),
.B(n_4286),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4424),
.Y(n_4571)
);

OAI22xp33_ASAP7_75t_L g4572 ( 
.A1(n_4443),
.A2(n_4384),
.B1(n_4395),
.B2(n_4380),
.Y(n_4572)
);

INVx3_ASAP7_75t_L g4573 ( 
.A(n_4427),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4464),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4491),
.Y(n_4575)
);

INVx2_ASAP7_75t_SL g4576 ( 
.A(n_4478),
.Y(n_4576)
);

AOI22xp33_ASAP7_75t_L g4577 ( 
.A1(n_4453),
.A2(n_4459),
.B1(n_4440),
.B2(n_4466),
.Y(n_4577)
);

AOI33xp33_ASAP7_75t_L g4578 ( 
.A1(n_4577),
.A2(n_4442),
.A3(n_4502),
.B1(n_4305),
.B2(n_4281),
.B3(n_4467),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_4544),
.B(n_4394),
.Y(n_4579)
);

INVx2_ASAP7_75t_L g4580 ( 
.A(n_4516),
.Y(n_4580)
);

INVx2_ASAP7_75t_L g4581 ( 
.A(n_4521),
.Y(n_4581)
);

INVx3_ASAP7_75t_L g4582 ( 
.A(n_4510),
.Y(n_4582)
);

INVx2_ASAP7_75t_L g4583 ( 
.A(n_4521),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4553),
.B(n_4407),
.Y(n_4584)
);

AND2x2_ASAP7_75t_L g4585 ( 
.A(n_4546),
.B(n_4412),
.Y(n_4585)
);

INVx4_ASAP7_75t_L g4586 ( 
.A(n_4510),
.Y(n_4586)
);

AO21x2_ASAP7_75t_L g4587 ( 
.A1(n_4545),
.A2(n_4420),
.B(n_4451),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4514),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4556),
.Y(n_4589)
);

NAND4xp25_ASAP7_75t_L g4590 ( 
.A(n_4577),
.B(n_4449),
.C(n_4468),
.D(n_4486),
.Y(n_4590)
);

AND2x2_ASAP7_75t_L g4591 ( 
.A(n_4528),
.B(n_4499),
.Y(n_4591)
);

BUFx3_ASAP7_75t_L g4592 ( 
.A(n_4576),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4559),
.B(n_4394),
.Y(n_4593)
);

NAND2xp5_ASAP7_75t_L g4594 ( 
.A(n_4559),
.B(n_4394),
.Y(n_4594)
);

INVx2_ASAP7_75t_L g4595 ( 
.A(n_4538),
.Y(n_4595)
);

INVx4_ASAP7_75t_L g4596 ( 
.A(n_4520),
.Y(n_4596)
);

INVxp67_ASAP7_75t_L g4597 ( 
.A(n_4529),
.Y(n_4597)
);

OAI21x1_ASAP7_75t_L g4598 ( 
.A1(n_4573),
.A2(n_4399),
.B(n_4299),
.Y(n_4598)
);

INVx2_ASAP7_75t_SL g4599 ( 
.A(n_4517),
.Y(n_4599)
);

HB1xp67_ASAP7_75t_L g4600 ( 
.A(n_4506),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4507),
.B(n_4287),
.Y(n_4601)
);

INVx5_ASAP7_75t_SL g4602 ( 
.A(n_4522),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4547),
.B(n_4290),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4527),
.B(n_4302),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4518),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4523),
.Y(n_4606)
);

INVx2_ASAP7_75t_L g4607 ( 
.A(n_4535),
.Y(n_4607)
);

OR2x2_ASAP7_75t_L g4608 ( 
.A(n_4511),
.B(n_4356),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4530),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4543),
.Y(n_4610)
);

NOR2x1_ASAP7_75t_R g4611 ( 
.A(n_4552),
.B(n_4460),
.Y(n_4611)
);

OAI31xp33_ASAP7_75t_L g4612 ( 
.A1(n_4572),
.A2(n_4545),
.A3(n_4565),
.B(n_4555),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4543),
.Y(n_4613)
);

INVxp67_ASAP7_75t_L g4614 ( 
.A(n_4533),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4519),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4535),
.Y(n_4616)
);

INVxp67_ASAP7_75t_SL g4617 ( 
.A(n_4573),
.Y(n_4617)
);

AOI22xp33_ASAP7_75t_L g4618 ( 
.A1(n_4575),
.A2(n_4505),
.B1(n_4496),
.B2(n_4390),
.Y(n_4618)
);

INVx3_ASAP7_75t_L g4619 ( 
.A(n_4564),
.Y(n_4619)
);

HB1xp67_ASAP7_75t_L g4620 ( 
.A(n_4509),
.Y(n_4620)
);

AOI221xp5_ASAP7_75t_L g4621 ( 
.A1(n_4572),
.A2(n_4493),
.B1(n_4053),
.B2(n_3931),
.C(n_3969),
.Y(n_4621)
);

OR2x2_ASAP7_75t_L g4622 ( 
.A(n_4540),
.B(n_4311),
.Y(n_4622)
);

AOI22xp5_ASAP7_75t_L g4623 ( 
.A1(n_4555),
.A2(n_4542),
.B1(n_4536),
.B2(n_4539),
.Y(n_4623)
);

OAI321xp33_ASAP7_75t_L g4624 ( 
.A1(n_4536),
.A2(n_4403),
.A3(n_4342),
.B1(n_4331),
.B2(n_4314),
.C(n_4340),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4519),
.Y(n_4625)
);

OR2x2_ASAP7_75t_L g4626 ( 
.A(n_4532),
.B(n_4317),
.Y(n_4626)
);

OR2x2_ASAP7_75t_L g4627 ( 
.A(n_4532),
.B(n_4365),
.Y(n_4627)
);

BUFx2_ASAP7_75t_L g4628 ( 
.A(n_4562),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_4542),
.B(n_4390),
.Y(n_4629)
);

NAND2x1p5_ASAP7_75t_L g4630 ( 
.A(n_4562),
.B(n_4327),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4554),
.B(n_4436),
.Y(n_4631)
);

OR2x2_ASAP7_75t_L g4632 ( 
.A(n_4537),
.B(n_4361),
.Y(n_4632)
);

INVx2_ASAP7_75t_L g4633 ( 
.A(n_4557),
.Y(n_4633)
);

OR2x2_ASAP7_75t_L g4634 ( 
.A(n_4531),
.B(n_4361),
.Y(n_4634)
);

NAND3xp33_ASAP7_75t_L g4635 ( 
.A(n_4551),
.B(n_4195),
.C(n_4403),
.Y(n_4635)
);

AND2x2_ASAP7_75t_L g4636 ( 
.A(n_4515),
.B(n_4498),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4541),
.B(n_4497),
.Y(n_4637)
);

AND2x4_ASAP7_75t_L g4638 ( 
.A(n_4560),
.B(n_4403),
.Y(n_4638)
);

AND2x2_ASAP7_75t_L g4639 ( 
.A(n_4549),
.B(n_4501),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_4615),
.B(n_4551),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4580),
.Y(n_4641)
);

OR2x2_ASAP7_75t_L g4642 ( 
.A(n_4634),
.B(n_4531),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4610),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4610),
.Y(n_4644)
);

NAND3xp33_ASAP7_75t_L g4645 ( 
.A(n_4612),
.B(n_4567),
.C(n_4566),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4619),
.B(n_4525),
.Y(n_4646)
);

INVx3_ASAP7_75t_L g4647 ( 
.A(n_4602),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4613),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4613),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4619),
.B(n_4525),
.Y(n_4650)
);

HB1xp67_ASAP7_75t_L g4651 ( 
.A(n_4600),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4596),
.B(n_4550),
.Y(n_4652)
);

OR2x2_ASAP7_75t_L g4653 ( 
.A(n_4632),
.B(n_4557),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4626),
.Y(n_4654)
);

AND2x2_ASAP7_75t_L g4655 ( 
.A(n_4596),
.B(n_4571),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4602),
.B(n_4513),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4627),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4628),
.B(n_4508),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4605),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4605),
.Y(n_4660)
);

HB1xp67_ASAP7_75t_L g4661 ( 
.A(n_4581),
.Y(n_4661)
);

AND2x2_ASAP7_75t_L g4662 ( 
.A(n_4631),
.B(n_4548),
.Y(n_4662)
);

OR2x2_ASAP7_75t_L g4663 ( 
.A(n_4579),
.B(n_4615),
.Y(n_4663)
);

AND2x2_ASAP7_75t_L g4664 ( 
.A(n_4582),
.B(n_4599),
.Y(n_4664)
);

AND2x2_ASAP7_75t_L g4665 ( 
.A(n_4582),
.B(n_4563),
.Y(n_4665)
);

NOR2xp33_ASAP7_75t_L g4666 ( 
.A(n_4611),
.B(n_4475),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4625),
.B(n_4567),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_4625),
.B(n_4566),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4614),
.B(n_4568),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_4629),
.B(n_4574),
.Y(n_4670)
);

INVx2_ASAP7_75t_L g4671 ( 
.A(n_4583),
.Y(n_4671)
);

INVxp67_ASAP7_75t_SL g4672 ( 
.A(n_4593),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4586),
.B(n_4570),
.Y(n_4673)
);

OR2x2_ASAP7_75t_L g4674 ( 
.A(n_4608),
.B(n_4620),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4606),
.Y(n_4675)
);

AND2x2_ASAP7_75t_L g4676 ( 
.A(n_4647),
.B(n_4586),
.Y(n_4676)
);

AND2x2_ASAP7_75t_L g4677 ( 
.A(n_4647),
.B(n_4592),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4659),
.Y(n_4678)
);

NAND2xp5_ASAP7_75t_L g4679 ( 
.A(n_4651),
.B(n_4623),
.Y(n_4679)
);

NAND2xp5_ASAP7_75t_L g4680 ( 
.A(n_4672),
.B(n_4618),
.Y(n_4680)
);

NOR3xp33_ASAP7_75t_L g4681 ( 
.A(n_4645),
.B(n_4590),
.C(n_4578),
.Y(n_4681)
);

BUFx3_ASAP7_75t_L g4682 ( 
.A(n_4666),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4654),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4664),
.B(n_4636),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_4674),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4660),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4665),
.B(n_4617),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_4672),
.B(n_4594),
.Y(n_4688)
);

OR2x2_ASAP7_75t_L g4689 ( 
.A(n_4642),
.B(n_4633),
.Y(n_4689)
);

AND2x2_ASAP7_75t_L g4690 ( 
.A(n_4646),
.B(n_4591),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4650),
.B(n_4607),
.Y(n_4691)
);

INVx2_ASAP7_75t_L g4692 ( 
.A(n_4641),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4657),
.B(n_4670),
.Y(n_4693)
);

AND2x2_ASAP7_75t_L g4694 ( 
.A(n_4655),
.B(n_4616),
.Y(n_4694)
);

INVx2_ASAP7_75t_L g4695 ( 
.A(n_4671),
.Y(n_4695)
);

OR2x2_ASAP7_75t_L g4696 ( 
.A(n_4663),
.B(n_4622),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4675),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4652),
.Y(n_4698)
);

AND2x2_ASAP7_75t_L g4699 ( 
.A(n_4673),
.B(n_4597),
.Y(n_4699)
);

OR2x2_ASAP7_75t_L g4700 ( 
.A(n_4640),
.B(n_4589),
.Y(n_4700)
);

NAND2x1_ASAP7_75t_L g4701 ( 
.A(n_4656),
.B(n_4624),
.Y(n_4701)
);

OR2x6_ASAP7_75t_L g4702 ( 
.A(n_4645),
.B(n_4630),
.Y(n_4702)
);

INVxp67_ASAP7_75t_L g4703 ( 
.A(n_4662),
.Y(n_4703)
);

AOI21xp33_ASAP7_75t_L g4704 ( 
.A1(n_4670),
.A2(n_4587),
.B(n_4635),
.Y(n_4704)
);

INVx2_ASAP7_75t_L g4705 ( 
.A(n_4653),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4643),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4644),
.Y(n_4707)
);

INVxp67_ASAP7_75t_SL g4708 ( 
.A(n_4661),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4640),
.B(n_4606),
.Y(n_4709)
);

AOI22xp5_ASAP7_75t_L g4710 ( 
.A1(n_4669),
.A2(n_4639),
.B1(n_4621),
.B2(n_4584),
.Y(n_4710)
);

AND2x2_ASAP7_75t_L g4711 ( 
.A(n_4658),
.B(n_4585),
.Y(n_4711)
);

AND2x2_ASAP7_75t_L g4712 ( 
.A(n_4661),
.B(n_4637),
.Y(n_4712)
);

AND2x4_ASAP7_75t_L g4713 ( 
.A(n_4648),
.B(n_4649),
.Y(n_4713)
);

HB1xp67_ASAP7_75t_L g4714 ( 
.A(n_4668),
.Y(n_4714)
);

INVx2_ASAP7_75t_L g4715 ( 
.A(n_4667),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4667),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4668),
.B(n_4609),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4651),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4651),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4651),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_L g4721 ( 
.A(n_4651),
.B(n_4609),
.Y(n_4721)
);

AOI222xp33_ASAP7_75t_L g4722 ( 
.A1(n_4645),
.A2(n_4588),
.B1(n_4595),
.B2(n_4603),
.C1(n_4638),
.C2(n_4601),
.Y(n_4722)
);

OR2x2_ASAP7_75t_L g4723 ( 
.A(n_4693),
.B(n_4604),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4676),
.B(n_4638),
.Y(n_4724)
);

NAND3xp33_ASAP7_75t_L g4725 ( 
.A(n_4681),
.B(n_4210),
.C(n_3963),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4708),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4718),
.Y(n_4727)
);

HB1xp67_ASAP7_75t_L g4728 ( 
.A(n_4719),
.Y(n_4728)
);

AND2x2_ASAP7_75t_L g4729 ( 
.A(n_4682),
.B(n_4558),
.Y(n_4729)
);

OR2x2_ASAP7_75t_L g4730 ( 
.A(n_4688),
.B(n_4598),
.Y(n_4730)
);

XOR2x2_ASAP7_75t_L g4731 ( 
.A(n_4677),
.B(n_608),
.Y(n_4731)
);

AND2x2_ASAP7_75t_L g4732 ( 
.A(n_4684),
.B(n_4561),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_L g4733 ( 
.A(n_4720),
.B(n_4524),
.Y(n_4733)
);

OAI31xp33_ASAP7_75t_L g4734 ( 
.A1(n_4704),
.A2(n_4526),
.A3(n_4534),
.B(n_4569),
.Y(n_4734)
);

OAI21xp33_ASAP7_75t_L g4735 ( 
.A1(n_4702),
.A2(n_4722),
.B(n_4679),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4685),
.Y(n_4736)
);

XOR2xp5_ASAP7_75t_L g4737 ( 
.A(n_4710),
.B(n_4512),
.Y(n_4737)
);

BUFx12f_ASAP7_75t_L g4738 ( 
.A(n_4702),
.Y(n_4738)
);

OR2x2_ASAP7_75t_L g4739 ( 
.A(n_4705),
.B(n_3738),
.Y(n_4739)
);

AOI32xp33_ASAP7_75t_L g4740 ( 
.A1(n_4680),
.A2(n_4699),
.A3(n_4716),
.B1(n_4687),
.B2(n_4698),
.Y(n_4740)
);

OR2x2_ASAP7_75t_L g4741 ( 
.A(n_4683),
.B(n_4512),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_4690),
.B(n_4512),
.Y(n_4742)
);

INVx2_ASAP7_75t_SL g4743 ( 
.A(n_4712),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4714),
.B(n_3899),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4716),
.B(n_3899),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4703),
.B(n_4405),
.Y(n_4746)
);

AND2x2_ASAP7_75t_L g4747 ( 
.A(n_4711),
.B(n_3808),
.Y(n_4747)
);

AOI21xp5_ASAP7_75t_L g4748 ( 
.A1(n_4701),
.A2(n_4721),
.B(n_4709),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4678),
.Y(n_4749)
);

INVx1_ASAP7_75t_SL g4750 ( 
.A(n_4700),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4715),
.B(n_4713),
.Y(n_4751)
);

NOR2xp33_ASAP7_75t_L g4752 ( 
.A(n_4717),
.B(n_609),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4689),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4678),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4686),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4686),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4691),
.B(n_3808),
.Y(n_4757)
);

AND2x2_ASAP7_75t_L g4758 ( 
.A(n_4694),
.B(n_4341),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4697),
.Y(n_4759)
);

HB1xp67_ASAP7_75t_L g4760 ( 
.A(n_4706),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4692),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4697),
.Y(n_4762)
);

NAND3xp33_ASAP7_75t_L g4763 ( 
.A(n_4706),
.B(n_3971),
.C(n_3942),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4707),
.Y(n_4764)
);

INVx1_ASAP7_75t_SL g4765 ( 
.A(n_4696),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4707),
.Y(n_4766)
);

OR2x6_ASAP7_75t_L g4767 ( 
.A(n_4695),
.B(n_3970),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4713),
.Y(n_4768)
);

AND2x2_ASAP7_75t_L g4769 ( 
.A(n_4676),
.B(n_3764),
.Y(n_4769)
);

OR2x2_ASAP7_75t_L g4770 ( 
.A(n_4693),
.B(n_609),
.Y(n_4770)
);

NAND2x1_ASAP7_75t_SL g4771 ( 
.A(n_4676),
.B(n_3796),
.Y(n_4771)
);

AND2x2_ASAP7_75t_L g4772 ( 
.A(n_4676),
.B(n_3792),
.Y(n_4772)
);

AOI22xp33_ASAP7_75t_L g4773 ( 
.A1(n_4738),
.A2(n_4183),
.B1(n_4207),
.B2(n_3984),
.Y(n_4773)
);

INVxp67_ASAP7_75t_L g4774 ( 
.A(n_4752),
.Y(n_4774)
);

NOR2xp33_ASAP7_75t_L g4775 ( 
.A(n_4735),
.B(n_609),
.Y(n_4775)
);

INVx2_ASAP7_75t_L g4776 ( 
.A(n_4753),
.Y(n_4776)
);

AOI22xp33_ASAP7_75t_L g4777 ( 
.A1(n_4750),
.A2(n_3805),
.B1(n_3785),
.B2(n_3991),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4765),
.B(n_610),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4743),
.Y(n_4779)
);

OR4x1_ASAP7_75t_L g4780 ( 
.A(n_4726),
.B(n_4727),
.C(n_4754),
.D(n_4749),
.Y(n_4780)
);

AND2x4_ASAP7_75t_L g4781 ( 
.A(n_4724),
.B(n_610),
.Y(n_4781)
);

OAI21xp33_ASAP7_75t_L g4782 ( 
.A1(n_4740),
.A2(n_3820),
.B(n_3821),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4726),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4742),
.B(n_610),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4728),
.B(n_4736),
.Y(n_4785)
);

AOI22xp5_ASAP7_75t_L g4786 ( 
.A1(n_4725),
.A2(n_3791),
.B1(n_3751),
.B2(n_3903),
.Y(n_4786)
);

OAI22xp33_ASAP7_75t_L g4787 ( 
.A1(n_4768),
.A2(n_3828),
.B1(n_3633),
.B2(n_3653),
.Y(n_4787)
);

INVx2_ASAP7_75t_L g4788 ( 
.A(n_4761),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4760),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4749),
.Y(n_4790)
);

NOR3xp33_ASAP7_75t_L g4791 ( 
.A(n_4748),
.B(n_3824),
.C(n_3337),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4754),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4755),
.Y(n_4793)
);

AOI22xp5_ASAP7_75t_L g4794 ( 
.A1(n_4737),
.A2(n_4042),
.B1(n_4044),
.B2(n_4026),
.Y(n_4794)
);

AOI21xp5_ASAP7_75t_L g4795 ( 
.A1(n_4731),
.A2(n_3586),
.B(n_3839),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4755),
.Y(n_4796)
);

BUFx2_ASAP7_75t_L g4797 ( 
.A(n_4741),
.Y(n_4797)
);

AOI221xp5_ASAP7_75t_L g4798 ( 
.A1(n_4734),
.A2(n_4751),
.B1(n_4746),
.B2(n_4759),
.C(n_4756),
.Y(n_4798)
);

AOI21xp33_ASAP7_75t_L g4799 ( 
.A1(n_4770),
.A2(n_611),
.B(n_612),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4762),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4776),
.Y(n_4801)
);

INVxp67_ASAP7_75t_L g4802 ( 
.A(n_4784),
.Y(n_4802)
);

INVx2_ASAP7_75t_L g4803 ( 
.A(n_4779),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4785),
.Y(n_4804)
);

AOI22xp33_ASAP7_75t_SL g4805 ( 
.A1(n_4775),
.A2(n_4730),
.B1(n_4729),
.B2(n_4764),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4778),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4797),
.B(n_4732),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4783),
.Y(n_4808)
);

NAND2x1_ASAP7_75t_L g4809 ( 
.A(n_4788),
.B(n_4766),
.Y(n_4809)
);

INVx2_ASAP7_75t_L g4810 ( 
.A(n_4781),
.Y(n_4810)
);

INVx2_ASAP7_75t_SL g4811 ( 
.A(n_4781),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4789),
.Y(n_4812)
);

OR2x2_ASAP7_75t_L g4813 ( 
.A(n_4774),
.B(n_4744),
.Y(n_4813)
);

NAND2xp5_ASAP7_75t_SL g4814 ( 
.A(n_4798),
.B(n_4739),
.Y(n_4814)
);

BUFx3_ASAP7_75t_L g4815 ( 
.A(n_4800),
.Y(n_4815)
);

AOI22xp5_ASAP7_75t_L g4816 ( 
.A1(n_4782),
.A2(n_4772),
.B1(n_4769),
.B2(n_4733),
.Y(n_4816)
);

NAND2xp5_ASAP7_75t_L g4817 ( 
.A(n_4773),
.B(n_4747),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4780),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4790),
.Y(n_4819)
);

NAND2xp5_ASAP7_75t_L g4820 ( 
.A(n_4799),
.B(n_4791),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4792),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4796),
.Y(n_4822)
);

AOI22xp5_ASAP7_75t_L g4823 ( 
.A1(n_4793),
.A2(n_4767),
.B1(n_4745),
.B2(n_4757),
.Y(n_4823)
);

INVx1_ASAP7_75t_SL g4824 ( 
.A(n_4794),
.Y(n_4824)
);

INVx2_ASAP7_75t_L g4825 ( 
.A(n_4786),
.Y(n_4825)
);

OAI21xp5_ASAP7_75t_SL g4826 ( 
.A1(n_4795),
.A2(n_4763),
.B(n_4758),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4777),
.B(n_4723),
.Y(n_4827)
);

OR2x6_ASAP7_75t_L g4828 ( 
.A(n_4787),
.B(n_4767),
.Y(n_4828)
);

AO21x1_ASAP7_75t_L g4829 ( 
.A1(n_4775),
.A2(n_4771),
.B(n_4054),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_4797),
.B(n_611),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_L g4831 ( 
.A(n_4775),
.B(n_611),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4785),
.Y(n_4832)
);

INVx2_ASAP7_75t_L g4833 ( 
.A(n_4779),
.Y(n_4833)
);

OAI21xp33_ASAP7_75t_L g4834 ( 
.A1(n_4775),
.A2(n_4045),
.B(n_3960),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_4775),
.B(n_612),
.Y(n_4835)
);

NAND2x1_ASAP7_75t_L g4836 ( 
.A(n_4797),
.B(n_3612),
.Y(n_4836)
);

NOR2xp33_ASAP7_75t_L g4837 ( 
.A(n_4818),
.B(n_612),
.Y(n_4837)
);

AND2x2_ASAP7_75t_L g4838 ( 
.A(n_4807),
.B(n_613),
.Y(n_4838)
);

INVx1_ASAP7_75t_SL g4839 ( 
.A(n_4830),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4801),
.B(n_613),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4801),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4803),
.Y(n_4842)
);

AOI22xp33_ASAP7_75t_L g4843 ( 
.A1(n_4833),
.A2(n_4825),
.B1(n_4824),
.B2(n_4804),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4832),
.Y(n_4844)
);

OAI22xp33_ASAP7_75t_L g4845 ( 
.A1(n_4811),
.A2(n_3633),
.B1(n_3653),
.B2(n_3612),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4815),
.Y(n_4846)
);

OAI221xp5_ASAP7_75t_L g4847 ( 
.A1(n_4805),
.A2(n_616),
.B1(n_614),
.B2(n_615),
.C(n_617),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4810),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4802),
.B(n_615),
.Y(n_4849)
);

OAI31xp33_ASAP7_75t_L g4850 ( 
.A1(n_4820),
.A2(n_619),
.A3(n_616),
.B(n_618),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_SL g4851 ( 
.A(n_4812),
.B(n_3633),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4831),
.Y(n_4852)
);

OAI221xp5_ASAP7_75t_L g4853 ( 
.A1(n_4826),
.A2(n_620),
.B1(n_616),
.B2(n_618),
.C(n_621),
.Y(n_4853)
);

OAI21xp33_ASAP7_75t_SL g4854 ( 
.A1(n_4814),
.A2(n_3964),
.B(n_3959),
.Y(n_4854)
);

AND2x2_ASAP7_75t_L g4855 ( 
.A(n_4806),
.B(n_618),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4835),
.B(n_4817),
.Y(n_4856)
);

AOI222xp33_ASAP7_75t_L g4857 ( 
.A1(n_4808),
.A2(n_3863),
.B1(n_622),
.B2(n_624),
.C1(n_620),
.C2(n_621),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4809),
.Y(n_4858)
);

AOI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4827),
.A2(n_3833),
.B(n_3832),
.Y(n_4859)
);

BUFx8_ASAP7_75t_SL g4860 ( 
.A(n_4828),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4816),
.B(n_620),
.Y(n_4861)
);

INVxp33_ASAP7_75t_L g4862 ( 
.A(n_4813),
.Y(n_4862)
);

AOI22xp5_ASAP7_75t_L g4863 ( 
.A1(n_4829),
.A2(n_3825),
.B1(n_3660),
.B2(n_3680),
.Y(n_4863)
);

INVxp67_ASAP7_75t_SL g4864 ( 
.A(n_4819),
.Y(n_4864)
);

INVx1_ASAP7_75t_SL g4865 ( 
.A(n_4821),
.Y(n_4865)
);

OAI322xp33_ASAP7_75t_L g4866 ( 
.A1(n_4822),
.A2(n_628),
.A3(n_627),
.B1(n_625),
.B2(n_623),
.C1(n_624),
.C2(n_626),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4834),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_SL g4868 ( 
.A(n_4823),
.B(n_3653),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4828),
.B(n_4836),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4830),
.Y(n_4870)
);

INVx2_ASAP7_75t_L g4871 ( 
.A(n_4803),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4838),
.B(n_623),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_4837),
.B(n_625),
.Y(n_4873)
);

OAI221xp5_ASAP7_75t_L g4874 ( 
.A1(n_4853),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.C(n_628),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4843),
.B(n_629),
.Y(n_4875)
);

BUFx12f_ASAP7_75t_L g4876 ( 
.A(n_4849),
.Y(n_4876)
);

NOR2xp33_ASAP7_75t_L g4877 ( 
.A(n_4860),
.B(n_4862),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4871),
.Y(n_4878)
);

NAND4xp25_ASAP7_75t_L g4879 ( 
.A(n_4856),
.B(n_631),
.C(n_629),
.D(n_630),
.Y(n_4879)
);

NOR2xp33_ASAP7_75t_L g4880 ( 
.A(n_4847),
.B(n_629),
.Y(n_4880)
);

OAI22xp33_ASAP7_75t_L g4881 ( 
.A1(n_4869),
.A2(n_4846),
.B1(n_4839),
.B2(n_4842),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_L g4882 ( 
.A(n_4839),
.B(n_630),
.Y(n_4882)
);

NOR3xp33_ASAP7_75t_L g4883 ( 
.A(n_4866),
.B(n_631),
.C(n_632),
.Y(n_4883)
);

NAND4xp25_ASAP7_75t_L g4884 ( 
.A(n_4848),
.B(n_634),
.C(n_632),
.D(n_633),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_SL g4885 ( 
.A(n_4858),
.B(n_3660),
.Y(n_4885)
);

NOR2x1_ASAP7_75t_L g4886 ( 
.A(n_4840),
.B(n_632),
.Y(n_4886)
);

AND2x2_ASAP7_75t_L g4887 ( 
.A(n_4861),
.B(n_633),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_L g4888 ( 
.A(n_4850),
.B(n_634),
.Y(n_4888)
);

NOR2xp33_ASAP7_75t_L g4889 ( 
.A(n_4870),
.B(n_635),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4841),
.Y(n_4890)
);

NAND3xp33_ASAP7_75t_L g4891 ( 
.A(n_4844),
.B(n_635),
.C(n_636),
.Y(n_4891)
);

AOI21xp33_ASAP7_75t_SL g4892 ( 
.A1(n_4867),
.A2(n_4852),
.B(n_4855),
.Y(n_4892)
);

AND2x2_ASAP7_75t_L g4893 ( 
.A(n_4864),
.B(n_636),
.Y(n_4893)
);

OAI211xp5_ASAP7_75t_L g4894 ( 
.A1(n_4865),
.A2(n_638),
.B(n_636),
.C(n_637),
.Y(n_4894)
);

NOR3xp33_ASAP7_75t_L g4895 ( 
.A(n_4854),
.B(n_4865),
.C(n_4845),
.Y(n_4895)
);

AND4x1_ASAP7_75t_L g4896 ( 
.A(n_4857),
.B(n_639),
.C(n_637),
.D(n_638),
.Y(n_4896)
);

AOI22xp5_ASAP7_75t_L g4897 ( 
.A1(n_4868),
.A2(n_3680),
.B1(n_3725),
.B2(n_3660),
.Y(n_4897)
);

AOI322xp5_ASAP7_75t_L g4898 ( 
.A1(n_4851),
.A2(n_3967),
.A3(n_3663),
.B1(n_644),
.B2(n_641),
.C1(n_643),
.C2(n_639),
.Y(n_4898)
);

INVx2_ASAP7_75t_L g4899 ( 
.A(n_4863),
.Y(n_4899)
);

O2A1O1Ixp33_ASAP7_75t_SL g4900 ( 
.A1(n_4859),
.A2(n_642),
.B(n_640),
.C(n_641),
.Y(n_4900)
);

OAI211xp5_ASAP7_75t_SL g4901 ( 
.A1(n_4843),
.A2(n_643),
.B(n_640),
.C(n_642),
.Y(n_4901)
);

OAI21xp33_ASAP7_75t_SL g4902 ( 
.A1(n_4843),
.A2(n_640),
.B(n_642),
.Y(n_4902)
);

NAND2xp5_ASAP7_75t_L g4903 ( 
.A(n_4838),
.B(n_643),
.Y(n_4903)
);

NOR2xp33_ASAP7_75t_L g4904 ( 
.A(n_4860),
.B(n_644),
.Y(n_4904)
);

NOR3xp33_ASAP7_75t_L g4905 ( 
.A(n_4853),
.B(n_644),
.C(n_645),
.Y(n_4905)
);

AOI222xp33_ASAP7_75t_L g4906 ( 
.A1(n_4837),
.A2(n_647),
.B1(n_649),
.B2(n_645),
.C1(n_646),
.C2(n_648),
.Y(n_4906)
);

AND2x2_ASAP7_75t_L g4907 ( 
.A(n_4838),
.B(n_646),
.Y(n_4907)
);

OAI22xp5_ASAP7_75t_L g4908 ( 
.A1(n_4843),
.A2(n_3725),
.B1(n_3732),
.B2(n_3680),
.Y(n_4908)
);

NAND4xp25_ASAP7_75t_SL g4909 ( 
.A(n_4843),
.B(n_649),
.C(n_647),
.D(n_648),
.Y(n_4909)
);

AOI321xp33_ASAP7_75t_L g4910 ( 
.A1(n_4877),
.A2(n_649),
.A3(n_651),
.B1(n_647),
.B2(n_648),
.C(n_650),
.Y(n_4910)
);

AOI221xp5_ASAP7_75t_L g4911 ( 
.A1(n_4881),
.A2(n_652),
.B1(n_650),
.B2(n_651),
.C(n_653),
.Y(n_4911)
);

XOR2xp5_ASAP7_75t_L g4912 ( 
.A(n_4909),
.B(n_650),
.Y(n_4912)
);

AOI221xp5_ASAP7_75t_L g4913 ( 
.A1(n_4902),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.C(n_655),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_4904),
.B(n_652),
.Y(n_4914)
);

AOI221xp5_ASAP7_75t_L g4915 ( 
.A1(n_4892),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.C(n_656),
.Y(n_4915)
);

AOI221xp5_ASAP7_75t_L g4916 ( 
.A1(n_4883),
.A2(n_657),
.B1(n_655),
.B2(n_656),
.C(n_658),
.Y(n_4916)
);

AOI211x1_ASAP7_75t_SL g4917 ( 
.A1(n_4901),
.A2(n_659),
.B(n_657),
.C(n_658),
.Y(n_4917)
);

AOI21xp5_ASAP7_75t_L g4918 ( 
.A1(n_4875),
.A2(n_658),
.B(n_659),
.Y(n_4918)
);

AOI321xp33_ASAP7_75t_L g4919 ( 
.A1(n_4878),
.A2(n_662),
.A3(n_664),
.B1(n_660),
.B2(n_661),
.C(n_663),
.Y(n_4919)
);

AOI22xp5_ASAP7_75t_L g4920 ( 
.A1(n_4905),
.A2(n_4880),
.B1(n_4887),
.B2(n_4879),
.Y(n_4920)
);

O2A1O1Ixp33_ASAP7_75t_L g4921 ( 
.A1(n_4882),
.A2(n_662),
.B(n_660),
.C(n_661),
.Y(n_4921)
);

AOI21xp5_ASAP7_75t_L g4922 ( 
.A1(n_4888),
.A2(n_662),
.B(n_663),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4907),
.Y(n_4923)
);

AOI21xp33_ASAP7_75t_SL g4924 ( 
.A1(n_4891),
.A2(n_663),
.B(n_664),
.Y(n_4924)
);

OAI21xp33_ASAP7_75t_L g4925 ( 
.A1(n_4889),
.A2(n_664),
.B(n_665),
.Y(n_4925)
);

NOR4xp75_ASAP7_75t_L g4926 ( 
.A(n_4874),
.B(n_667),
.C(n_665),
.D(n_666),
.Y(n_4926)
);

AOI221x1_ASAP7_75t_L g4927 ( 
.A1(n_4890),
.A2(n_668),
.B1(n_665),
.B2(n_666),
.C(n_704),
.Y(n_4927)
);

AOI22xp33_ASAP7_75t_L g4928 ( 
.A1(n_4876),
.A2(n_3732),
.B1(n_3725),
.B2(n_666),
.Y(n_4928)
);

AOI221xp5_ASAP7_75t_L g4929 ( 
.A1(n_4900),
.A2(n_4895),
.B1(n_4893),
.B2(n_4884),
.C(n_4894),
.Y(n_4929)
);

O2A1O1Ixp33_ASAP7_75t_L g4930 ( 
.A1(n_4873),
.A2(n_668),
.B(n_706),
.C(n_705),
.Y(n_4930)
);

INVxp67_ASAP7_75t_L g4931 ( 
.A(n_4872),
.Y(n_4931)
);

AOI21xp5_ASAP7_75t_L g4932 ( 
.A1(n_4903),
.A2(n_705),
.B(n_708),
.Y(n_4932)
);

NAND4xp25_ASAP7_75t_SL g4933 ( 
.A(n_4906),
.B(n_710),
.C(n_708),
.D(n_709),
.Y(n_4933)
);

AOI221xp5_ASAP7_75t_L g4934 ( 
.A1(n_4916),
.A2(n_4884),
.B1(n_4885),
.B2(n_4899),
.C(n_4908),
.Y(n_4934)
);

CKINVDCx5p33_ASAP7_75t_R g4935 ( 
.A(n_4914),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4913),
.B(n_4896),
.Y(n_4936)
);

INVxp67_ASAP7_75t_L g4937 ( 
.A(n_4912),
.Y(n_4937)
);

AOI322xp5_ASAP7_75t_L g4938 ( 
.A1(n_4929),
.A2(n_4886),
.A3(n_4897),
.B1(n_4898),
.B2(n_3663),
.C1(n_715),
.C2(n_718),
.Y(n_4938)
);

AOI21xp5_ASAP7_75t_L g4939 ( 
.A1(n_4932),
.A2(n_711),
.B(n_714),
.Y(n_4939)
);

AOI31xp33_ASAP7_75t_L g4940 ( 
.A1(n_4911),
.A2(n_717),
.A3(n_711),
.B(n_716),
.Y(n_4940)
);

OAI211xp5_ASAP7_75t_L g4941 ( 
.A1(n_4915),
.A2(n_720),
.B(n_718),
.C(n_719),
.Y(n_4941)
);

BUFx6f_ASAP7_75t_L g4942 ( 
.A(n_4923),
.Y(n_4942)
);

AO22x2_ASAP7_75t_L g4943 ( 
.A1(n_4922),
.A2(n_721),
.B1(n_719),
.B2(n_720),
.Y(n_4943)
);

AOI322xp5_ASAP7_75t_L g4944 ( 
.A1(n_4920),
.A2(n_4931),
.A3(n_4925),
.B1(n_4928),
.B2(n_4917),
.C1(n_4910),
.C2(n_4926),
.Y(n_4944)
);

AOI221xp5_ASAP7_75t_L g4945 ( 
.A1(n_4933),
.A2(n_3732),
.B1(n_723),
.B2(n_721),
.C(n_722),
.Y(n_4945)
);

AOI22xp33_ASAP7_75t_L g4946 ( 
.A1(n_4918),
.A2(n_725),
.B1(n_723),
.B2(n_724),
.Y(n_4946)
);

AOI222xp33_ASAP7_75t_L g4947 ( 
.A1(n_4919),
.A2(n_728),
.B1(n_730),
.B2(n_724),
.C1(n_727),
.C2(n_729),
.Y(n_4947)
);

NAND4xp25_ASAP7_75t_L g4948 ( 
.A(n_4921),
.B(n_730),
.C(n_728),
.D(n_729),
.Y(n_4948)
);

NAND3xp33_ASAP7_75t_SL g4949 ( 
.A(n_4930),
.B(n_731),
.C(n_732),
.Y(n_4949)
);

AOI22xp5_ASAP7_75t_L g4950 ( 
.A1(n_4924),
.A2(n_3663),
.B1(n_734),
.B2(n_732),
.Y(n_4950)
);

OAI22xp33_ASAP7_75t_SL g4951 ( 
.A1(n_4927),
.A2(n_735),
.B1(n_733),
.B2(n_734),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_4916),
.B(n_733),
.Y(n_4952)
);

OAI221xp5_ASAP7_75t_L g4953 ( 
.A1(n_4910),
.A2(n_737),
.B1(n_735),
.B2(n_736),
.C(n_738),
.Y(n_4953)
);

XNOR2x1_ASAP7_75t_L g4954 ( 
.A(n_4926),
.B(n_736),
.Y(n_4954)
);

NOR2xp33_ASAP7_75t_L g4955 ( 
.A(n_4912),
.B(n_737),
.Y(n_4955)
);

AOI322xp5_ASAP7_75t_L g4956 ( 
.A1(n_4929),
.A2(n_738),
.A3(n_739),
.B1(n_740),
.B2(n_741),
.C1(n_742),
.C2(n_743),
.Y(n_4956)
);

OAI211xp5_ASAP7_75t_SL g4957 ( 
.A1(n_4929),
.A2(n_742),
.B(n_739),
.C(n_740),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4943),
.Y(n_4958)
);

NAND4xp75_ASAP7_75t_L g4959 ( 
.A(n_4945),
.B(n_745),
.C(n_743),
.D(n_744),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4954),
.Y(n_4960)
);

NAND4xp75_ASAP7_75t_L g4961 ( 
.A(n_4939),
.B(n_746),
.C(n_744),
.D(n_745),
.Y(n_4961)
);

NAND2xp5_ASAP7_75t_L g4962 ( 
.A(n_4956),
.B(n_746),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4936),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4952),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4955),
.Y(n_4965)
);

OR2x2_ASAP7_75t_L g4966 ( 
.A(n_4948),
.B(n_747),
.Y(n_4966)
);

XNOR2xp5_ASAP7_75t_L g4967 ( 
.A(n_4953),
.B(n_748),
.Y(n_4967)
);

AND2x4_ASAP7_75t_L g4968 ( 
.A(n_4942),
.B(n_748),
.Y(n_4968)
);

INVx1_ASAP7_75t_SL g4969 ( 
.A(n_4942),
.Y(n_4969)
);

OAI211xp5_ASAP7_75t_L g4970 ( 
.A1(n_4947),
.A2(n_752),
.B(n_749),
.C(n_751),
.Y(n_4970)
);

NOR2xp33_ASAP7_75t_L g4971 ( 
.A(n_4937),
.B(n_751),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4951),
.Y(n_4972)
);

NOR2xp33_ASAP7_75t_L g4973 ( 
.A(n_4957),
.B(n_752),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4968),
.Y(n_4974)
);

AOI322xp5_ASAP7_75t_L g4975 ( 
.A1(n_4969),
.A2(n_4949),
.A3(n_4934),
.B1(n_4935),
.B2(n_4946),
.C1(n_4950),
.C2(n_4944),
.Y(n_4975)
);

OAI221xp5_ASAP7_75t_L g4976 ( 
.A1(n_4970),
.A2(n_4941),
.B1(n_4938),
.B2(n_4940),
.C(n_755),
.Y(n_4976)
);

AND2x2_ASAP7_75t_L g4977 ( 
.A(n_4972),
.B(n_753),
.Y(n_4977)
);

NAND3xp33_ASAP7_75t_L g4978 ( 
.A(n_4971),
.B(n_4967),
.C(n_4963),
.Y(n_4978)
);

OR3x2_ASAP7_75t_L g4979 ( 
.A(n_4966),
.B(n_754),
.C(n_756),
.Y(n_4979)
);

HB1xp67_ASAP7_75t_L g4980 ( 
.A(n_4968),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_SL g4981 ( 
.A(n_4962),
.B(n_754),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_4958),
.B(n_756),
.Y(n_4982)
);

NAND3xp33_ASAP7_75t_L g4983 ( 
.A(n_4960),
.B(n_757),
.C(n_758),
.Y(n_4983)
);

AOI222xp33_ASAP7_75t_L g4984 ( 
.A1(n_4973),
.A2(n_760),
.B1(n_762),
.B2(n_757),
.C1(n_759),
.C2(n_761),
.Y(n_4984)
);

AOI22xp5_ASAP7_75t_L g4985 ( 
.A1(n_4959),
.A2(n_4964),
.B1(n_4965),
.B2(n_4961),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4968),
.Y(n_4986)
);

OAI221xp5_ASAP7_75t_L g4987 ( 
.A1(n_4976),
.A2(n_4982),
.B1(n_4983),
.B2(n_4985),
.C(n_4978),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4977),
.B(n_939),
.Y(n_4988)
);

NOR2x1_ASAP7_75t_L g4989 ( 
.A(n_4981),
.B(n_759),
.Y(n_4989)
);

INVx1_ASAP7_75t_L g4990 ( 
.A(n_4980),
.Y(n_4990)
);

XOR2xp5_ASAP7_75t_L g4991 ( 
.A(n_4979),
.B(n_762),
.Y(n_4991)
);

AOI22xp5_ASAP7_75t_L g4992 ( 
.A1(n_4984),
.A2(n_766),
.B1(n_764),
.B2(n_765),
.Y(n_4992)
);

A2O1A1Ixp33_ASAP7_75t_L g4993 ( 
.A1(n_4975),
.A2(n_766),
.B(n_764),
.C(n_765),
.Y(n_4993)
);

AOI22xp5_ASAP7_75t_L g4994 ( 
.A1(n_4990),
.A2(n_4986),
.B1(n_4974),
.B2(n_770),
.Y(n_4994)
);

AOI22xp5_ASAP7_75t_L g4995 ( 
.A1(n_4991),
.A2(n_771),
.B1(n_767),
.B2(n_768),
.Y(n_4995)
);

AOI31xp33_ASAP7_75t_L g4996 ( 
.A1(n_4993),
.A2(n_772),
.A3(n_767),
.B(n_771),
.Y(n_4996)
);

OAI22x1_ASAP7_75t_L g4997 ( 
.A1(n_4992),
.A2(n_774),
.B1(n_772),
.B2(n_773),
.Y(n_4997)
);

CKINVDCx20_ASAP7_75t_R g4998 ( 
.A(n_4988),
.Y(n_4998)
);

OAI22x1_ASAP7_75t_L g4999 ( 
.A1(n_4989),
.A2(n_776),
.B1(n_773),
.B2(n_774),
.Y(n_4999)
);

BUFx2_ASAP7_75t_SL g5000 ( 
.A(n_4998),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4996),
.Y(n_5001)
);

NOR2x1_ASAP7_75t_L g5002 ( 
.A(n_4994),
.B(n_4987),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_5002),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_5000),
.B(n_4995),
.Y(n_5004)
);

AOI22xp5_ASAP7_75t_L g5005 ( 
.A1(n_5003),
.A2(n_5001),
.B1(n_5004),
.B2(n_4997),
.Y(n_5005)
);

OAI21xp5_ASAP7_75t_L g5006 ( 
.A1(n_5003),
.A2(n_4999),
.B(n_777),
.Y(n_5006)
);

AOI22xp33_ASAP7_75t_SL g5007 ( 
.A1(n_5006),
.A2(n_781),
.B1(n_778),
.B2(n_780),
.Y(n_5007)
);

AOI21xp5_ASAP7_75t_L g5008 ( 
.A1(n_5005),
.A2(n_783),
.B(n_784),
.Y(n_5008)
);

NOR2x2_ASAP7_75t_L g5009 ( 
.A(n_5007),
.B(n_783),
.Y(n_5009)
);

OA21x2_ASAP7_75t_L g5010 ( 
.A1(n_5008),
.A2(n_784),
.B(n_785),
.Y(n_5010)
);

AOI22xp5_ASAP7_75t_SL g5011 ( 
.A1(n_5010),
.A2(n_788),
.B1(n_786),
.B2(n_787),
.Y(n_5011)
);

AOI22x1_ASAP7_75t_L g5012 ( 
.A1(n_5009),
.A2(n_789),
.B1(n_786),
.B2(n_787),
.Y(n_5012)
);

OAI221xp5_ASAP7_75t_L g5013 ( 
.A1(n_5011),
.A2(n_793),
.B1(n_791),
.B2(n_792),
.C(n_794),
.Y(n_5013)
);

AOI211xp5_ASAP7_75t_L g5014 ( 
.A1(n_5013),
.A2(n_5012),
.B(n_796),
.C(n_795),
.Y(n_5014)
);


endmodule