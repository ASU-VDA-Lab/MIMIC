module fake_aes_107_n_1646 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_381, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_379, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_380, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1646);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_381;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_379;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_380;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1646;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_1627;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1618;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_1619;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_1631;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_1620;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_1623;
wire n_556;
wire n_1214;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_1613;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1582;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_1639;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_994;
wire n_930;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_510;
wire n_1075;
wire n_1615;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1628;
wire n_1533;
wire n_1611;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_1563;
wire n_1642;
wire n_824;
wire n_793;
wire n_753;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1602;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1361;
wire n_1333;
wire n_1557;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1625;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_1629;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_1643;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1608;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_1593;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_1621;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_1638;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1645;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_1633;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1626;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1641;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_1583;
wire n_606;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_1634;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_659;
wire n_432;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1460;
wire n_1372;
wire n_1640;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_1635;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1576;
wire n_1609;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1610;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_1622;
wire n_1614;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1612;
wire n_1636;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1130;
wire n_584;
wire n_1042;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_1624;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1616;
wire n_1378;
wire n_1570;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_401;
wire n_481;
wire n_443;
wire n_694;
wire n_1601;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1644;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_1630;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1637;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1617;
wire n_1632;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_1607;
wire n_906;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_600;
wire n_1531;
wire n_1548;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
CKINVDCx16_ASAP7_75t_R g382 ( .A(n_239), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_333), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_81), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_46), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_199), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_201), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_287), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_43), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_219), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_274), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_186), .Y(n_392) );
NOR2xp67_ASAP7_75t_L g393 ( .A(n_215), .B(n_148), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_292), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_212), .Y(n_395) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_327), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_180), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_224), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_131), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_57), .Y(n_400) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_300), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_159), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_31), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_137), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_273), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_118), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_52), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_375), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_92), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_307), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_240), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_146), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_268), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_60), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_253), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_95), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_255), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_291), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_230), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_211), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_100), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_338), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_206), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_26), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_313), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_351), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_209), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_39), .Y(n_428) );
INVx2_ASAP7_75t_SL g429 ( .A(n_138), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_288), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_277), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_228), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_266), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_158), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g435 ( .A(n_111), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g436 ( .A(n_376), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_39), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_205), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_297), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_129), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_139), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_128), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_82), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_147), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_29), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_285), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_249), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_17), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_173), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_329), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_276), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_373), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_130), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_135), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_167), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_257), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_145), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_81), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_59), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_223), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_11), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_9), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_187), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_82), .Y(n_464) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_203), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_86), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_55), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_190), .Y(n_468) );
BUFx3_ASAP7_75t_L g469 ( .A(n_58), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_55), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_310), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_176), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_368), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_189), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_2), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_171), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_43), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_192), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_197), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_340), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_62), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_5), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_78), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_86), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_62), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_232), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_283), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_33), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_335), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_357), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_120), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_346), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_14), .Y(n_493) );
BUFx10_ASAP7_75t_L g494 ( .A(n_378), .Y(n_494) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_73), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_251), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_302), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_262), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_80), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_244), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_325), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_69), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_143), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_52), .Y(n_504) );
CKINVDCx14_ASAP7_75t_R g505 ( .A(n_272), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_108), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_301), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_352), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_30), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_37), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_365), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_341), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_77), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_160), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_207), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_299), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_104), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_204), .Y(n_518) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_331), .Y(n_519) );
INVxp33_ASAP7_75t_L g520 ( .A(n_349), .Y(n_520) );
INVxp33_ASAP7_75t_L g521 ( .A(n_229), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_367), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_132), .Y(n_523) );
INVxp67_ASAP7_75t_SL g524 ( .A(n_140), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_242), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_57), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_354), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_366), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_116), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_194), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_36), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_217), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_269), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_144), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_2), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_164), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_183), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_348), .Y(n_538) );
CKINVDCx16_ASAP7_75t_R g539 ( .A(n_58), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_225), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_381), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_265), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_170), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_4), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_20), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_151), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_31), .Y(n_547) );
INVxp33_ASAP7_75t_L g548 ( .A(n_35), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_121), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_214), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_172), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_250), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_353), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_90), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_185), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_8), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_289), .Y(n_557) );
NOR2xp67_ASAP7_75t_L g558 ( .A(n_70), .B(n_56), .Y(n_558) );
BUFx3_ASAP7_75t_L g559 ( .A(n_179), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_256), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_22), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_108), .Y(n_562) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_45), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_169), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_308), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_296), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_320), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_317), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_28), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_67), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_12), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_48), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_494), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_459), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_401), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_494), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_401), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_401), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_429), .B(n_0), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_444), .B(n_0), .Y(n_580) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_401), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_459), .Y(n_582) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_419), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_422), .B(n_1), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_460), .B(n_1), .Y(n_585) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_419), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_419), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_419), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_462), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_420), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_416), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_420), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_520), .B(n_3), .Y(n_593) );
INVx6_ASAP7_75t_L g594 ( .A(n_494), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_462), .Y(n_595) );
BUFx2_ASAP7_75t_L g596 ( .A(n_421), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_548), .B(n_3), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_435), .A2(n_458), .B1(n_539), .B2(n_517), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_389), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_424), .Y(n_600) );
INVx6_ASAP7_75t_L g601 ( .A(n_559), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_464), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_420), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_548), .B(n_4), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_443), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_389), .B(n_5), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_464), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_469), .B(n_6), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_384), .B(n_6), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_484), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_382), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_481), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_420), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_469), .B(n_7), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_481), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_573), .B(n_502), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_575), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_599), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_573), .B(n_576), .Y(n_619) );
CKINVDCx14_ASAP7_75t_R g620 ( .A(n_611), .Y(n_620) );
NOR2x1p5_ASAP7_75t_L g621 ( .A(n_573), .B(n_576), .Y(n_621) );
INVx3_ASAP7_75t_L g622 ( .A(n_606), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_599), .Y(n_623) );
OR2x6_ASAP7_75t_L g624 ( .A(n_597), .B(n_558), .Y(n_624) );
INVxp67_ASAP7_75t_L g625 ( .A(n_610), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_596), .B(n_520), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_594), .B(n_521), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_594), .B(n_521), .Y(n_628) );
AND2x6_ASAP7_75t_L g629 ( .A(n_606), .B(n_559), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_599), .Y(n_630) );
BUFx3_ASAP7_75t_L g631 ( .A(n_601), .Y(n_631) );
NAND2x1p5_ASAP7_75t_L g632 ( .A(n_606), .B(n_383), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_606), .Y(n_633) );
INVx4_ASAP7_75t_L g634 ( .A(n_608), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_599), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_575), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_596), .B(n_505), .Y(n_637) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_581), .Y(n_638) );
CKINVDCx11_ASAP7_75t_R g639 ( .A(n_608), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_594), .B(n_390), .Y(n_640) );
INVx4_ASAP7_75t_L g641 ( .A(n_608), .Y(n_641) );
BUFx3_ASAP7_75t_L g642 ( .A(n_601), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_608), .Y(n_643) );
NAND2xp33_ASAP7_75t_L g644 ( .A(n_573), .B(n_426), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_614), .Y(n_645) );
AND2x6_ASAP7_75t_L g646 ( .A(n_614), .B(n_386), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_575), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_576), .B(n_436), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_576), .B(n_502), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_614), .B(n_478), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_591), .Y(n_651) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_581), .Y(n_652) );
INVx4_ASAP7_75t_L g653 ( .A(n_614), .Y(n_653) );
INVx4_ASAP7_75t_L g654 ( .A(n_601), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_594), .B(n_480), .Y(n_655) );
INVx3_ASAP7_75t_L g656 ( .A(n_601), .Y(n_656) );
INVx8_ASAP7_75t_L g657 ( .A(n_594), .Y(n_657) );
CKINVDCx16_ASAP7_75t_R g658 ( .A(n_598), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_577), .Y(n_659) );
INVx4_ASAP7_75t_L g660 ( .A(n_601), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_577), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_621), .B(n_597), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_627), .B(n_605), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_634), .B(n_580), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_634), .B(n_580), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_621), .B(n_604), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_616), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_628), .B(n_600), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_651), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_620), .Y(n_670) );
INVxp67_ASAP7_75t_L g671 ( .A(n_637), .Y(n_671) );
BUFx8_ASAP7_75t_L g672 ( .A(n_626), .Y(n_672) );
NAND2x1p5_ASAP7_75t_L g673 ( .A(n_634), .B(n_385), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_616), .Y(n_674) );
INVx3_ASAP7_75t_L g675 ( .A(n_634), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_639), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_616), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_637), .B(n_593), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_626), .B(n_598), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_641), .B(n_388), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_649), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_649), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_641), .B(n_391), .Y(n_683) );
NAND3xp33_ASAP7_75t_SL g684 ( .A(n_625), .B(n_404), .C(n_402), .Y(n_684) );
INVx2_ASAP7_75t_SL g685 ( .A(n_648), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_640), .B(n_604), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_655), .B(n_579), .Y(n_687) );
OR2x2_ASAP7_75t_SL g688 ( .A(n_658), .B(n_569), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_632), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_649), .B(n_584), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_632), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_649), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_641), .B(n_585), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_624), .B(n_609), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_618), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_653), .B(n_387), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_650), .B(n_609), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_618), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_646), .A2(n_402), .B1(n_441), .B2(n_404), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_653), .B(n_392), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_623), .Y(n_701) );
INVx4_ASAP7_75t_L g702 ( .A(n_657), .Y(n_702) );
BUFx3_ASAP7_75t_L g703 ( .A(n_657), .Y(n_703) );
BUFx2_ASAP7_75t_L g704 ( .A(n_629), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_623), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_646), .A2(n_442), .B1(n_449), .B2(n_441), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_653), .B(n_657), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_630), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_619), .A2(n_445), .B(n_499), .C(n_484), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_630), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_653), .B(n_394), .Y(n_711) );
AND2x4_ASAP7_75t_L g712 ( .A(n_624), .B(n_442), .Y(n_712) );
INVx3_ASAP7_75t_L g713 ( .A(n_622), .Y(n_713) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_646), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_632), .Y(n_715) );
INVx1_ASAP7_75t_SL g716 ( .A(n_629), .Y(n_716) );
INVx4_ASAP7_75t_L g717 ( .A(n_657), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_657), .B(n_394), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_646), .B(n_399), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_635), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_646), .B(n_399), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_635), .Y(n_722) );
CKINVDCx6p67_ASAP7_75t_R g723 ( .A(n_624), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_631), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_643), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_643), .B(n_395), .Y(n_726) );
O2A1O1Ixp33_ASAP7_75t_L g727 ( .A1(n_645), .A2(n_582), .B(n_589), .C(n_574), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_646), .B(n_410), .Y(n_728) );
NAND3xp33_ASAP7_75t_SL g729 ( .A(n_645), .B(n_457), .C(n_449), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_622), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g731 ( .A1(n_622), .A2(n_582), .B(n_589), .C(n_574), .Y(n_731) );
BUFx3_ASAP7_75t_L g732 ( .A(n_642), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_617), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_617), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_622), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_624), .B(n_535), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_646), .A2(n_602), .B1(n_607), .B2(n_595), .Y(n_737) );
INVxp67_ASAP7_75t_L g738 ( .A(n_624), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_633), .B(n_595), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_633), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_633), .B(n_397), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_629), .B(n_410), .Y(n_742) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_633), .A2(n_569), .B1(n_486), .B2(n_487), .Y(n_743) );
NOR2xp33_ASAP7_75t_R g744 ( .A(n_629), .B(n_457), .Y(n_744) );
AOI211xp5_ASAP7_75t_L g745 ( .A1(n_644), .A2(n_545), .B(n_554), .C(n_535), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_636), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g747 ( .A1(n_659), .A2(n_607), .B(n_612), .C(n_602), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_629), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_656), .B(n_545), .Y(n_749) );
AND2x4_ASAP7_75t_L g750 ( .A(n_629), .B(n_486), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_713), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_730), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_713), .Y(n_753) );
BUFx6f_ASAP7_75t_L g754 ( .A(n_714), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_735), .Y(n_755) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_714), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_662), .B(n_629), .Y(n_757) );
NOR2xp67_ASAP7_75t_L g758 ( .A(n_669), .B(n_554), .Y(n_758) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_714), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_694), .A2(n_505), .B1(n_497), .B2(n_487), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_667), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_669), .B(n_497), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_691), .A2(n_540), .B1(n_538), .B2(n_571), .Y(n_763) );
INVx3_ASAP7_75t_L g764 ( .A(n_675), .Y(n_764) );
INVx3_ASAP7_75t_L g765 ( .A(n_675), .Y(n_765) );
INVx1_ASAP7_75t_SL g766 ( .A(n_749), .Y(n_766) );
AO21x1_ASAP7_75t_L g767 ( .A1(n_739), .A2(n_405), .B(n_398), .Y(n_767) );
A2O1A1Ixp33_ASAP7_75t_L g768 ( .A1(n_697), .A2(n_403), .B(n_407), .C(n_400), .Y(n_768) );
BUFx3_ASAP7_75t_L g769 ( .A(n_672), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_750), .A2(n_538), .B1(n_540), .B2(n_571), .Y(n_770) );
BUFx12f_ASAP7_75t_L g771 ( .A(n_670), .Y(n_771) );
BUFx8_ASAP7_75t_L g772 ( .A(n_712), .Y(n_772) );
AND2x4_ASAP7_75t_L g773 ( .A(n_685), .B(n_495), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_676), .Y(n_774) );
AND2x4_ASAP7_75t_L g775 ( .A(n_691), .B(n_563), .Y(n_775) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_714), .Y(n_776) );
INVx3_ASAP7_75t_L g777 ( .A(n_702), .Y(n_777) );
INVx5_ASAP7_75t_L g778 ( .A(n_689), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_698), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_750), .A2(n_556), .B1(n_477), .B2(n_440), .Y(n_780) );
INVx3_ASAP7_75t_L g781 ( .A(n_702), .Y(n_781) );
BUFx6f_ASAP7_75t_SL g782 ( .A(n_712), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_674), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_698), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_L g785 ( .A1(n_697), .A2(n_414), .B(n_428), .C(n_409), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_740), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_677), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_705), .Y(n_788) );
AND2x4_ASAP7_75t_SL g789 ( .A(n_715), .B(n_654), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_705), .Y(n_790) );
XOR2x2_ASAP7_75t_SL g791 ( .A(n_699), .B(n_437), .Y(n_791) );
A2O1A1Ixp33_ASAP7_75t_L g792 ( .A1(n_725), .A2(n_461), .B(n_466), .C(n_448), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_671), .B(n_654), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_722), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_738), .B(n_654), .Y(n_795) );
AND2x4_ASAP7_75t_L g796 ( .A(n_715), .B(n_467), .Y(n_796) );
AOI222xp33_ASAP7_75t_L g797 ( .A1(n_679), .A2(n_615), .B1(n_612), .B2(n_475), .C1(n_482), .C2(n_485), .Y(n_797) );
O2A1O1Ixp33_ASAP7_75t_L g798 ( .A1(n_731), .A2(n_483), .B(n_488), .C(n_470), .Y(n_798) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_703), .Y(n_799) );
OAI22x1_ASAP7_75t_L g800 ( .A1(n_706), .A2(n_418), .B1(n_489), .B2(n_440), .Y(n_800) );
O2A1O1Ixp33_ASAP7_75t_L g801 ( .A1(n_731), .A2(n_504), .B(n_506), .C(n_493), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_662), .B(n_666), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_722), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_694), .A2(n_489), .B1(n_503), .B2(n_418), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_666), .B(n_654), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_681), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_673), .Y(n_807) );
A2O1A1Ixp33_ASAP7_75t_L g808 ( .A1(n_727), .A2(n_510), .B(n_526), .C(n_513), .Y(n_808) );
CKINVDCx6p67_ASAP7_75t_R g809 ( .A(n_723), .Y(n_809) );
A2O1A1Ixp33_ASAP7_75t_L g810 ( .A1(n_739), .A2(n_529), .B(n_544), .C(n_531), .Y(n_810) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_672), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_668), .B(n_660), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_736), .A2(n_522), .B1(n_523), .B2(n_503), .Y(n_813) );
INVx3_ASAP7_75t_L g814 ( .A(n_717), .Y(n_814) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_703), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_686), .B(n_663), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_664), .A2(n_660), .B(n_631), .Y(n_817) );
AOI21x1_ASAP7_75t_L g818 ( .A1(n_680), .A2(n_659), .B(n_647), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_682), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_695), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_673), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_737), .A2(n_522), .B1(n_525), .B2(n_523), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_692), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_701), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_678), .B(n_660), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_704), .A2(n_547), .B1(n_562), .B2(n_561), .Y(n_826) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_744), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_708), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_710), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_690), .B(n_525), .Y(n_830) );
A2O1A1Ixp33_ASAP7_75t_L g831 ( .A1(n_720), .A2(n_570), .B(n_656), .C(n_615), .Y(n_831) );
BUFx6f_ASAP7_75t_L g832 ( .A(n_717), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_724), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_743), .Y(n_834) );
INVx5_ASAP7_75t_L g835 ( .A(n_732), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_745), .B(n_532), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_744), .B(n_509), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_729), .A2(n_533), .B1(n_534), .B2(n_532), .Y(n_838) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_732), .Y(n_839) );
A2O1A1Ixp33_ASAP7_75t_L g840 ( .A1(n_747), .A2(n_656), .B(n_572), .C(n_509), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_737), .B(n_533), .Y(n_841) );
O2A1O1Ixp33_ASAP7_75t_SL g842 ( .A1(n_747), .A2(n_408), .B(n_412), .C(n_406), .Y(n_842) );
INVxp33_ASAP7_75t_SL g843 ( .A(n_748), .Y(n_843) );
BUFx3_ASAP7_75t_L g844 ( .A(n_688), .Y(n_844) );
OR2x2_ASAP7_75t_L g845 ( .A(n_684), .B(n_572), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_665), .Y(n_846) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_707), .Y(n_847) );
A2O1A1Ixp33_ASAP7_75t_L g848 ( .A1(n_693), .A2(n_656), .B(n_415), .C(n_417), .Y(n_848) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_733), .Y(n_849) );
OAI21x1_ASAP7_75t_L g850 ( .A1(n_741), .A2(n_450), .B(n_411), .Y(n_850) );
HAxp5_ASAP7_75t_L g851 ( .A(n_709), .B(n_7), .CON(n_851), .SN(n_851) );
NOR2xp67_ASAP7_75t_SL g852 ( .A(n_742), .B(n_534), .Y(n_852) );
INVx3_ASAP7_75t_L g853 ( .A(n_716), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_665), .Y(n_854) );
OR2x6_ASAP7_75t_L g855 ( .A(n_680), .B(n_393), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_726), .Y(n_856) );
BUFx6f_ASAP7_75t_L g857 ( .A(n_733), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_696), .B(n_536), .Y(n_858) );
BUFx12f_ASAP7_75t_L g859 ( .A(n_741), .Y(n_859) );
INVx4_ASAP7_75t_L g860 ( .A(n_746), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_734), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_726), .Y(n_862) );
AND2x4_ASAP7_75t_L g863 ( .A(n_683), .B(n_642), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_683), .A2(n_423), .B1(n_425), .B2(n_413), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_687), .A2(n_542), .B1(n_536), .B2(n_465), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_734), .Y(n_866) );
BUFx6f_ASAP7_75t_L g867 ( .A(n_746), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_711), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_700), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_700), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_719), .Y(n_871) );
INVx1_ASAP7_75t_SL g872 ( .A(n_721), .Y(n_872) );
AOI21xp5_ASAP7_75t_L g873 ( .A1(n_728), .A2(n_519), .B(n_396), .Y(n_873) );
INVxp67_ASAP7_75t_L g874 ( .A(n_718), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_713), .Y(n_875) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_669), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_750), .A2(n_542), .B1(n_524), .B2(n_427), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_667), .Y(n_878) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_669), .Y(n_879) );
A2O1A1Ixp33_ASAP7_75t_L g880 ( .A1(n_697), .A2(n_430), .B(n_432), .C(n_431), .Y(n_880) );
BUFx12f_ASAP7_75t_L g881 ( .A(n_670), .Y(n_881) );
AND2x4_ASAP7_75t_L g882 ( .A(n_685), .B(n_553), .Y(n_882) );
OR2x6_ASAP7_75t_L g883 ( .A(n_743), .B(n_433), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_662), .B(n_555), .Y(n_884) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_714), .Y(n_885) );
AOI21xp5_ASAP7_75t_L g886 ( .A1(n_664), .A2(n_438), .B(n_434), .Y(n_886) );
BUFx12f_ASAP7_75t_L g887 ( .A(n_670), .Y(n_887) );
INVx4_ASAP7_75t_L g888 ( .A(n_714), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_730), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_691), .A2(n_439), .B1(n_447), .B2(n_446), .Y(n_890) );
INVx4_ASAP7_75t_L g891 ( .A(n_714), .Y(n_891) );
NOR2xp67_ASAP7_75t_L g892 ( .A(n_778), .B(n_119), .Y(n_892) );
OAI21x1_ASAP7_75t_L g893 ( .A1(n_850), .A2(n_818), .B(n_817), .Y(n_893) );
O2A1O1Ixp33_ASAP7_75t_L g894 ( .A1(n_768), .A2(n_453), .B(n_455), .C(n_451), .Y(n_894) );
INVx2_ASAP7_75t_SL g895 ( .A(n_769), .Y(n_895) );
NAND3xp33_ASAP7_75t_L g896 ( .A(n_880), .B(n_583), .C(n_581), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_860), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_860), .Y(n_898) );
AOI21x1_ASAP7_75t_L g899 ( .A1(n_767), .A2(n_472), .B(n_468), .Y(n_899) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_876), .Y(n_900) );
INVx2_ASAP7_75t_L g901 ( .A(n_779), .Y(n_901) );
OAI21x1_ASAP7_75t_L g902 ( .A1(n_820), .A2(n_472), .B(n_468), .Y(n_902) );
OAI21x1_ASAP7_75t_L g903 ( .A1(n_820), .A2(n_463), .B(n_456), .Y(n_903) );
O2A1O1Ixp5_ASAP7_75t_L g904 ( .A1(n_848), .A2(n_473), .B(n_474), .C(n_471), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_784), .Y(n_905) );
NAND2x1_ASAP7_75t_L g906 ( .A(n_832), .B(n_476), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_828), .A2(n_490), .B1(n_491), .B2(n_479), .Y(n_907) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_828), .A2(n_498), .B1(n_500), .B2(n_492), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_802), .A2(n_501), .B1(n_508), .B2(n_507), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_762), .B(n_496), .Y(n_910) );
OA21x2_ASAP7_75t_L g911 ( .A1(n_840), .A2(n_512), .B(n_511), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g912 ( .A1(n_763), .A2(n_454), .B1(n_452), .B2(n_565), .Y(n_912) );
OAI21x1_ASAP7_75t_L g913 ( .A1(n_788), .A2(n_515), .B(n_514), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_802), .A2(n_518), .B1(n_527), .B2(n_516), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_790), .Y(n_915) );
OAI21x1_ASAP7_75t_L g916 ( .A1(n_794), .A2(n_530), .B(n_528), .Y(n_916) );
O2A1O1Ixp5_ASAP7_75t_L g917 ( .A1(n_810), .A2(n_541), .B(n_543), .C(n_537), .Y(n_917) );
OR2x6_ASAP7_75t_L g918 ( .A(n_811), .B(n_546), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_816), .A2(n_550), .B1(n_551), .B2(n_549), .Y(n_919) );
BUFx6f_ASAP7_75t_L g920 ( .A(n_832), .Y(n_920) );
AND2x4_ASAP7_75t_L g921 ( .A(n_778), .B(n_552), .Y(n_921) );
AO31x2_ASAP7_75t_L g922 ( .A1(n_831), .A2(n_578), .A3(n_587), .B(n_577), .Y(n_922) );
AOI22xp33_ASAP7_75t_SL g923 ( .A1(n_834), .A2(n_560), .B1(n_564), .B2(n_557), .Y(n_923) );
BUFx6f_ASAP7_75t_L g924 ( .A(n_832), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_879), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_883), .A2(n_567), .B1(n_568), .B2(n_566), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_824), .B(n_636), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_846), .Y(n_928) );
INVx6_ASAP7_75t_L g929 ( .A(n_771), .Y(n_929) );
OAI21x1_ASAP7_75t_L g930 ( .A1(n_803), .A2(n_587), .B(n_578), .Y(n_930) );
OAI21x1_ASAP7_75t_L g931 ( .A1(n_752), .A2(n_587), .B(n_578), .Y(n_931) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_825), .A2(n_661), .B(n_647), .Y(n_932) );
OAI21x1_ASAP7_75t_L g933 ( .A1(n_752), .A2(n_590), .B(n_588), .Y(n_933) );
OAI21x1_ASAP7_75t_L g934 ( .A1(n_755), .A2(n_590), .B(n_588), .Y(n_934) );
OA21x2_ASAP7_75t_L g935 ( .A1(n_886), .A2(n_590), .B(n_588), .Y(n_935) );
NAND2x1p5_ASAP7_75t_L g936 ( .A(n_778), .B(n_592), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_766), .B(n_8), .Y(n_937) );
AOI21xp5_ASAP7_75t_L g938 ( .A1(n_842), .A2(n_661), .B(n_603), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_829), .Y(n_939) );
INVx3_ASAP7_75t_L g940 ( .A(n_777), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_854), .Y(n_941) );
OAI21x1_ASAP7_75t_L g942 ( .A1(n_755), .A2(n_603), .B(n_592), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_761), .B(n_9), .Y(n_943) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_796), .Y(n_944) );
A2O1A1Ixp33_ASAP7_75t_L g945 ( .A1(n_798), .A2(n_603), .B(n_613), .C(n_592), .Y(n_945) );
AOI221xp5_ASAP7_75t_L g946 ( .A1(n_785), .A2(n_613), .B1(n_586), .B2(n_583), .C(n_581), .Y(n_946) );
BUFx2_ASAP7_75t_L g947 ( .A(n_772), .Y(n_947) );
OAI21x1_ASAP7_75t_L g948 ( .A1(n_786), .A2(n_613), .B(n_583), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_783), .B(n_10), .Y(n_949) );
OAI21x1_ASAP7_75t_SL g950 ( .A1(n_807), .A2(n_10), .B(n_11), .Y(n_950) );
OR2x6_ASAP7_75t_L g951 ( .A(n_881), .B(n_12), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_861), .Y(n_952) );
CKINVDCx11_ASAP7_75t_R g953 ( .A(n_887), .Y(n_953) );
OA21x2_ASAP7_75t_L g954 ( .A1(n_889), .A2(n_583), .B(n_581), .Y(n_954) );
OAI21x1_ASAP7_75t_L g955 ( .A1(n_889), .A2(n_586), .B(n_583), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_787), .B(n_13), .Y(n_956) );
OR2x6_ASAP7_75t_L g957 ( .A(n_883), .B(n_13), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_796), .B(n_14), .Y(n_958) );
INVx1_ASAP7_75t_SL g959 ( .A(n_789), .Y(n_959) );
AOI21xp33_ASAP7_75t_SL g960 ( .A1(n_774), .A2(n_15), .B(n_16), .Y(n_960) );
AND2x4_ASAP7_75t_L g961 ( .A(n_758), .B(n_15), .Y(n_961) );
OAI21x1_ASAP7_75t_L g962 ( .A1(n_866), .A2(n_586), .B(n_123), .Y(n_962) );
BUFx2_ASAP7_75t_L g963 ( .A(n_772), .Y(n_963) );
NAND2x1p5_ASAP7_75t_L g964 ( .A(n_799), .B(n_815), .Y(n_964) );
OR2x6_ASAP7_75t_L g965 ( .A(n_859), .B(n_16), .Y(n_965) );
OR2x2_ASAP7_75t_L g966 ( .A(n_770), .B(n_760), .Y(n_966) );
OAI21x1_ASAP7_75t_L g967 ( .A1(n_833), .A2(n_586), .B(n_124), .Y(n_967) );
CKINVDCx16_ASAP7_75t_R g968 ( .A(n_782), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_806), .B(n_17), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_819), .Y(n_970) );
OA21x2_ASAP7_75t_L g971 ( .A1(n_792), .A2(n_586), .B(n_638), .Y(n_971) );
INVx4_ASAP7_75t_L g972 ( .A(n_799), .Y(n_972) );
A2O1A1Ixp33_ASAP7_75t_L g973 ( .A1(n_801), .A2(n_586), .B(n_652), .C(n_638), .Y(n_973) );
CKINVDCx5p33_ASAP7_75t_R g974 ( .A(n_809), .Y(n_974) );
OAI21x1_ASAP7_75t_L g975 ( .A1(n_821), .A2(n_125), .B(n_122), .Y(n_975) );
OR2x6_ASAP7_75t_L g976 ( .A(n_844), .B(n_18), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_823), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_849), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_849), .Y(n_979) );
OR3x4_ASAP7_75t_SL g980 ( .A(n_782), .B(n_18), .C(n_19), .Y(n_980) );
OAI21x1_ASAP7_75t_L g981 ( .A1(n_878), .A2(n_127), .B(n_126), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_845), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_797), .B(n_19), .Y(n_983) );
INVx3_ASAP7_75t_L g984 ( .A(n_777), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_837), .Y(n_985) );
OAI21x1_ASAP7_75t_L g986 ( .A1(n_853), .A2(n_134), .B(n_133), .Y(n_986) );
AOI21xp5_ASAP7_75t_L g987 ( .A1(n_873), .A2(n_652), .B(n_638), .Y(n_987) );
INVxp67_ASAP7_75t_SL g988 ( .A(n_791), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_773), .Y(n_989) );
OAI21x1_ASAP7_75t_L g990 ( .A1(n_853), .A2(n_141), .B(n_136), .Y(n_990) );
OR2x2_ASAP7_75t_L g991 ( .A(n_775), .B(n_21), .Y(n_991) );
BUFx2_ASAP7_75t_L g992 ( .A(n_799), .Y(n_992) );
O2A1O1Ixp5_ASAP7_75t_L g993 ( .A1(n_852), .A2(n_652), .B(n_638), .C(n_149), .Y(n_993) );
OAI21x1_ASAP7_75t_L g994 ( .A1(n_781), .A2(n_150), .B(n_142), .Y(n_994) );
INVx4_ASAP7_75t_SL g995 ( .A(n_815), .Y(n_995) );
OAI21xp5_ASAP7_75t_L g996 ( .A1(n_808), .A2(n_652), .B(n_638), .Y(n_996) );
NOR2xp33_ASAP7_75t_R g997 ( .A(n_815), .B(n_21), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_773), .B(n_22), .Y(n_998) );
AOI22xp33_ASAP7_75t_SL g999 ( .A1(n_827), .A2(n_25), .B1(n_23), .B2(n_24), .Y(n_999) );
AO31x2_ASAP7_75t_L g1000 ( .A1(n_890), .A2(n_652), .A3(n_25), .B(n_23), .Y(n_1000) );
OAI22xp33_ASAP7_75t_L g1001 ( .A1(n_838), .A2(n_27), .B1(n_24), .B2(n_26), .Y(n_1001) );
OA21x2_ASAP7_75t_L g1002 ( .A1(n_856), .A2(n_153), .B(n_152), .Y(n_1002) );
AOI21x1_ASAP7_75t_L g1003 ( .A1(n_855), .A2(n_155), .B(n_154), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_862), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_882), .B(n_27), .Y(n_1005) );
INVx2_ASAP7_75t_L g1006 ( .A(n_849), .Y(n_1006) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_874), .A2(n_30), .B1(n_28), .B2(n_29), .Y(n_1007) );
AO21x2_ASAP7_75t_L g1008 ( .A1(n_869), .A2(n_870), .B(n_858), .Y(n_1008) );
NAND2x1p5_ASAP7_75t_L g1009 ( .A(n_835), .B(n_32), .Y(n_1009) );
OAI21xp5_ASAP7_75t_L g1010 ( .A1(n_757), .A2(n_32), .B(n_33), .Y(n_1010) );
AND2x4_ASAP7_75t_L g1011 ( .A(n_781), .B(n_34), .Y(n_1011) );
OAI21x1_ASAP7_75t_L g1012 ( .A1(n_814), .A2(n_157), .B(n_156), .Y(n_1012) );
NAND2x1p5_ASAP7_75t_L g1013 ( .A(n_835), .B(n_34), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_857), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_868), .B(n_35), .Y(n_1015) );
AND2x4_ASAP7_75t_L g1016 ( .A(n_814), .B(n_36), .Y(n_1016) );
INVx4_ASAP7_75t_SL g1017 ( .A(n_882), .Y(n_1017) );
INVx8_ASAP7_75t_L g1018 ( .A(n_835), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_800), .Y(n_1019) );
BUFx2_ASAP7_75t_L g1020 ( .A(n_847), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_805), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_884), .Y(n_1022) );
AND2x4_ASAP7_75t_L g1023 ( .A(n_764), .B(n_37), .Y(n_1023) );
NOR2xp33_ASAP7_75t_SL g1024 ( .A(n_754), .B(n_161), .Y(n_1024) );
OAI21x1_ASAP7_75t_L g1025 ( .A1(n_751), .A2(n_163), .B(n_162), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_855), .A2(n_38), .B1(n_40), .B2(n_41), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_753), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_851), .B(n_38), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_875), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_857), .A2(n_40), .B1(n_41), .B2(n_42), .Y(n_1030) );
NAND3xp33_ASAP7_75t_L g1031 ( .A(n_877), .B(n_42), .C(n_44), .Y(n_1031) );
INVx8_ASAP7_75t_L g1032 ( .A(n_754), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_813), .B(n_44), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_872), .B(n_45), .Y(n_1034) );
AOI21xp5_ASAP7_75t_L g1035 ( .A1(n_830), .A2(n_166), .B(n_165), .Y(n_1035) );
NOR2xp67_ASAP7_75t_L g1036 ( .A(n_888), .B(n_168), .Y(n_1036) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_764), .B(n_46), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g1038 ( .A(n_780), .Y(n_1038) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_847), .Y(n_1039) );
AO21x1_ASAP7_75t_L g1040 ( .A1(n_812), .A2(n_175), .B(n_174), .Y(n_1040) );
AO21x2_ASAP7_75t_L g1041 ( .A1(n_841), .A2(n_178), .B(n_177), .Y(n_1041) );
OAI21xp5_ASAP7_75t_L g1042 ( .A1(n_871), .A2(n_47), .B(n_48), .Y(n_1042) );
OAI21x1_ASAP7_75t_L g1043 ( .A1(n_765), .A2(n_182), .B(n_181), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1044 ( .A(n_765), .B(n_47), .Y(n_1044) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_804), .B(n_49), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_847), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_1046) );
BUFx6f_ASAP7_75t_L g1047 ( .A(n_754), .Y(n_1047) );
INVx2_ASAP7_75t_L g1048 ( .A(n_857), .Y(n_1048) );
BUFx4f_ASAP7_75t_SL g1049 ( .A(n_839), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_867), .Y(n_1050) );
INVx2_ASAP7_75t_SL g1051 ( .A(n_839), .Y(n_1051) );
OAI21x1_ASAP7_75t_L g1052 ( .A1(n_864), .A2(n_188), .B(n_184), .Y(n_1052) );
INVx6_ASAP7_75t_L g1053 ( .A(n_839), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_826), .B(n_50), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_836), .Y(n_1055) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_822), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_867), .B(n_51), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_983), .B(n_865), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_925), .Y(n_1059) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_988), .A2(n_843), .B1(n_867), .B2(n_793), .Y(n_1060) );
AO21x2_ASAP7_75t_L g1061 ( .A1(n_996), .A2(n_795), .B(n_863), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_966), .A2(n_863), .B1(n_888), .B2(n_891), .Y(n_1062) );
A2O1A1Ixp33_ASAP7_75t_L g1063 ( .A1(n_1042), .A2(n_885), .B(n_776), .C(n_759), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_939), .Y(n_1064) );
OAI21x1_ASAP7_75t_L g1065 ( .A1(n_893), .A2(n_759), .B(n_756), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_957), .A2(n_891), .B1(n_885), .B2(n_776), .Y(n_1066) );
OAI21xp5_ASAP7_75t_L g1067 ( .A1(n_917), .A2(n_759), .B(n_756), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_957), .A2(n_885), .B1(n_776), .B2(n_756), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_983), .B(n_53), .Y(n_1069) );
AOI221xp5_ASAP7_75t_L g1070 ( .A1(n_1022), .A2(n_53), .B1(n_54), .B2(n_56), .C(n_59), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_957), .A2(n_54), .B1(n_60), .B2(n_61), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_1056), .A2(n_61), .B1(n_63), .B2(n_64), .Y(n_1072) );
A2O1A1Ixp33_ASAP7_75t_L g1073 ( .A1(n_1042), .A2(n_63), .B(n_64), .C(n_65), .Y(n_1073) );
AOI222xp33_ASAP7_75t_L g1074 ( .A1(n_1028), .A2(n_65), .B1(n_66), .B2(n_67), .C1(n_68), .C2(n_69), .Y(n_1074) );
OR2x6_ASAP7_75t_L g1075 ( .A(n_1018), .B(n_965), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_944), .B(n_66), .Y(n_1076) );
AND2x4_ASAP7_75t_L g1077 ( .A(n_1017), .B(n_68), .Y(n_1077) );
OAI22xp33_ASAP7_75t_L g1078 ( .A1(n_965), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_1033), .A2(n_71), .B1(n_72), .B2(n_73), .Y(n_1079) );
BUFx12f_ASAP7_75t_L g1080 ( .A(n_953), .Y(n_1080) );
OAI211xp5_ASAP7_75t_SL g1081 ( .A1(n_923), .A2(n_74), .B(n_75), .C(n_76), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_1038), .A2(n_74), .B1(n_75), .B2(n_76), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_985), .A2(n_77), .B1(n_78), .B2(n_79), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g1084 ( .A(n_900), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_901), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_982), .B(n_79), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1017), .B(n_80), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_1005), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_1045), .A2(n_1016), .B1(n_1011), .B2(n_910), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_989), .B(n_83), .Y(n_1090) );
AOI222xp33_ASAP7_75t_L g1091 ( .A1(n_947), .A2(n_84), .B1(n_85), .B2(n_87), .C1(n_88), .C2(n_89), .Y(n_1091) );
INVx2_ASAP7_75t_L g1092 ( .A(n_905), .Y(n_1092) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_919), .A2(n_87), .B1(n_88), .B2(n_89), .C(n_90), .Y(n_1093) );
OAI211xp5_ASAP7_75t_SL g1094 ( .A1(n_926), .A2(n_91), .B(n_92), .C(n_93), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1095 ( .A(n_918), .Y(n_1095) );
AO21x2_ASAP7_75t_L g1096 ( .A1(n_996), .A2(n_267), .B(n_379), .Y(n_1096) );
AOI221xp5_ASAP7_75t_L g1097 ( .A1(n_919), .A2(n_91), .B1(n_93), .B2(n_94), .C(n_95), .Y(n_1097) );
BUFx3_ASAP7_75t_L g1098 ( .A(n_963), .Y(n_1098) );
INVx5_ASAP7_75t_L g1099 ( .A(n_1018), .Y(n_1099) );
OAI221xp5_ASAP7_75t_SL g1100 ( .A1(n_951), .A2(n_94), .B1(n_96), .B2(n_97), .C(n_98), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_943), .Y(n_1101) );
AOI21xp5_ASAP7_75t_L g1102 ( .A1(n_987), .A2(n_271), .B(n_377), .Y(n_1102) );
OR2x4_ASAP7_75t_L g1103 ( .A(n_991), .B(n_1054), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_918), .A2(n_96), .B1(n_97), .B2(n_98), .Y(n_1104) );
AOI21xp5_ASAP7_75t_L g1105 ( .A1(n_987), .A2(n_275), .B(n_374), .Y(n_1105) );
INVx2_ASAP7_75t_L g1106 ( .A(n_915), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_1019), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_1107) );
INVx4_ASAP7_75t_SL g1108 ( .A(n_1049), .Y(n_1108) );
OAI221xp5_ASAP7_75t_L g1109 ( .A1(n_912), .A2(n_101), .B1(n_102), .B2(n_103), .C(n_104), .Y(n_1109) );
BUFx2_ASAP7_75t_R g1110 ( .A(n_974), .Y(n_1110) );
INVx3_ASAP7_75t_L g1111 ( .A(n_1018), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_943), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g1113 ( .A1(n_958), .A2(n_102), .B1(n_103), .B2(n_105), .Y(n_1113) );
INVxp67_ASAP7_75t_SL g1114 ( .A(n_1023), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_949), .Y(n_1115) );
AOI21xp33_ASAP7_75t_L g1116 ( .A1(n_894), .A2(n_105), .B(n_106), .Y(n_1116) );
AOI21xp5_ASAP7_75t_L g1117 ( .A1(n_1008), .A2(n_281), .B(n_372), .Y(n_1117) );
AOI21x1_ASAP7_75t_L g1118 ( .A1(n_899), .A2(n_280), .B(n_371), .Y(n_1118) );
OAI211xp5_ASAP7_75t_L g1119 ( .A1(n_960), .A2(n_106), .B(n_107), .C(n_109), .Y(n_1119) );
INVxp67_ASAP7_75t_L g1120 ( .A(n_937), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1121 ( .A1(n_998), .A2(n_107), .B1(n_109), .B2(n_110), .Y(n_1121) );
INVx2_ASAP7_75t_L g1122 ( .A(n_952), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_1055), .A2(n_110), .B1(n_111), .B2(n_112), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_976), .A2(n_112), .B1(n_113), .B2(n_114), .Y(n_1124) );
OAI22xp5_ASAP7_75t_L g1125 ( .A1(n_1007), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1126 ( .A1(n_965), .A2(n_115), .B1(n_116), .B2(n_117), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_949), .Y(n_1127) );
BUFx8_ASAP7_75t_L g1128 ( .A(n_895), .Y(n_1128) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_1007), .A2(n_117), .B1(n_191), .B2(n_193), .Y(n_1129) );
AOI221xp5_ASAP7_75t_L g1130 ( .A1(n_907), .A2(n_195), .B1(n_196), .B2(n_198), .C(n_200), .Y(n_1130) );
AO21x2_ASAP7_75t_L g1131 ( .A1(n_973), .A2(n_202), .B(n_208), .Y(n_1131) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_959), .A2(n_210), .B1(n_213), .B2(n_216), .Y(n_1132) );
OAI21xp5_ASAP7_75t_L g1133 ( .A1(n_904), .A2(n_218), .B(n_220), .Y(n_1133) );
OR2x6_ASAP7_75t_L g1134 ( .A(n_951), .B(n_221), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_976), .B(n_222), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_970), .B(n_226), .Y(n_1136) );
CKINVDCx5p33_ASAP7_75t_R g1137 ( .A(n_968), .Y(n_1137) );
INVx2_ASAP7_75t_L g1138 ( .A(n_977), .Y(n_1138) );
AOI21xp5_ASAP7_75t_L g1139 ( .A1(n_1008), .A2(n_227), .B(n_231), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1021), .Y(n_1140) );
INVx2_ASAP7_75t_L g1141 ( .A(n_928), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_976), .B(n_951), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_1023), .A2(n_233), .B1(n_234), .B2(n_235), .Y(n_1143) );
OAI21xp5_ASAP7_75t_L g1144 ( .A1(n_945), .A2(n_236), .B(n_237), .Y(n_1144) );
AOI221xp5_ASAP7_75t_L g1145 ( .A1(n_907), .A2(n_238), .B1(n_241), .B2(n_243), .C(n_245), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_1037), .A2(n_246), .B1(n_247), .B2(n_248), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g1147 ( .A1(n_961), .A2(n_252), .B1(n_254), .B2(n_258), .Y(n_1147) );
AOI221xp5_ASAP7_75t_L g1148 ( .A1(n_908), .A2(n_259), .B1(n_260), .B2(n_261), .C(n_263), .Y(n_1148) );
NOR2xp33_ASAP7_75t_SL g1149 ( .A(n_1009), .B(n_264), .Y(n_1149) );
INVx1_ASAP7_75t_SL g1150 ( .A(n_1020), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_1037), .A2(n_270), .B1(n_278), .B2(n_279), .Y(n_1151) );
OAI21xp33_ASAP7_75t_L g1152 ( .A1(n_1015), .A2(n_282), .B(n_284), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_1044), .A2(n_286), .B1(n_290), .B2(n_293), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_1044), .A2(n_294), .B1(n_295), .B2(n_298), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_1054), .A2(n_303), .B1(n_304), .B2(n_305), .Y(n_1155) );
AOI22xp33_ASAP7_75t_SL g1156 ( .A1(n_961), .A2(n_306), .B1(n_309), .B2(n_311), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1015), .B(n_312), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1158 ( .A1(n_908), .A2(n_314), .B1(n_315), .B2(n_316), .C(n_318), .Y(n_1158) );
AOI21xp5_ASAP7_75t_L g1159 ( .A1(n_927), .A2(n_319), .B(n_321), .Y(n_1159) );
AOI21xp5_ASAP7_75t_L g1160 ( .A1(n_927), .A2(n_322), .B(n_323), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1161 ( .A(n_959), .B(n_324), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_909), .B(n_326), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_956), .Y(n_1163) );
OA21x2_ASAP7_75t_L g1164 ( .A1(n_962), .A2(n_902), .B(n_967), .Y(n_1164) );
AND2x4_ASAP7_75t_L g1165 ( .A(n_995), .B(n_328), .Y(n_1165) );
CKINVDCx8_ASAP7_75t_R g1166 ( .A(n_980), .Y(n_1166) );
OA21x2_ASAP7_75t_L g1167 ( .A1(n_955), .A2(n_330), .B(n_332), .Y(n_1167) );
AOI222xp33_ASAP7_75t_L g1168 ( .A1(n_1026), .A2(n_334), .B1(n_336), .B2(n_337), .C1(n_339), .C2(n_342), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_921), .B(n_343), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_914), .B(n_344), .Y(n_1170) );
AOI22xp33_ASAP7_75t_SL g1171 ( .A1(n_997), .A2(n_345), .B1(n_347), .B2(n_350), .Y(n_1171) );
OAI22xp33_ASAP7_75t_L g1172 ( .A1(n_1026), .A2(n_355), .B1(n_356), .B2(n_358), .Y(n_1172) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_1009), .A2(n_359), .B1(n_360), .B2(n_361), .Y(n_1173) );
AND2x4_ASAP7_75t_L g1174 ( .A(n_920), .B(n_362), .Y(n_1174) );
NOR2xp33_ASAP7_75t_L g1175 ( .A(n_921), .B(n_363), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_1031), .A2(n_364), .B1(n_369), .B2(n_370), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_941), .Y(n_1177) );
OAI22xp33_ASAP7_75t_L g1178 ( .A1(n_1031), .A2(n_380), .B1(n_1013), .B2(n_1034), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_956), .B(n_969), .Y(n_1179) );
AOI221xp5_ASAP7_75t_L g1180 ( .A1(n_1001), .A2(n_1010), .B1(n_969), .B2(n_1030), .C(n_946), .Y(n_1180) );
AOI21xp5_ASAP7_75t_L g1181 ( .A1(n_932), .A2(n_935), .B(n_1040), .Y(n_1181) );
OR2x6_ASAP7_75t_L g1182 ( .A(n_929), .B(n_1013), .Y(n_1182) );
AND2x2_ASAP7_75t_SL g1183 ( .A(n_920), .B(n_924), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_1034), .A2(n_1010), .B1(n_999), .B2(n_1039), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1004), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1027), .B(n_1029), .Y(n_1186) );
INVx2_ASAP7_75t_L g1187 ( .A(n_924), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1030), .Y(n_1188) );
AOI22xp5_ASAP7_75t_SL g1189 ( .A1(n_929), .A2(n_936), .B1(n_940), .B2(n_984), .Y(n_1189) );
AOI21xp5_ASAP7_75t_L g1190 ( .A1(n_935), .A2(n_1035), .B(n_1002), .Y(n_1190) );
AOI221xp5_ASAP7_75t_L g1191 ( .A1(n_946), .A2(n_896), .B1(n_950), .B2(n_1046), .C(n_1057), .Y(n_1191) );
OAI22xp5_ASAP7_75t_L g1192 ( .A1(n_936), .A2(n_1057), .B1(n_898), .B2(n_897), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_992), .B(n_984), .Y(n_1193) );
OA21x2_ASAP7_75t_L g1194 ( .A1(n_986), .A2(n_990), .B(n_1025), .Y(n_1194) );
OAI21xp5_ASAP7_75t_L g1195 ( .A1(n_896), .A2(n_938), .B(n_903), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_940), .B(n_911), .Y(n_1196) );
INVx1_ASAP7_75t_SL g1197 ( .A(n_924), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1000), .Y(n_1198) );
BUFx3_ASAP7_75t_L g1199 ( .A(n_1053), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_911), .A2(n_972), .B1(n_1053), .B2(n_906), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1000), .Y(n_1201) );
A2O1A1Ixp33_ASAP7_75t_L g1202 ( .A1(n_913), .A2(n_916), .B(n_892), .C(n_938), .Y(n_1202) );
AND2x4_ASAP7_75t_L g1203 ( .A(n_972), .B(n_892), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_964), .A2(n_1051), .B1(n_1036), .B2(n_1050), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_964), .B(n_1006), .Y(n_1205) );
OA21x2_ASAP7_75t_L g1206 ( .A1(n_975), .A2(n_948), .B(n_981), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_978), .B(n_1014), .Y(n_1207) );
OAI211xp5_ASAP7_75t_L g1208 ( .A1(n_1003), .A2(n_971), .B(n_1002), .C(n_1036), .Y(n_1208) );
AOI21xp5_ASAP7_75t_L g1209 ( .A1(n_993), .A2(n_1024), .B(n_954), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_979), .A2(n_1048), .B1(n_1032), .B2(n_1047), .Y(n_1210) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_1041), .A2(n_1032), .B1(n_1024), .B2(n_971), .Y(n_1211) );
OAI211xp5_ASAP7_75t_L g1212 ( .A1(n_994), .A2(n_1012), .B(n_1052), .C(n_1043), .Y(n_1212) );
AO31x2_ASAP7_75t_L g1213 ( .A1(n_1041), .A2(n_922), .A3(n_1000), .B(n_954), .Y(n_1213) );
NOR2xp33_ASAP7_75t_L g1214 ( .A(n_1032), .B(n_1047), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_922), .B(n_1047), .Y(n_1215) );
OAI221xp5_ASAP7_75t_L g1216 ( .A1(n_1089), .A2(n_922), .B1(n_931), .B2(n_933), .C(n_934), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1114), .B(n_942), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1140), .B(n_930), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1058), .B(n_1069), .Y(n_1219) );
HB1xp67_ASAP7_75t_L g1220 ( .A(n_1084), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1085), .B(n_1092), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1106), .B(n_1122), .Y(n_1222) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1177), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1198), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1150), .B(n_1179), .Y(n_1225) );
AND2x4_ASAP7_75t_SL g1226 ( .A(n_1075), .B(n_1134), .Y(n_1226) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1185), .Y(n_1227) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1164), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1059), .Y(n_1229) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1150), .B(n_1101), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1064), .B(n_1112), .Y(n_1231) );
INVx2_ASAP7_75t_SL g1232 ( .A(n_1099), .Y(n_1232) );
HB1xp67_ASAP7_75t_L g1233 ( .A(n_1099), .Y(n_1233) );
AND2x4_ASAP7_75t_L g1234 ( .A(n_1099), .B(n_1182), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1201), .Y(n_1235) );
NOR2xp67_ASAP7_75t_L g1236 ( .A(n_1099), .B(n_1111), .Y(n_1236) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1164), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1115), .B(n_1127), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1163), .B(n_1138), .Y(n_1239) );
BUFx3_ASAP7_75t_L g1240 ( .A(n_1128), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1196), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1188), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1186), .B(n_1095), .Y(n_1243) );
BUFx2_ASAP7_75t_L g1244 ( .A(n_1182), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1215), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1207), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_1075), .A2(n_1134), .B1(n_1142), .B2(n_1081), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1103), .B(n_1120), .Y(n_1248) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1167), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1213), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1091), .B(n_1125), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1213), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1103), .B(n_1076), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1075), .B(n_1193), .Y(n_1254) );
INVx3_ASAP7_75t_SL g1255 ( .A(n_1108), .Y(n_1255) );
BUFx2_ASAP7_75t_L g1256 ( .A(n_1182), .Y(n_1256) );
BUFx2_ASAP7_75t_L g1257 ( .A(n_1183), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1086), .B(n_1074), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1213), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1091), .B(n_1125), .Y(n_1260) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1065), .Y(n_1261) );
AO21x2_ASAP7_75t_L g1262 ( .A1(n_1190), .A2(n_1195), .B(n_1181), .Y(n_1262) );
OR2x2_ASAP7_75t_L g1263 ( .A(n_1197), .B(n_1134), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1205), .Y(n_1264) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1197), .B(n_1090), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1074), .B(n_1168), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1168), .B(n_1073), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1187), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_1184), .A2(n_1094), .B1(n_1180), .B2(n_1129), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_1129), .A2(n_1078), .B1(n_1126), .B2(n_1109), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1136), .Y(n_1271) );
BUFx3_ASAP7_75t_L g1272 ( .A(n_1128), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1096), .Y(n_1273) );
INVxp67_ASAP7_75t_SL g1274 ( .A(n_1149), .Y(n_1274) );
HB1xp67_ASAP7_75t_L g1275 ( .A(n_1111), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1189), .B(n_1135), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1096), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1063), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1169), .B(n_1077), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1077), .B(n_1087), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1079), .B(n_1098), .Y(n_1281) );
INVxp67_ASAP7_75t_SL g1282 ( .A(n_1149), .Y(n_1282) );
INVxp33_ASAP7_75t_L g1283 ( .A(n_1214), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1071), .B(n_1072), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1157), .B(n_1174), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1174), .B(n_1083), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1121), .B(n_1113), .Y(n_1287) );
NOR3xp33_ASAP7_75t_L g1288 ( .A(n_1100), .B(n_1119), .C(n_1070), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1289 ( .A(n_1161), .B(n_1062), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1195), .Y(n_1290) );
NOR2x1_ASAP7_75t_SL g1291 ( .A(n_1173), .B(n_1192), .Y(n_1291) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1206), .Y(n_1292) );
NOR2xp33_ASAP7_75t_L g1293 ( .A(n_1166), .B(n_1137), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1199), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1093), .B(n_1097), .Y(n_1295) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1206), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1123), .B(n_1124), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1194), .Y(n_1298) );
HB1xp67_ASAP7_75t_L g1299 ( .A(n_1108), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1165), .B(n_1104), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_1116), .A2(n_1082), .B1(n_1088), .B2(n_1175), .Y(n_1301) );
BUFx3_ASAP7_75t_L g1302 ( .A(n_1165), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1194), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1304 ( .A1(n_1066), .A2(n_1068), .B1(n_1171), .B2(n_1060), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1107), .B(n_1061), .Y(n_1305) );
INVx2_ASAP7_75t_R g1306 ( .A(n_1208), .Y(n_1306) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1118), .Y(n_1307) );
INVx2_ASAP7_75t_L g1308 ( .A(n_1131), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1108), .Y(n_1309) );
BUFx3_ASAP7_75t_L g1310 ( .A(n_1080), .Y(n_1310) );
BUFx2_ASAP7_75t_L g1311 ( .A(n_1061), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1133), .B(n_1156), .Y(n_1312) );
OAI21x1_ASAP7_75t_L g1313 ( .A1(n_1209), .A2(n_1211), .B(n_1204), .Y(n_1313) );
HB1xp67_ASAP7_75t_L g1314 ( .A(n_1210), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1133), .B(n_1147), .Y(n_1315) );
INVx1_ASAP7_75t_SL g1316 ( .A(n_1110), .Y(n_1316) );
INVx2_ASAP7_75t_L g1317 ( .A(n_1131), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1212), .Y(n_1318) );
INVx3_ASAP7_75t_L g1319 ( .A(n_1203), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1203), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1067), .B(n_1200), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1067), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1202), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1172), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1178), .Y(n_1325) );
AND2x4_ASAP7_75t_L g1326 ( .A(n_1144), .B(n_1117), .Y(n_1326) );
BUFx6f_ASAP7_75t_L g1327 ( .A(n_1162), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1176), .Y(n_1328) );
BUFx2_ASAP7_75t_L g1329 ( .A(n_1144), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1143), .B(n_1153), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1146), .B(n_1154), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1152), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1139), .Y(n_1333) );
OAI211xp5_ASAP7_75t_L g1334 ( .A1(n_1130), .A2(n_1158), .B(n_1145), .C(n_1148), .Y(n_1334) );
INVx2_ASAP7_75t_L g1335 ( .A(n_1170), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g1336 ( .A(n_1132), .Y(n_1336) );
NOR2x1p5_ASAP7_75t_L g1337 ( .A(n_1151), .B(n_1155), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1191), .B(n_1102), .Y(n_1338) );
AND2x4_ASAP7_75t_L g1339 ( .A(n_1105), .B(n_1159), .Y(n_1339) );
INVx2_ASAP7_75t_L g1340 ( .A(n_1160), .Y(n_1340) );
INVx2_ASAP7_75t_L g1341 ( .A(n_1141), .Y(n_1341) );
BUFx3_ASAP7_75t_L g1342 ( .A(n_1240), .Y(n_1342) );
OR2x2_ASAP7_75t_L g1343 ( .A(n_1243), .B(n_1225), .Y(n_1343) );
NAND4xp25_ASAP7_75t_L g1344 ( .A(n_1269), .B(n_1247), .C(n_1248), .D(n_1270), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1229), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1227), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1280), .B(n_1221), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1227), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1239), .Y(n_1349) );
OR2x2_ASAP7_75t_L g1350 ( .A(n_1243), .B(n_1225), .Y(n_1350) );
INVx4_ASAP7_75t_L g1351 ( .A(n_1302), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1239), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1280), .B(n_1221), .Y(n_1353) );
AND2x4_ASAP7_75t_L g1354 ( .A(n_1242), .B(n_1245), .Y(n_1354) );
BUFx12f_ASAP7_75t_L g1355 ( .A(n_1240), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1356 ( .A(n_1230), .B(n_1220), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1238), .B(n_1231), .Y(n_1357) );
OR2x2_ASAP7_75t_L g1358 ( .A(n_1230), .B(n_1223), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1222), .B(n_1279), .Y(n_1359) );
INVx2_ASAP7_75t_L g1360 ( .A(n_1228), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1238), .B(n_1231), .Y(n_1361) );
INVx3_ASAP7_75t_L g1362 ( .A(n_1234), .Y(n_1362) );
NAND4xp25_ASAP7_75t_SL g1363 ( .A(n_1316), .B(n_1251), .C(n_1260), .D(n_1266), .Y(n_1363) );
OR2x2_ASAP7_75t_L g1364 ( .A(n_1341), .B(n_1264), .Y(n_1364) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1219), .B(n_1251), .Y(n_1365) );
INVx2_ASAP7_75t_SL g1366 ( .A(n_1234), .Y(n_1366) );
INVxp67_ASAP7_75t_L g1367 ( .A(n_1245), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1222), .Y(n_1368) );
OAI321xp33_ASAP7_75t_L g1369 ( .A1(n_1266), .A2(n_1260), .A3(n_1267), .B1(n_1304), .B2(n_1258), .C(n_1318), .Y(n_1369) );
NAND4xp25_ASAP7_75t_L g1370 ( .A(n_1253), .B(n_1288), .C(n_1301), .D(n_1281), .Y(n_1370) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1237), .Y(n_1371) );
INVx4_ASAP7_75t_L g1372 ( .A(n_1302), .Y(n_1372) );
INVx2_ASAP7_75t_L g1373 ( .A(n_1237), .Y(n_1373) );
INVxp67_ASAP7_75t_L g1374 ( .A(n_1263), .Y(n_1374) );
INVx4_ASAP7_75t_L g1375 ( .A(n_1226), .Y(n_1375) );
NAND2xp5_ASAP7_75t_SL g1376 ( .A(n_1312), .B(n_1315), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1279), .B(n_1283), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1233), .B(n_1232), .Y(n_1378) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1298), .Y(n_1379) );
NAND3xp33_ASAP7_75t_L g1380 ( .A(n_1318), .B(n_1242), .C(n_1325), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1232), .B(n_1276), .Y(n_1381) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1246), .Y(n_1382) );
INVxp67_ASAP7_75t_SL g1383 ( .A(n_1274), .Y(n_1383) );
AND2x4_ASAP7_75t_L g1384 ( .A(n_1224), .B(n_1235), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1276), .B(n_1226), .Y(n_1385) );
BUFx2_ASAP7_75t_L g1386 ( .A(n_1234), .Y(n_1386) );
BUFx3_ASAP7_75t_L g1387 ( .A(n_1272), .Y(n_1387) );
AND2x4_ASAP7_75t_L g1388 ( .A(n_1224), .B(n_1235), .Y(n_1388) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1298), .Y(n_1389) );
NAND3xp33_ASAP7_75t_L g1390 ( .A(n_1325), .B(n_1267), .C(n_1338), .Y(n_1390) );
INVx3_ASAP7_75t_L g1391 ( .A(n_1319), .Y(n_1391) );
OR2x2_ASAP7_75t_L g1392 ( .A(n_1264), .B(n_1254), .Y(n_1392) );
HB1xp67_ASAP7_75t_L g1393 ( .A(n_1241), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1275), .B(n_1294), .Y(n_1394) );
INVx1_ASAP7_75t_SL g1395 ( .A(n_1272), .Y(n_1395) );
INVx2_ASAP7_75t_L g1396 ( .A(n_1303), .Y(n_1396) );
OAI221xp5_ASAP7_75t_SL g1397 ( .A1(n_1287), .A2(n_1295), .B1(n_1300), .B2(n_1284), .C(n_1244), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1236), .B(n_1244), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1256), .B(n_1246), .Y(n_1399) );
OR2x2_ASAP7_75t_L g1400 ( .A(n_1254), .B(n_1263), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1268), .Y(n_1401) );
INVx2_ASAP7_75t_SL g1402 ( .A(n_1256), .Y(n_1402) );
INVx5_ASAP7_75t_L g1403 ( .A(n_1319), .Y(n_1403) );
INVx2_ASAP7_75t_L g1404 ( .A(n_1303), .Y(n_1404) );
AND2x4_ASAP7_75t_L g1405 ( .A(n_1320), .B(n_1319), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1295), .B(n_1284), .Y(n_1406) );
INVxp67_ASAP7_75t_L g1407 ( .A(n_1241), .Y(n_1407) );
INVxp67_ASAP7_75t_SL g1408 ( .A(n_1282), .Y(n_1408) );
INVx5_ASAP7_75t_SL g1409 ( .A(n_1255), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1257), .B(n_1297), .Y(n_1410) );
OR2x6_ASAP7_75t_L g1411 ( .A(n_1257), .B(n_1300), .Y(n_1411) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1268), .Y(n_1412) );
BUFx6f_ASAP7_75t_L g1413 ( .A(n_1255), .Y(n_1413) );
OAI321xp33_ASAP7_75t_L g1414 ( .A1(n_1324), .A2(n_1329), .A3(n_1305), .B1(n_1311), .B2(n_1321), .C(n_1289), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1297), .B(n_1285), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1285), .B(n_1286), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1265), .Y(n_1417) );
INVx3_ASAP7_75t_L g1418 ( .A(n_1255), .Y(n_1418) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1265), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1309), .Y(n_1420) );
BUFx2_ASAP7_75t_L g1421 ( .A(n_1299), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1422 ( .A1(n_1324), .A2(n_1286), .B1(n_1337), .B2(n_1305), .Y(n_1422) );
AOI22xp33_ASAP7_75t_SL g1423 ( .A1(n_1291), .A2(n_1329), .B1(n_1336), .B2(n_1330), .Y(n_1423) );
OAI211xp5_ASAP7_75t_L g1424 ( .A1(n_1293), .A2(n_1320), .B(n_1334), .C(n_1314), .Y(n_1424) );
INVx2_ASAP7_75t_L g1425 ( .A(n_1292), .Y(n_1425) );
INVx2_ASAP7_75t_L g1426 ( .A(n_1296), .Y(n_1426) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1218), .Y(n_1427) );
INVx2_ASAP7_75t_L g1428 ( .A(n_1296), .Y(n_1428) );
OR2x2_ASAP7_75t_L g1429 ( .A(n_1289), .B(n_1217), .Y(n_1429) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1218), .Y(n_1430) );
HB1xp67_ASAP7_75t_L g1431 ( .A(n_1393), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_1427), .B(n_1250), .Y(n_1432) );
BUFx3_ASAP7_75t_L g1433 ( .A(n_1413), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1349), .B(n_1271), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_1352), .B(n_1271), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1430), .B(n_1259), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1384), .Y(n_1437) );
AND2x4_ASAP7_75t_L g1438 ( .A(n_1354), .B(n_1252), .Y(n_1438) );
INVx1_ASAP7_75t_SL g1439 ( .A(n_1421), .Y(n_1439) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1384), .Y(n_1440) );
BUFx3_ASAP7_75t_L g1441 ( .A(n_1413), .Y(n_1441) );
OR2x2_ASAP7_75t_L g1442 ( .A(n_1429), .B(n_1290), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1354), .B(n_1290), .Y(n_1443) );
INVxp67_ASAP7_75t_SL g1444 ( .A(n_1393), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1354), .B(n_1311), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1384), .Y(n_1446) );
NOR2x1_ASAP7_75t_L g1447 ( .A(n_1375), .B(n_1418), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1388), .B(n_1321), .Y(n_1448) );
INVxp67_ASAP7_75t_SL g1449 ( .A(n_1407), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1450 ( .A(n_1417), .B(n_1328), .Y(n_1450) );
NOR2xp33_ASAP7_75t_L g1451 ( .A(n_1395), .B(n_1342), .Y(n_1451) );
INVx2_ASAP7_75t_L g1452 ( .A(n_1379), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1388), .B(n_1322), .Y(n_1453) );
INVx2_ASAP7_75t_L g1454 ( .A(n_1379), .Y(n_1454) );
OR2x2_ASAP7_75t_L g1455 ( .A(n_1343), .B(n_1322), .Y(n_1455) );
INVx2_ASAP7_75t_L g1456 ( .A(n_1389), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1388), .B(n_1323), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1389), .Y(n_1458) );
AND2x4_ASAP7_75t_L g1459 ( .A(n_1396), .B(n_1313), .Y(n_1459) );
INVx1_ASAP7_75t_SL g1460 ( .A(n_1378), .Y(n_1460) );
BUFx2_ASAP7_75t_L g1461 ( .A(n_1386), .Y(n_1461) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1404), .Y(n_1462) );
AND2x4_ASAP7_75t_L g1463 ( .A(n_1404), .B(n_1313), .Y(n_1463) );
INVx2_ASAP7_75t_L g1464 ( .A(n_1360), .Y(n_1464) );
AND2x4_ASAP7_75t_L g1465 ( .A(n_1362), .B(n_1261), .Y(n_1465) );
AND2x4_ASAP7_75t_L g1466 ( .A(n_1362), .B(n_1261), .Y(n_1466) );
OR2x2_ASAP7_75t_L g1467 ( .A(n_1350), .B(n_1262), .Y(n_1467) );
AOI21xp33_ASAP7_75t_L g1468 ( .A1(n_1424), .A2(n_1278), .B(n_1328), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1347), .B(n_1262), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1353), .B(n_1273), .Y(n_1470) );
CKINVDCx16_ASAP7_75t_R g1471 ( .A(n_1355), .Y(n_1471) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1419), .B(n_1330), .Y(n_1472) );
NAND2xp5_ASAP7_75t_L g1473 ( .A(n_1368), .B(n_1331), .Y(n_1473) );
NAND2xp5_ASAP7_75t_L g1474 ( .A(n_1357), .B(n_1331), .Y(n_1474) );
NAND2xp5_ASAP7_75t_L g1475 ( .A(n_1361), .B(n_1335), .Y(n_1475) );
BUFx2_ASAP7_75t_L g1476 ( .A(n_1351), .Y(n_1476) );
OR2x2_ASAP7_75t_L g1477 ( .A(n_1400), .B(n_1278), .Y(n_1477) );
NAND3xp33_ASAP7_75t_L g1478 ( .A(n_1370), .B(n_1333), .C(n_1273), .Y(n_1478) );
HB1xp67_ASAP7_75t_L g1479 ( .A(n_1356), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1365), .B(n_1335), .Y(n_1480) );
INVx4_ASAP7_75t_L g1481 ( .A(n_1375), .Y(n_1481) );
INVxp67_ASAP7_75t_L g1482 ( .A(n_1387), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1359), .B(n_1277), .Y(n_1483) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1374), .B(n_1277), .Y(n_1484) );
OR2x2_ASAP7_75t_L g1485 ( .A(n_1358), .B(n_1317), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1376), .B(n_1306), .Y(n_1486) );
NOR2xp33_ASAP7_75t_L g1487 ( .A(n_1387), .B(n_1310), .Y(n_1487) );
AOI221xp5_ASAP7_75t_L g1488 ( .A1(n_1369), .A2(n_1216), .B1(n_1333), .B2(n_1326), .C(n_1339), .Y(n_1488) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1406), .B(n_1291), .Y(n_1489) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1346), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1376), .B(n_1306), .Y(n_1491) );
INVxp67_ASAP7_75t_L g1492 ( .A(n_1377), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1348), .Y(n_1493) );
INVx2_ASAP7_75t_L g1494 ( .A(n_1371), .Y(n_1494) );
NAND3xp33_ASAP7_75t_SL g1495 ( .A(n_1423), .B(n_1332), .C(n_1308), .Y(n_1495) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1410), .B(n_1249), .Y(n_1496) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1479), .Y(n_1497) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1431), .Y(n_1498) );
INVx2_ASAP7_75t_L g1499 ( .A(n_1452), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1500 ( .A(n_1474), .B(n_1390), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1501 ( .A(n_1469), .B(n_1428), .Y(n_1501) );
OAI31xp33_ASAP7_75t_L g1502 ( .A1(n_1476), .A2(n_1363), .A3(n_1344), .B(n_1397), .Y(n_1502) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1449), .Y(n_1503) );
NAND2xp5_ASAP7_75t_L g1504 ( .A(n_1470), .B(n_1422), .Y(n_1504) );
NAND2xp5_ASAP7_75t_L g1505 ( .A(n_1470), .B(n_1422), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1469), .B(n_1428), .Y(n_1506) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1448), .B(n_1373), .Y(n_1507) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1490), .Y(n_1508) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1483), .B(n_1345), .Y(n_1509) );
AND3x1_ASAP7_75t_L g1510 ( .A(n_1487), .B(n_1385), .C(n_1355), .Y(n_1510) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1490), .Y(n_1511) );
INVx2_ASAP7_75t_SL g1512 ( .A(n_1476), .Y(n_1512) );
OR2x2_ASAP7_75t_L g1513 ( .A(n_1460), .B(n_1407), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1448), .B(n_1426), .Y(n_1514) );
OR2x6_ASAP7_75t_L g1515 ( .A(n_1481), .B(n_1375), .Y(n_1515) );
NAND2xp5_ASAP7_75t_L g1516 ( .A(n_1483), .B(n_1415), .Y(n_1516) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1443), .B(n_1426), .Y(n_1517) );
INVxp67_ASAP7_75t_L g1518 ( .A(n_1439), .Y(n_1518) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1493), .Y(n_1519) );
AOI21xp33_ASAP7_75t_SL g1520 ( .A1(n_1471), .A2(n_1397), .B(n_1418), .Y(n_1520) );
INVx2_ASAP7_75t_L g1521 ( .A(n_1452), .Y(n_1521) );
OR2x6_ASAP7_75t_L g1522 ( .A(n_1481), .B(n_1411), .Y(n_1522) );
AOI221xp5_ASAP7_75t_L g1523 ( .A1(n_1492), .A2(n_1414), .B1(n_1382), .B2(n_1420), .C(n_1416), .Y(n_1523) );
AND2x4_ASAP7_75t_L g1524 ( .A(n_1437), .B(n_1383), .Y(n_1524) );
INVx1_ASAP7_75t_SL g1525 ( .A(n_1471), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1443), .B(n_1373), .Y(n_1526) );
NAND2xp5_ASAP7_75t_L g1527 ( .A(n_1473), .B(n_1367), .Y(n_1527) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1493), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1529 ( .A(n_1453), .B(n_1425), .Y(n_1529) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1444), .Y(n_1530) );
INVxp67_ASAP7_75t_SL g1531 ( .A(n_1447), .Y(n_1531) );
NAND2xp5_ASAP7_75t_L g1532 ( .A(n_1472), .B(n_1367), .Y(n_1532) );
NAND2xp5_ASAP7_75t_L g1533 ( .A(n_1439), .B(n_1399), .Y(n_1533) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1434), .Y(n_1534) );
HB1xp67_ASAP7_75t_L g1535 ( .A(n_1461), .Y(n_1535) );
AND2x4_ASAP7_75t_L g1536 ( .A(n_1437), .B(n_1408), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_1453), .B(n_1425), .Y(n_1537) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1435), .Y(n_1538) );
NAND2xp5_ASAP7_75t_L g1539 ( .A(n_1477), .B(n_1392), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_1460), .B(n_1381), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_1477), .B(n_1401), .Y(n_1541) );
AND2x4_ASAP7_75t_SL g1542 ( .A(n_1481), .B(n_1413), .Y(n_1542) );
OR2x2_ASAP7_75t_L g1543 ( .A(n_1442), .B(n_1411), .Y(n_1543) );
INVx2_ASAP7_75t_SL g1544 ( .A(n_1447), .Y(n_1544) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1432), .Y(n_1545) );
NOR2xp33_ASAP7_75t_L g1546 ( .A(n_1489), .B(n_1482), .Y(n_1546) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1432), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1436), .Y(n_1548) );
NAND2xp5_ASAP7_75t_L g1549 ( .A(n_1534), .B(n_1467), .Y(n_1549) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1498), .Y(n_1550) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1503), .Y(n_1551) );
AOI221xp5_ASAP7_75t_L g1552 ( .A1(n_1520), .A2(n_1478), .B1(n_1468), .B2(n_1446), .C(n_1440), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1553 ( .A(n_1509), .B(n_1467), .Y(n_1553) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1540), .B(n_1445), .Y(n_1554) );
AND2x4_ASAP7_75t_L g1555 ( .A(n_1512), .B(n_1440), .Y(n_1555) );
OAI22x1_ASAP7_75t_L g1556 ( .A1(n_1525), .A2(n_1481), .B1(n_1461), .B2(n_1451), .Y(n_1556) );
NAND2x1_ASAP7_75t_L g1557 ( .A(n_1515), .B(n_1351), .Y(n_1557) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1545), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1559 ( .A(n_1500), .B(n_1436), .Y(n_1559) );
OR2x2_ASAP7_75t_L g1560 ( .A(n_1539), .B(n_1455), .Y(n_1560) );
AOI22xp33_ASAP7_75t_SL g1561 ( .A1(n_1515), .A2(n_1372), .B1(n_1351), .B2(n_1366), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1507), .B(n_1445), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1507), .B(n_1457), .Y(n_1563) );
CKINVDCx20_ASAP7_75t_R g1564 ( .A(n_1533), .Y(n_1564) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1538), .B(n_1484), .Y(n_1565) );
INVx2_ASAP7_75t_L g1566 ( .A(n_1513), .Y(n_1566) );
AOI22xp5_ASAP7_75t_L g1567 ( .A1(n_1510), .A2(n_1438), .B1(n_1480), .B2(n_1491), .Y(n_1567) );
OAI321xp33_ASAP7_75t_L g1568 ( .A1(n_1515), .A2(n_1495), .A3(n_1478), .B1(n_1486), .B2(n_1491), .C(n_1488), .Y(n_1568) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1547), .Y(n_1569) );
OAI22xp5_ASAP7_75t_L g1570 ( .A1(n_1515), .A2(n_1372), .B1(n_1366), .B2(n_1446), .Y(n_1570) );
OAI21xp5_ASAP7_75t_L g1571 ( .A1(n_1502), .A2(n_1380), .B(n_1372), .Y(n_1571) );
AOI221xp5_ASAP7_75t_L g1572 ( .A1(n_1523), .A2(n_1450), .B1(n_1394), .B2(n_1475), .C(n_1486), .Y(n_1572) );
OR2x2_ASAP7_75t_L g1573 ( .A(n_1516), .B(n_1455), .Y(n_1573) );
INVx2_ASAP7_75t_L g1574 ( .A(n_1535), .Y(n_1574) );
AOI22xp33_ASAP7_75t_SL g1575 ( .A1(n_1531), .A2(n_1398), .B1(n_1441), .B2(n_1433), .Y(n_1575) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1548), .Y(n_1576) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1497), .Y(n_1577) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1530), .B(n_1484), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1579 ( .A(n_1501), .B(n_1458), .Y(n_1579) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1508), .Y(n_1580) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1511), .Y(n_1581) );
OAI22xp5_ASAP7_75t_L g1582 ( .A1(n_1522), .A2(n_1409), .B1(n_1438), .B2(n_1403), .Y(n_1582) );
AOI211xp5_ASAP7_75t_L g1583 ( .A1(n_1571), .A2(n_1546), .B(n_1505), .C(n_1504), .Y(n_1583) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1578), .Y(n_1584) );
AOI322xp5_ASAP7_75t_L g1585 ( .A1(n_1572), .A2(n_1518), .A3(n_1546), .B1(n_1535), .B2(n_1514), .C1(n_1527), .C2(n_1541), .Y(n_1585) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1549), .B(n_1514), .Y(n_1586) );
OAI21xp33_ASAP7_75t_SL g1587 ( .A1(n_1567), .A2(n_1522), .B(n_1544), .Y(n_1587) );
INVx2_ASAP7_75t_L g1588 ( .A(n_1574), .Y(n_1588) );
NOR2x1p5_ASAP7_75t_L g1589 ( .A(n_1557), .B(n_1413), .Y(n_1589) );
INVxp67_ASAP7_75t_L g1590 ( .A(n_1556), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1554), .B(n_1501), .Y(n_1591) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1578), .Y(n_1592) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1551), .Y(n_1593) );
NAND2xp5_ASAP7_75t_L g1594 ( .A(n_1558), .B(n_1517), .Y(n_1594) );
AOI21xp5_ASAP7_75t_L g1595 ( .A1(n_1571), .A2(n_1522), .B(n_1542), .Y(n_1595) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1579), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1562), .B(n_1506), .Y(n_1597) );
OAI221xp5_ASAP7_75t_L g1598 ( .A1(n_1552), .A2(n_1532), .B1(n_1543), .B2(n_1528), .C(n_1519), .Y(n_1598) );
INVx1_ASAP7_75t_SL g1599 ( .A(n_1564), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1569), .B(n_1526), .Y(n_1600) );
CKINVDCx14_ASAP7_75t_R g1601 ( .A(n_1582), .Y(n_1601) );
AOI22xp5_ASAP7_75t_L g1602 ( .A1(n_1559), .A2(n_1517), .B1(n_1537), .B2(n_1526), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1566), .B(n_1506), .Y(n_1603) );
NAND2xp5_ASAP7_75t_L g1604 ( .A(n_1576), .B(n_1537), .Y(n_1604) );
NAND2xp5_ASAP7_75t_L g1605 ( .A(n_1577), .B(n_1529), .Y(n_1605) );
OAI21xp33_ASAP7_75t_L g1606 ( .A1(n_1585), .A2(n_1565), .B(n_1575), .Y(n_1606) );
OA22x2_ASAP7_75t_L g1607 ( .A1(n_1590), .A2(n_1582), .B1(n_1570), .B2(n_1542), .Y(n_1607) );
INVx2_ASAP7_75t_L g1608 ( .A(n_1588), .Y(n_1608) );
AOI22xp5_ASAP7_75t_L g1609 ( .A1(n_1601), .A2(n_1561), .B1(n_1570), .B2(n_1550), .Y(n_1609) );
O2A1O1Ixp33_ASAP7_75t_L g1610 ( .A1(n_1598), .A2(n_1568), .B(n_1565), .C(n_1560), .Y(n_1610) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1596), .Y(n_1611) );
AOI22xp5_ASAP7_75t_L g1612 ( .A1(n_1601), .A2(n_1555), .B1(n_1553), .B2(n_1573), .Y(n_1612) );
O2A1O1Ixp33_ASAP7_75t_L g1613 ( .A1(n_1583), .A2(n_1581), .B(n_1580), .C(n_1408), .Y(n_1613) );
AOI222xp33_ASAP7_75t_L g1614 ( .A1(n_1587), .A2(n_1555), .B1(n_1579), .B2(n_1563), .C1(n_1536), .C2(n_1524), .Y(n_1614) );
OAI211xp5_ASAP7_75t_SL g1615 ( .A1(n_1599), .A2(n_1391), .B(n_1412), .C(n_1383), .Y(n_1615) );
OAI22xp5_ASAP7_75t_SL g1616 ( .A1(n_1589), .A2(n_1441), .B1(n_1433), .B2(n_1403), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_1597), .B(n_1536), .Y(n_1617) );
XOR2x2_ASAP7_75t_L g1618 ( .A(n_1595), .B(n_1524), .Y(n_1618) );
OAI22xp5_ASAP7_75t_L g1619 ( .A1(n_1602), .A2(n_1409), .B1(n_1441), .B2(n_1433), .Y(n_1619) );
AOI221xp5_ASAP7_75t_SL g1620 ( .A1(n_1606), .A2(n_1592), .B1(n_1584), .B2(n_1605), .C(n_1593), .Y(n_1620) );
AOI22xp5_ASAP7_75t_L g1621 ( .A1(n_1609), .A2(n_1604), .B1(n_1600), .B2(n_1594), .Y(n_1621) );
AOI21xp33_ASAP7_75t_SL g1622 ( .A1(n_1607), .A2(n_1588), .B(n_1586), .Y(n_1622) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1610), .B(n_1591), .Y(n_1623) );
INVx1_ASAP7_75t_SL g1624 ( .A(n_1618), .Y(n_1624) );
AOI221xp5_ASAP7_75t_L g1625 ( .A1(n_1613), .A2(n_1591), .B1(n_1597), .B2(n_1603), .C(n_1438), .Y(n_1625) );
NAND3xp33_ASAP7_75t_L g1626 ( .A(n_1609), .B(n_1614), .C(n_1612), .Y(n_1626) );
O2A1O1Ixp33_ASAP7_75t_L g1627 ( .A1(n_1615), .A2(n_1402), .B(n_1391), .C(n_1603), .Y(n_1627) );
O2A1O1Ixp33_ASAP7_75t_L g1628 ( .A1(n_1619), .A2(n_1402), .B(n_1391), .C(n_1332), .Y(n_1628) );
OR2x2_ASAP7_75t_L g1629 ( .A(n_1623), .B(n_1611), .Y(n_1629) );
AND3x4_ASAP7_75t_L g1630 ( .A(n_1624), .B(n_1616), .C(n_1608), .Y(n_1630) );
AOI211xp5_ASAP7_75t_L g1631 ( .A1(n_1626), .A2(n_1617), .B(n_1405), .C(n_1326), .Y(n_1631) );
XNOR2xp5_ASAP7_75t_L g1632 ( .A(n_1621), .B(n_1405), .Y(n_1632) );
OAI21xp5_ASAP7_75t_L g1633 ( .A1(n_1620), .A2(n_1403), .B(n_1405), .Y(n_1633) );
OAI222xp33_ASAP7_75t_L g1634 ( .A1(n_1627), .A2(n_1364), .B1(n_1485), .B2(n_1521), .C1(n_1499), .C2(n_1458), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1622), .B(n_1496), .Y(n_1635) );
NAND3xp33_ASAP7_75t_SL g1636 ( .A(n_1630), .B(n_1625), .C(n_1628), .Y(n_1636) );
OAI222xp33_ASAP7_75t_L g1637 ( .A1(n_1629), .A2(n_1628), .B1(n_1485), .B2(n_1499), .C1(n_1521), .C2(n_1462), .Y(n_1637) );
OAI21xp5_ASAP7_75t_L g1638 ( .A1(n_1636), .A2(n_1631), .B(n_1632), .Y(n_1638) );
OAI22x1_ASAP7_75t_L g1639 ( .A1(n_1637), .A2(n_1635), .B1(n_1634), .B2(n_1633), .Y(n_1639) );
INVx2_ASAP7_75t_L g1640 ( .A(n_1639), .Y(n_1640) );
OAI22xp5_ASAP7_75t_SL g1641 ( .A1(n_1638), .A2(n_1339), .B1(n_1340), .B2(n_1307), .Y(n_1641) );
INVx2_ASAP7_75t_L g1642 ( .A(n_1640), .Y(n_1642) );
AOI22xp33_ASAP7_75t_L g1643 ( .A1(n_1641), .A2(n_1466), .B1(n_1465), .B2(n_1463), .Y(n_1643) );
OR2x2_ASAP7_75t_L g1644 ( .A(n_1642), .B(n_1456), .Y(n_1644) );
OAI22xp33_ASAP7_75t_L g1645 ( .A1(n_1644), .A2(n_1643), .B1(n_1327), .B2(n_1456), .Y(n_1645) );
AOI222xp33_ASAP7_75t_L g1646 ( .A1(n_1645), .A2(n_1459), .B1(n_1463), .B2(n_1454), .C1(n_1494), .C2(n_1464), .Y(n_1646) );
endmodule