module fake_jpeg_14830_n_150 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_150);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_28),
.B(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_15),
.B(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_30),
.Y(n_44)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_43),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_14),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_18),
.B1(n_26),
.B2(n_29),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_34),
.B1(n_32),
.B2(n_13),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_59),
.B1(n_17),
.B2(n_24),
.Y(n_75)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_13),
.B1(n_21),
.B2(n_36),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_21),
.B1(n_36),
.B2(n_30),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_41),
.B1(n_50),
.B2(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_64),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_33),
.C(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_46),
.B(n_33),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_71),
.C(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_78),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_58),
.B1(n_57),
.B2(n_52),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_24),
.C(n_23),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_37),
.B(n_27),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_31),
.B(n_41),
.C(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_76),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_48),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_57),
.Y(n_85)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_77),
.C(n_73),
.Y(n_96)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_52),
.B1(n_17),
.B2(n_55),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_74),
.B(n_22),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_45),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_87),
.C(n_81),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_71),
.B1(n_77),
.B2(n_69),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_87),
.B(n_92),
.Y(n_112)
);

NOR4xp25_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_78),
.C(n_54),
.D(n_75),
.Y(n_100)
);

NOR4xp25_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_91),
.C(n_106),
.D(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_104),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_31),
.B1(n_48),
.B2(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_54),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_115),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_112),
.B(n_114),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_37),
.C(n_86),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_107),
.B1(n_102),
.B2(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_45),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_116),
.B(n_117),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g117 ( 
.A(n_97),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_19),
.B(n_1),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_118),
.A2(n_0),
.B(n_1),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_86),
.B(n_37),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_127),
.B(n_2),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_99),
.B1(n_10),
.B2(n_12),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_12),
.C(n_25),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_129),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_122),
.B(n_27),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_2),
.B(n_3),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_134),
.C(n_133),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_119),
.C(n_123),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_136),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_25),
.C(n_27),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_3),
.B(n_4),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_139),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_31),
.C(n_6),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_5),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_143),
.C(n_140),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_6),
.A3(n_7),
.B1(n_9),
.B2(n_142),
.C1(n_146),
.C2(n_147),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_9),
.Y(n_150)
);


endmodule