module fake_jpeg_25115_n_106 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_SL g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_50),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_38),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_56),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_34),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_45),
.B1(n_44),
.B2(n_41),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_43),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_39),
.Y(n_69)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_72),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_9),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_19),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_3),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_13),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_21),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_87),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_SL g82 ( 
.A(n_79),
.B(n_4),
.C(n_7),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_86),
.B(n_89),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_10),
.B(n_11),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_14),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_16),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_67),
.C(n_76),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_80),
.C(n_22),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_77),
.B1(n_65),
.B2(n_27),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_88),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_84),
.B(n_83),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_95),
.C(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_97),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_94),
.B(n_28),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_17),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_29),
.Y(n_106)
);


endmodule