module fake_netlist_1_12530_n_14 (n_1, n_2, n_4, n_3, n_5, n_0, n_14);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_9;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_SL g6 ( .A(n_0), .Y(n_6) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_5), .B(n_4), .Y(n_7) );
AOI22xp33_ASAP7_75t_L g8 ( .A1(n_2), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_8) );
BUFx2_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
INVx1_ASAP7_75t_SL g11 ( .A(n_10), .Y(n_11) );
AOI22xp33_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_9), .B1(n_8), .B2(n_2), .Y(n_12) );
OR2x6_ASAP7_75t_L g13 ( .A(n_12), .B(n_9), .Y(n_13) );
NAND2xp5_ASAP7_75t_SL g14 ( .A(n_13), .B(n_1), .Y(n_14) );
endmodule