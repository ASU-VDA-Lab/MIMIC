module fake_ariane_2125_n_192 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_192);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_192;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_30;
wire n_178;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_188;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_87;
wire n_81;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

INVxp67_ASAP7_75t_SL g31 ( 
.A(n_24),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVxp33_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_0),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_R g63 ( 
.A(n_38),
.B(n_14),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_46),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_46),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_32),
.B1(n_45),
.B2(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_40),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

AO22x2_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_87),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_62),
.B(n_66),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_52),
.B(n_62),
.C(n_71),
.Y(n_94)
);

OR2x2_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_64),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_63),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_65),
.B1(n_67),
.B2(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_72),
.B(n_71),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

BUFx2_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

OAI21x1_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_92),
.B(n_97),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_84),
.B1(n_78),
.B2(n_72),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

AO21x2_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_86),
.B(n_88),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_73),
.B(n_30),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_87),
.C(n_73),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_96),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_102),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_100),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_81),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_99),
.Y(n_116)
);

AO31x2_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_94),
.A3(n_93),
.B(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_107),
.B(n_98),
.C(n_86),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_113),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_110),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_110),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_110),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_112),
.Y(n_134)
);

NAND3x1_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_102),
.C(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_84),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_128),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_125),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_124),
.B(n_127),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_131),
.B1(n_112),
.B2(n_110),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_131),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_125),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_148),
.B(n_74),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

AOI222xp33_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_74),
.B1(n_107),
.B2(n_84),
.C1(n_146),
.C2(n_70),
.Y(n_158)
);

OAI211xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_145),
.B(n_71),
.C(n_70),
.Y(n_159)
);

AOI221xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_84),
.B1(n_71),
.B2(n_69),
.C(n_81),
.Y(n_160)
);

NAND4xp25_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_149),
.C(n_69),
.D(n_81),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_135),
.B1(n_146),
.B2(n_69),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_114),
.Y(n_163)
);

OAI21x1_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_114),
.B(n_2),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_88),
.Y(n_166)
);

AOI321xp33_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_151),
.A3(n_80),
.B1(n_79),
.B2(n_77),
.C(n_7),
.Y(n_167)
);

OAI211xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_158),
.B(n_159),
.C(n_165),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_163),
.B1(n_164),
.B2(n_160),
.Y(n_169)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.C(n_5),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_106),
.B(n_103),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_106),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_0),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_174)
);

OAI211xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_4),
.B(n_8),
.C(n_9),
.Y(n_175)
);

AOI221xp5_ASAP7_75t_SL g176 ( 
.A1(n_173),
.A2(n_9),
.B1(n_12),
.B2(n_16),
.C(n_18),
.Y(n_176)
);

OR3x2_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_19),
.C(n_21),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_172),
.Y(n_180)
);

NAND4xp75_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_50),
.C(n_27),
.D(n_28),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_182),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_175),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_177),
.B1(n_181),
.B2(n_111),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_185),
.B1(n_188),
.B2(n_187),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_185),
.B1(n_186),
.B2(n_183),
.C(n_177),
.Y(n_192)
);


endmodule