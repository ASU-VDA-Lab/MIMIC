module fake_jpeg_177_n_193 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_193);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g85 ( 
.A(n_75),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_65),
.B1(n_52),
.B2(n_68),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_76),
.B1(n_64),
.B2(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_76),
.A2(n_57),
.B1(n_62),
.B2(n_50),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_55),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_93),
.B1(n_94),
.B2(n_62),
.Y(n_107)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_70),
.B1(n_71),
.B2(n_60),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_60),
.B1(n_54),
.B2(n_63),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_49),
.A3(n_66),
.B1(n_53),
.B2(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_104),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_50),
.C(n_51),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_19),
.C(n_45),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_50),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_57),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_106),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_89),
.B1(n_82),
.B2(n_51),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_122),
.B1(n_32),
.B2(n_44),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_89),
.B1(n_56),
.B2(n_69),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_125),
.B1(n_121),
.B2(n_120),
.Y(n_147)
);

BUFx24_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_116),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_0),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_11),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_10),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_56),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_126),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_48),
.B1(n_22),
.B2(n_24),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_18),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_131),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_4),
.C(n_5),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_8),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_8),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_134),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_9),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_137),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_10),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_140),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_11),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_122),
.B(n_121),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_146),
.B(n_12),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_12),
.B(n_13),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

AOI221xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_161),
.B1(n_34),
.B2(n_35),
.C(n_36),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_33),
.C(n_43),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_162),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_136),
.B1(n_144),
.B2(n_127),
.C(n_147),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_47),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_30),
.C(n_37),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_25),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_160),
.A2(n_140),
.B(n_141),
.C(n_146),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_170),
.B(n_164),
.C(n_148),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_168),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_169),
.B(n_171),
.Y(n_178)
);

FAx1_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_13),
.CI(n_14),
.CON(n_170),
.SN(n_170)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_174),
.B1(n_158),
.B2(n_163),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_180),
.B1(n_181),
.B2(n_166),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_162),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_179),
.C(n_152),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_156),
.C(n_151),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_155),
.B(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_175),
.B(n_166),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_178),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_185),
.B(n_176),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_187),
.A2(n_188),
.B1(n_182),
.B2(n_149),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_186),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_41),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_17),
.C(n_15),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_16),
.Y(n_193)
);


endmodule