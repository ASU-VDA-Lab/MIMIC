module fake_jpeg_20781_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_26),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_29),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_53),
.C(n_44),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_29),
.B1(n_34),
.B2(n_31),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_34),
.B1(n_30),
.B2(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_19),
.B1(n_24),
.B2(n_26),
.Y(n_96)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_27),
.Y(n_87)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_24),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_45),
.B1(n_39),
.B2(n_33),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

NAND2x1p5_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_32),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_23),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_36),
.B(n_37),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_71),
.A2(n_77),
.B(n_109),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_81),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_28),
.B1(n_27),
.B2(n_39),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_75),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_1),
.Y(n_134)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_17),
.Y(n_79)
);

NOR2x1_ASAP7_75t_R g137 ( 
.A(n_79),
.B(n_2),
.Y(n_137)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_86),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_104),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_21),
.C(n_22),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_90),
.A2(n_97),
.B(n_0),
.Y(n_133)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_45),
.B1(n_19),
.B2(n_28),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_23),
.C(n_22),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_26),
.B(n_16),
.C(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_22),
.A3(n_21),
.B1(n_23),
.B2(n_19),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_19),
.B1(n_43),
.B2(n_38),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_101),
.A2(n_89),
.B1(n_79),
.B2(n_86),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_25),
.B1(n_17),
.B2(n_35),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_107),
.B1(n_2),
.B2(n_3),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_43),
.C(n_35),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_112),
.C(n_65),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_25),
.B1(n_17),
.B2(n_35),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_50),
.B(n_25),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_43),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_38),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_113),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_133),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_71),
.A2(n_20),
.B(n_18),
.C(n_35),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_132),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_0),
.C(n_1),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_77),
.C(n_88),
.Y(n_150)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_74),
.B(n_0),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_85),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_142),
.B1(n_110),
.B2(n_99),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_83),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_143),
.B1(n_91),
.B2(n_80),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_144),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_167),
.B1(n_175),
.B2(n_119),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_77),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_160),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_104),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_152),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_103),
.C(n_112),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_159),
.C(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_78),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_136),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_100),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_112),
.C(n_109),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_81),
.Y(n_160)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_164),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_116),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_98),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_73),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_109),
.C(n_101),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_130),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_174),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_114),
.B(n_111),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_132),
.B(n_141),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_114),
.B(n_92),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_143),
.A3(n_122),
.B1(n_138),
.B2(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_137),
.B(n_132),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_177),
.A2(n_194),
.B(n_204),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_172),
.B1(n_171),
.B2(n_159),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_8),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_169),
.A2(n_134),
.B1(n_124),
.B2(n_122),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_184),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_230)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_168),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_186),
.B(n_196),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_127),
.C(n_115),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_8),
.C(n_9),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_127),
.B1(n_126),
.B2(n_120),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_192),
.B1(n_207),
.B2(n_160),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_126),
.B1(n_120),
.B2(n_106),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_146),
.A2(n_82),
.B(n_123),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_173),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_123),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_198),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_150),
.B(n_123),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_161),
.A2(n_94),
.B1(n_78),
.B2(n_73),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_203),
.B1(n_157),
.B2(n_149),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_146),
.A2(n_72),
.B1(n_110),
.B2(n_118),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_5),
.B(n_6),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_72),
.B1(n_118),
.B2(n_7),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_151),
.A2(n_118),
.B(n_6),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_210),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_178),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_216),
.B1(n_201),
.B2(n_203),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_212),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_206),
.B(n_145),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_213),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_145),
.B1(n_170),
.B2(n_164),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_226),
.B1(n_228),
.B2(n_235),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_174),
.B1(n_168),
.B2(n_162),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_162),
.Y(n_221)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_149),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_230),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_157),
.B1(n_6),
.B2(n_7),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_204),
.Y(n_246)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_202),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_182),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_235),
.A2(n_187),
.B1(n_194),
.B2(n_183),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_224),
.B1(n_199),
.B2(n_223),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_190),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_251),
.C(n_257),
.Y(n_260)
);

NAND2x1_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_196),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_236),
.C(n_219),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_226),
.B1(n_179),
.B2(n_216),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_246),
.B(n_257),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_197),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_239),
.B1(n_243),
.B2(n_248),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_272),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_261),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_256),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_266),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_223),
.B(n_177),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_276),
.B(n_277),
.Y(n_286)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_224),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_265),
.B(n_267),
.Y(n_290)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_254),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_179),
.C(n_184),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_244),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_251),
.B(n_231),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_245),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_182),
.B1(n_205),
.B2(n_207),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_238),
.A2(n_219),
.B(n_205),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_234),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_284),
.Y(n_296)
);

OAI32xp33_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_250),
.A3(n_249),
.B1(n_253),
.B2(n_255),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_283),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_277),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_225),
.B1(n_222),
.B2(n_229),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_232),
.B1(n_222),
.B2(n_200),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_289),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_264),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_237),
.B1(n_246),
.B2(n_209),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_241),
.B1(n_237),
.B2(n_230),
.Y(n_291)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_208),
.B1(n_215),
.B2(n_11),
.Y(n_292)
);

OAI22x1_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_267),
.B1(n_263),
.B2(n_268),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_286),
.A2(n_265),
.B(n_269),
.Y(n_295)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_287),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_271),
.B(n_264),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_272),
.B(n_260),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_301),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_8),
.C(n_9),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_11),
.B(n_12),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_302),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_292),
.B1(n_290),
.B2(n_281),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_305),
.A2(n_307),
.B1(n_294),
.B2(n_302),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_290),
.B1(n_280),
.B2(n_284),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_288),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_309),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_304),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_278),
.C(n_303),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_315),
.B(n_311),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_282),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_318),
.B(n_297),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_305),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_306),
.B1(n_307),
.B2(n_303),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_322),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_316),
.B(n_293),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_309),
.Y(n_326)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_320),
.B(n_324),
.Y(n_327)
);

OAI321xp33_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_301),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_11),
.Y(n_328)
);

O2A1O1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_13),
.B(n_14),
.C(n_247),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_13),
.Y(n_330)
);


endmodule