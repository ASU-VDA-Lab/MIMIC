module fake_jpeg_4958_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_20),
.B(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_40),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_1),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_31),
.C(n_28),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_20),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_59),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_20),
.B1(n_30),
.B2(n_23),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_61),
.B1(n_21),
.B2(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_28),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_24),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_63),
.B(n_27),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_23),
.B1(n_30),
.B2(n_21),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_64),
.B(n_55),
.C(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_22),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_23),
.B1(n_31),
.B2(n_28),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_24),
.B(n_16),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_19),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_73),
.B1(n_64),
.B2(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_71),
.Y(n_88)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_69),
.B(n_70),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_29),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_82),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_32),
.B1(n_29),
.B2(n_17),
.Y(n_73)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_32),
.B1(n_45),
.B2(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_51),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_59),
.B(n_47),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_50),
.B(n_22),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_55),
.B1(n_62),
.B2(n_49),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_92),
.B1(n_97),
.B2(n_79),
.Y(n_117)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_93),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_63),
.C(n_57),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_95),
.C(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_45),
.B1(n_51),
.B2(n_58),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_74),
.B1(n_68),
.B2(n_25),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_95),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_80),
.B(n_29),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_108),
.C(n_115),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_73),
.C(n_78),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_73),
.B(n_70),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_121),
.B(n_86),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_66),
.B1(n_51),
.B2(n_49),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_119),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_117),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_77),
.C(n_62),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_49),
.B1(n_77),
.B2(n_27),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_102),
.B1(n_101),
.B2(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_137),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_135),
.B(n_138),
.Y(n_155)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_136),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_85),
.C(n_99),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_132),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_133),
.B1(n_138),
.B2(n_136),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_91),
.C(n_102),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_89),
.B(n_84),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_96),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_125),
.B(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_46),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_2),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_114),
.A3(n_121),
.B1(n_112),
.B2(n_122),
.C1(n_119),
.C2(n_111),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_SL g168 ( 
.A(n_144),
.B(n_127),
.C(n_11),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_112),
.B1(n_110),
.B2(n_62),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_149),
.B1(n_128),
.B2(n_134),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_110),
.B1(n_107),
.B2(n_17),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_151),
.B(n_153),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_80),
.B(n_18),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_162),
.B(n_2),
.Y(n_178)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_157),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_29),
.B(n_17),
.C(n_18),
.D(n_46),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_130),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_60),
.B1(n_46),
.B2(n_100),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_60),
.B1(n_18),
.B2(n_5),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_29),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_171),
.B(n_172),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_168),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_127),
.B1(n_100),
.B2(n_18),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_60),
.C(n_46),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_175),
.C(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_150),
.B1(n_148),
.B2(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_60),
.C(n_15),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.C(n_6),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

AOI321xp33_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_155),
.A3(n_160),
.B1(n_157),
.B2(n_162),
.C(n_9),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_4),
.C(n_7),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_155),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_189),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_186),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_190),
.B(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_187),
.C(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_196),
.C(n_198),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_168),
.B1(n_166),
.B2(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_195),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_184),
.B(n_13),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_179),
.B(n_189),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_10),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_200),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_4),
.Y(n_200)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_197),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_180),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_207),
.B(n_194),
.Y(n_210)
);

NOR2x1_ASAP7_75t_SL g207 ( 
.A(n_198),
.B(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_211),
.B(n_213),
.C(n_10),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_8),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_205),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_8),
.B(n_10),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_215),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_204),
.C(n_209),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_220),
.C(n_219),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_204),
.B(n_203),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_221),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_218),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_222),
.Y(n_224)
);


endmodule