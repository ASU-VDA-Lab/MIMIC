module real_jpeg_7400_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_1),
.A2(n_26),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_1),
.A2(n_40),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_1),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_1),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_1),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_1),
.A2(n_182),
.B1(n_231),
.B2(n_234),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_1),
.A2(n_263),
.B(n_266),
.C(n_269),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_1),
.B(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_1),
.B(n_102),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_1),
.B(n_121),
.C(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_1),
.B(n_90),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_1),
.B(n_86),
.C(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_1),
.B(n_33),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_2),
.A2(n_92),
.B1(n_93),
.B2(n_97),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_2),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_2),
.A2(n_80),
.B1(n_92),
.B2(n_124),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_2),
.A2(n_92),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_3),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_64),
.B1(n_147),
.B2(n_151),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_3),
.A2(n_64),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_4),
.Y(n_108)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_4),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_5),
.Y(n_389)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_7),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_7),
.Y(n_175)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_7),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_7),
.Y(n_277)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_10),
.A2(n_28),
.B1(n_154),
.B2(n_158),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_10),
.A2(n_28),
.B1(n_202),
.B2(n_205),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_10),
.A2(n_28),
.B1(n_171),
.B2(n_275),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_11),
.Y(n_271)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_12),
.Y(n_385)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_13),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_384),
.B(n_386),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_189),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_188),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_138),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_19),
.B(n_138),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_130),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_128),
.B2(n_129),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_56),
.B2(n_57),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_23),
.A2(n_24),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_23),
.A2(n_24),
.B1(n_152),
.B2(n_338),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_24),
.B(n_197),
.C(n_219),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_24),
.B(n_152),
.C(n_261),
.Y(n_260)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B1(n_52),
.B2(n_55),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_25),
.A2(n_32),
.B1(n_52),
.B2(n_55),
.Y(n_128)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_32),
.A2(n_52),
.B(n_55),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_42),
.Y(n_32)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_35),
.Y(n_137)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_40),
.Y(n_268)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_99),
.B2(n_127),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_66),
.B1(n_90),
.B2(n_91),
.Y(n_59)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_66),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_67),
.A2(n_78),
.B1(n_135),
.B2(n_153),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_67),
.A2(n_78),
.B1(n_135),
.B2(n_153),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_67),
.B(n_78),
.Y(n_238)
);

NAND2x1_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_78),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_74),
.Y(n_320)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_78),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

AOI22x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_82),
.Y(n_186)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_84),
.Y(n_322)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_128),
.C(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_127),
.B1(n_131),
.B2(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_126),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_100),
.B(n_179),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_115),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_101),
.A2(n_115),
.B1(n_200),
.B2(n_206),
.Y(n_199)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_102),
.A2(n_116),
.B1(n_126),
.B2(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_102),
.A2(n_146),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_102),
.B(n_201),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_109),
.B2(n_113),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g211 ( 
.A(n_108),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_108),
.Y(n_233)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_122),
.B2(n_124),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_119),
.Y(n_301)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_128),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_129),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_128),
.B(n_224),
.C(n_237),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_128),
.A2(n_129),
.B1(n_237),
.B2(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_128),
.A2(n_129),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_128),
.B(n_219),
.C(n_348),
.Y(n_365)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_134),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g266 ( 
.A1(n_136),
.A2(n_264),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_160),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_139),
.A2(n_143),
.B1(n_144),
.B2(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_139),
.Y(n_381)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_144),
.A2(n_145),
.B(n_152),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_152),
.A2(n_334),
.B1(n_335),
.B2(n_338),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_152),
.Y(n_338)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_160),
.B(n_380),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B(n_187),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_161),
.B(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_176),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_162),
.A2(n_176),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_162),
.A2(n_187),
.B1(n_222),
.B2(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_165),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_165),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_168),
.B(n_230),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_208),
.B1(n_213),
.B2(n_214),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_169),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_170),
.A2(n_230),
.B1(n_274),
.B2(n_277),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_170),
.A2(n_230),
.B1(n_274),
.B2(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_171),
.Y(n_289)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_174),
.Y(n_292)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_178),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_378),
.B(n_383),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI211xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_278),
.B(n_372),
.C(n_377),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_250),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_194),
.A2(n_250),
.B(n_373),
.C(n_376),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_239),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_195),
.B(n_239),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_220),
.C(n_223),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_196),
.B(n_220),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_217),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_207),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_198),
.A2(n_199),
.B1(n_207),
.B2(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_198),
.A2(n_199),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_198),
.A2(n_199),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_199),
.B(n_273),
.C(n_310),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_199),
.B(n_330),
.C(n_332),
.Y(n_343)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_218),
.A2(n_219),
.B1(n_235),
.B2(n_299),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_218),
.B(n_299),
.C(n_317),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_218),
.A2(n_219),
.B1(n_348),
.B2(n_349),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_252),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_235),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_226),
.A2(n_235),
.B1(n_299),
.B2(n_364),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_226),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_235),
.A2(n_299),
.B1(n_300),
.B2(n_304),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_235),
.Y(n_299)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_248),
.B2(n_249),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_241)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_245),
.B(n_247),
.C(n_249),
.Y(n_382)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_251),
.B(n_253),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.C(n_260),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_255),
.B(n_258),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_260),
.B(n_371),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_261),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_272),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_262),
.A2(n_272),
.B1(n_273),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_262),
.Y(n_355)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_272),
.A2(n_273),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_273),
.B(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_294),
.Y(n_295)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_357),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_342),
.B(n_356),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_327),
.B(n_341),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_314),
.B(n_326),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_306),
.B(n_313),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_296),
.B(n_305),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_293),
.B(n_295),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_291),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_291),
.A2(n_297),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_297),
.B(n_336),
.C(n_338),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_304),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_300),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_312),
.Y(n_313)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_316),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_325),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_323),
.B2(n_324),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_324),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_340),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_340),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_332),
.B1(n_333),
.B2(n_339),
.Y(n_328)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_329),
.Y(n_339)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_330),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_343),
.B(n_344),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_352),
.C(n_353),
.Y(n_366)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_348),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NOR2x1_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_367),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_366),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_366),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_360),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_363),
.B(n_365),
.C(n_369),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_367),
.A2(n_374),
.B(n_375),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_368),
.B(n_370),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_382),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_382),
.Y(n_383)
);

INVx8_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx13_ASAP7_75t_L g388 ( 
.A(n_385),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);


endmodule