module fake_jpeg_28177_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_3),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_17),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_18),
.Y(n_34)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_28),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_22),
.C(n_18),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_11),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_20),
.B1(n_13),
.B2(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_18),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_10),
.C(n_25),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_42),
.Y(n_55)
);

AND2x6_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_8),
.Y(n_47)
);

OAI322xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_4),
.A3(n_7),
.B1(n_15),
.B2(n_0),
.C1(n_1),
.C2(n_3),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_21),
.B1(n_25),
.B2(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_24),
.B1(n_37),
.B2(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_54),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_38),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_57),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_51),
.Y(n_58)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_47),
.B(n_46),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_45),
.C(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_7),
.Y(n_66)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_63),
.B(n_65),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_62),
.B(n_65),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_24),
.B1(n_1),
.B2(n_3),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_0),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_68),
.Y(n_72)
);

AOI221xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_24),
.B1(n_60),
.B2(n_71),
.C(n_67),
.Y(n_73)
);


endmodule