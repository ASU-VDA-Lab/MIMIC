module fake_aes_7805_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g10 ( .A(n_2), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_4), .B(n_7), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_4), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
A2O1A1Ixp33_ASAP7_75t_L g18 ( .A1(n_11), .A2(n_1), .B(n_2), .C(n_3), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_10), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_12), .B(n_3), .Y(n_20) );
INVxp67_ASAP7_75t_SL g21 ( .A(n_14), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_10), .B1(n_13), .B2(n_15), .Y(n_22) );
NOR2xp33_ASAP7_75t_R g23 ( .A(n_17), .B(n_16), .Y(n_23) );
NOR2x1_ASAP7_75t_SL g24 ( .A(n_20), .B(n_10), .Y(n_24) );
AND3x1_ASAP7_75t_L g25 ( .A(n_18), .B(n_5), .C(n_6), .Y(n_25) );
NAND2x1p5_ASAP7_75t_L g26 ( .A(n_25), .B(n_20), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
HB1xp67_ASAP7_75t_L g28 ( .A(n_23), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_26), .A2(n_22), .B1(n_25), .B2(n_19), .Y(n_30) );
AOI211xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_28), .B(n_26), .C(n_19), .Y(n_31) );
OAI211xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_17), .B(n_24), .C(n_5), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_31), .Y(n_33) );
INVx1_ASAP7_75t_SL g34 ( .A(n_32), .Y(n_34) );
CKINVDCx20_ASAP7_75t_R g35 ( .A(n_33), .Y(n_35) );
AOI22xp33_ASAP7_75t_SL g36 ( .A1(n_35), .A2(n_34), .B1(n_8), .B2(n_9), .Y(n_36) );
endmodule