module real_jpeg_16542_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_518),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_0),
.B(n_519),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_1),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_1),
.B(n_94),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_1),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_1),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_1),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_1),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_SL g328 ( 
.A(n_1),
.B(n_329),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_2),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_2),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_2),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_3),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_3),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_3),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_3),
.B(n_294),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_3),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_3),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_3),
.B(n_436),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_3),
.B(n_466),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_4),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_5),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_5),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_5),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_5),
.Y(n_292)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_5),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_6),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_6),
.B(n_111),
.Y(n_110)
);

AND2x4_ASAP7_75t_SL g139 ( 
.A(n_6),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_6),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_6),
.B(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_7),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_7),
.Y(n_233)
);

BUFx4f_ASAP7_75t_L g495 ( 
.A(n_7),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_8),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_8),
.B(n_213),
.Y(n_212)
);

AOI22x1_ASAP7_75t_SL g259 ( 
.A1(n_8),
.A2(n_17),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_8),
.B(n_67),
.Y(n_333)
);

AOI31xp33_ASAP7_75t_L g369 ( 
.A1(n_8),
.A2(n_259),
.A3(n_370),
.B(n_375),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_8),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_8),
.B(n_448),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_8),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_8),
.B(n_37),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_9),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_9),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_9),
.B(n_94),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_9),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_9),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_9),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_9),
.B(n_373),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_10),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_10),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_10),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_10),
.B(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_11),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_11),
.B(n_220),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_11),
.B(n_240),
.Y(n_239)
);

AND2x4_ASAP7_75t_SL g284 ( 
.A(n_11),
.B(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_11),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_11),
.B(n_382),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_11),
.B(n_330),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_12),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_12),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_13),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_14),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_14),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_14),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_14),
.B(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_14),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_14),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_14),
.B(n_493),
.Y(n_492)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_15),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_15),
.Y(n_119)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_15),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_15),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_16),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_17),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_17),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_17),
.B(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_17),
.B(n_231),
.Y(n_230)
);

NAND2x1_ASAP7_75t_L g234 ( 
.A(n_17),
.B(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_17),
.Y(n_371)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_18),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_18),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_196),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_195),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_165),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_24),
.B(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_114),
.C(n_129),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_25),
.A2(n_26),
.B1(n_114),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_72),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_54),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_28),
.B(n_167),
.C(n_168),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_43),
.C(n_49),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_29),
.A2(n_30),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_36),
.C(n_39),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_31),
.A2(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_31),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_31),
.A2(n_36),
.B1(n_83),
.B2(n_148),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_32),
.B(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_34),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_36),
.B(n_135),
.C(n_139),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_36),
.Y(n_148)
);

AOI22x1_ASAP7_75t_L g209 ( 
.A1(n_36),
.A2(n_139),
.B1(n_148),
.B2(n_210),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_39),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_39),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_39),
.A2(n_145),
.B1(n_272),
.B2(n_322),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_41),
.Y(n_188)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_42),
.Y(n_152)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_42),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_43),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_44),
.B(n_49),
.Y(n_163)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_45),
.B(n_227),
.C(n_230),
.Y(n_226)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_47),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_49),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_49),
.A2(n_158),
.B1(n_161),
.B2(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_52),
.Y(n_241)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_53),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g407 ( 
.A(n_53),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_54),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_55),
.B(n_65),
.C(n_71),
.Y(n_194)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_70),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_84),
.C(n_98),
.Y(n_72)
);

XNOR2x2_ASAP7_75t_SL g204 ( 
.A(n_73),
.B(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_80),
.C(n_83),
.Y(n_127)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_80),
.B1(n_117),
.B2(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g175 ( 
.A(n_80),
.B(n_117),
.C(n_121),
.Y(n_175)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_81),
.Y(n_432)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_82),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_84),
.B(n_98),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.C(n_93),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_87),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_88),
.Y(n_286)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_97),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_104),
.C(n_110),
.Y(n_128)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_102),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_110),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_114),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_126),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_115),
.B(n_127),
.C(n_128),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_117),
.A2(n_120),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_129),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_149),
.C(n_162),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_144),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_132),
.B(n_134),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_135),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

BUFx2_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_143),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_144),
.B(n_304),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_145),
.B(n_267),
.C(n_272),
.Y(n_266)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_162),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.C(n_161),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_150),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_157),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_151),
.B(n_157),
.Y(n_224)
);

XOR2x1_ASAP7_75t_SL g223 ( 
.A(n_153),
.B(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_158),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_160),
.Y(n_283)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_185),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

XOR2x1_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_182),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_194),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_192),
.Y(n_295)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_192),
.Y(n_378)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_515),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_249),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_246),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_200),
.B(n_246),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.C(n_206),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g349 ( 
.A(n_202),
.B(n_204),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_206),
.B(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_225),
.C(n_242),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_207),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_223),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_208),
.B(n_211),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.C(n_218),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_212),
.A2(n_218),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_212),
.Y(n_346)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_215),
.B(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_218),
.B(n_404),
.C(n_408),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_218),
.A2(n_345),
.B1(n_404),
.B2(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_219),
.Y(n_345)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_223),
.B(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_225),
.B(n_243),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.C(n_238),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_226),
.B(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_230),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_228),
.Y(n_466)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_229),
.Y(n_331)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_233),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_233),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_234),
.A2(n_238),
.B1(n_239),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_234),
.Y(n_299)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_238),
.A2(n_239),
.B1(n_385),
.B2(n_386),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_239),
.B(n_380),
.C(n_385),
.Y(n_379)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AO21x2_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_354),
.B(n_512),
.Y(n_249)
);

NOR2xp67_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_347),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_307),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_252),
.B(n_307),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_300),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_253),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_275),
.C(n_296),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_255),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.C(n_266),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_256),
.B(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_258),
.A2(n_259),
.B1(n_266),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_266),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_267),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_269),
.Y(n_446)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_274),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_276),
.A2(n_296),
.B1(n_297),
.B2(n_312),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_276),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_287),
.C(n_293),
.Y(n_276)
);

XOR2x2_ASAP7_75t_L g341 ( 
.A(n_277),
.B(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_282),
.C(n_284),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_278),
.A2(n_284),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_278),
.Y(n_368)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_282),
.B(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_284),
.Y(n_367)
);

XNOR2x1_ASAP7_75t_L g458 ( 
.A(n_284),
.B(n_459),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_286),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_293),
.Y(n_342)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_291),
.Y(n_450)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_300)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_303),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_305),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.C(n_316),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_309),
.A2(n_310),
.B1(n_314),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_358),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_341),
.C(n_343),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_318),
.B(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.C(n_332),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g413 ( 
.A(n_320),
.B(n_414),
.Y(n_413)
);

XNOR2x1_ASAP7_75t_L g414 ( 
.A(n_323),
.B(n_332),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_324),
.B(n_328),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.C(n_339),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_333),
.A2(n_334),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_334),
.A2(n_401),
.B1(n_482),
.B2(n_483),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_334),
.B(n_478),
.C(n_482),
.Y(n_502)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_339),
.B(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_343),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_347),
.A2(n_513),
.B(n_514),
.Y(n_512)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_348),
.B(n_350),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.C(n_353),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_417),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_360),
.C(n_392),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_357),
.B(n_361),
.Y(n_511)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.C(n_388),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_362),
.B(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_364),
.B(n_389),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_369),
.C(n_379),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_369),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_367),
.B(n_445),
.C(n_447),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_380),
.B(n_427),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_381),
.B(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_381),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_381),
.A2(n_475),
.B1(n_476),
.B2(n_490),
.Y(n_489)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_415),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_415),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.C(n_413),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_394),
.B(n_509),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_397),
.B(n_413),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_402),
.C(n_411),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_440),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_403),
.B(n_412),
.Y(n_440)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_407),
.Y(n_406)
);

XOR2x1_ASAP7_75t_L g452 ( 
.A(n_408),
.B(n_453),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NAND3xp33_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.C(n_511),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_420),
.A2(n_506),
.B(n_510),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_455),
.B(n_505),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_441),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_422),
.B(n_441),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_438),
.B2(n_439),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_428),
.B2(n_429),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_425),
.B(n_429),
.C(n_438),
.Y(n_507)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

MAJx2_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.C(n_433),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_431),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_433),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

AO22x1_ASAP7_75t_SL g467 ( 
.A1(n_434),
.A2(n_435),
.B1(n_437),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_437),
.Y(n_468)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.C(n_451),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_470),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_452),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_447),
.Y(n_459)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

OAI21x1_ASAP7_75t_SL g455 ( 
.A1(n_456),
.A2(n_471),
.B(n_504),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_469),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_469),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.C(n_467),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_458),
.B(n_500),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_460),
.A2(n_461),
.B1(n_467),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_465),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_462),
.B(n_465),
.Y(n_479)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_467),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_492),
.Y(n_491)
);

AOI21x1_ASAP7_75t_SL g471 ( 
.A1(n_472),
.A2(n_498),
.B(n_503),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_473),
.A2(n_485),
.B(n_497),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_477),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_477),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_476),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_480),
.B2(n_481),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_491),
.B(n_496),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_489),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_489),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_502),
.Y(n_498)
);

NOR2x1_ASAP7_75t_SL g503 ( 
.A(n_499),
.B(n_502),
.Y(n_503)
);

NOR2xp67_ASAP7_75t_SL g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_507),
.B(n_508),
.Y(n_510)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);


endmodule