module fake_jpeg_12960_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_10),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_52),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_49),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_17),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_53),
.B(n_59),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_64),
.Y(n_107)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_28),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_62),
.Y(n_138)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_66),
.B(n_76),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_18),
.B(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_68),
.B(n_89),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_73),
.Y(n_106)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_78),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_79),
.Y(n_119)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_82),
.Y(n_130)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_87),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_85),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_31),
.B(n_15),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_91),
.Y(n_124)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_42),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_69),
.B1(n_67),
.B2(n_61),
.Y(n_96)
);

AO22x2_ASAP7_75t_L g172 ( 
.A1(n_96),
.A2(n_121),
.B1(n_140),
.B2(n_109),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_43),
.C(n_38),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_141),
.C(n_114),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_39),
.B1(n_29),
.B2(n_40),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_132),
.B1(n_117),
.B2(n_94),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_70),
.B1(n_88),
.B2(n_86),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_110),
.A2(n_117),
.B1(n_132),
.B2(n_144),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_58),
.A2(n_39),
.B1(n_29),
.B2(n_40),
.Y(n_117)
);

AO22x1_ASAP7_75t_SL g121 ( 
.A1(n_65),
.A2(n_43),
.B1(n_38),
.B2(n_41),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_141),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_56),
.B(n_42),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_143),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_55),
.B(n_41),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_128),
.B(n_131),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g129 ( 
.A1(n_60),
.A2(n_31),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_114),
.B(n_130),
.C(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_54),
.B(n_1),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_85),
.B1(n_82),
.B2(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_14),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_135),
.B(n_136),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_54),
.B(n_14),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_80),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_126),
.B1(n_97),
.B2(n_124),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_74),
.B(n_9),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_74),
.B(n_13),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_142),
.B(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_92),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_76),
.A2(n_58),
.B1(n_88),
.B2(n_86),
.Y(n_144)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_148),
.B1(n_113),
.B2(n_159),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_155),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_144),
.B1(n_133),
.B2(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_94),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_151),
.Y(n_214)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_103),
.B1(n_137),
.B2(n_100),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_169),
.Y(n_194)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_180),
.C(n_181),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_161),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_98),
.B(n_122),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_158),
.B(n_164),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_99),
.B(n_107),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_172),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_165),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_121),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_114),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_176),
.Y(n_206)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_95),
.A2(n_121),
.B1(n_105),
.B2(n_111),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_148),
.B1(n_146),
.B2(n_172),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_171),
.C(n_182),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_125),
.C(n_96),
.Y(n_171)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_127),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_177),
.Y(n_192)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_106),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_106),
.B(n_130),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_106),
.B(n_133),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_125),
.B(n_134),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_96),
.Y(n_182)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_113),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_183),
.Y(n_216)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_185),
.Y(n_212)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_113),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_214),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_199),
.Y(n_227)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_173),
.B(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_170),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_171),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_186),
.B(n_147),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_206),
.B(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_167),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_217),
.Y(n_235)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_165),
.A2(n_183),
.B(n_162),
.C(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_217),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_174),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_187),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_220),
.B(n_225),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_184),
.B(n_185),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_222),
.A2(n_224),
.B(n_209),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_145),
.C(n_150),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_230),
.C(n_232),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_189),
.B(n_199),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_197),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_240),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_214),
.C(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_239),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_189),
.B(n_192),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_SL g249 ( 
.A1(n_236),
.A2(n_225),
.A3(n_227),
.B1(n_234),
.B2(n_230),
.C1(n_238),
.C2(n_231),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_204),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_196),
.B1(n_191),
.B2(n_215),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_221),
.B1(n_219),
.B2(n_239),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_205),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_187),
.B(n_192),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_198),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_252),
.C(n_223),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_221),
.B1(n_219),
.B2(n_224),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_249),
.B(n_228),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_204),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_222),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

OAI322xp33_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_260),
.A3(n_262),
.B1(n_243),
.B2(n_265),
.C1(n_247),
.C2(n_241),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_227),
.B1(n_236),
.B2(n_228),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_241),
.B1(n_245),
.B2(n_244),
.Y(n_274)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_251),
.B(n_254),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_207),
.C(n_201),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_268),
.Y(n_273)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_207),
.C(n_201),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_216),
.C(n_212),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_269),
.A2(n_216),
.B(n_188),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_251),
.B(n_256),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_277),
.B(n_276),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_242),
.B1(n_246),
.B2(n_255),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_279),
.B1(n_257),
.B2(n_266),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_263),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_278),
.A2(n_267),
.B1(n_269),
.B2(n_260),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_286),
.B1(n_273),
.B2(n_277),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_273),
.C(n_268),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_290),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_278),
.B1(n_271),
.B2(n_279),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_280),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g292 ( 
.A1(n_288),
.A2(n_272),
.B(n_283),
.C(n_280),
.Y(n_292)
);

OAI22x1_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_287),
.B1(n_209),
.B2(n_255),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_289),
.Y(n_296)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_290),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_293),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_211),
.C(n_226),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_299),
.A2(n_210),
.B(n_226),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_300),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_210),
.Y(n_303)
);


endmodule