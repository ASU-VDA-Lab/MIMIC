module fake_jpeg_25892_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_9),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_20),
.B1(n_24),
.B2(n_23),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_17),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_37),
.B(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_40),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_22),
.B1(n_16),
.B2(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_37),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_32),
.B1(n_19),
.B2(n_23),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_32),
.B1(n_19),
.B2(n_24),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_36),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_64),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_61),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_38),
.B1(n_35),
.B2(n_31),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_84),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_35),
.C(n_36),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_87),
.C(n_36),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_66),
.Y(n_107)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_36),
.B1(n_28),
.B2(n_31),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_86),
.B1(n_59),
.B2(n_58),
.Y(n_106)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_17),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_86),
.B(n_63),
.C(n_82),
.Y(n_108)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_72),
.Y(n_109)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_27),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_85),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_88),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_21),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_51),
.B(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_92),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_49),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_114),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_56),
.B1(n_52),
.B2(n_21),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_74),
.B1(n_53),
.B2(n_72),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_108),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_56),
.C(n_25),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_74),
.C(n_53),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_68),
.B1(n_78),
.B2(n_77),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_39),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_102),
.Y(n_125)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_39),
.Y(n_114)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_79),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_123),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_94),
.B1(n_106),
.B2(n_114),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_118),
.A2(n_119),
.B1(n_134),
.B2(n_113),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_59),
.B1(n_86),
.B2(n_85),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_62),
.B1(n_75),
.B2(n_61),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_120),
.A2(n_127),
.B1(n_110),
.B2(n_93),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_60),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_138),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_126),
.B(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_84),
.B1(n_69),
.B2(n_73),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_137),
.B1(n_126),
.B2(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_132),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_0),
.B(n_1),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_0),
.B(n_1),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_90),
.C(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_89),
.B(n_9),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_39),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_145),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_29),
.B1(n_53),
.B2(n_8),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_53),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_53),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_2),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_7),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_90),
.B(n_100),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_2),
.B(n_3),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_149),
.A2(n_161),
.B(n_170),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_101),
.B(n_97),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_165),
.C(n_167),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_131),
.C(n_10),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_116),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_159),
.Y(n_181)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_109),
.B(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_115),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_115),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_173),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_53),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_168),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_93),
.B1(n_110),
.B2(n_2),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_176),
.B1(n_11),
.B2(n_14),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_10),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_120),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_7),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_140),
.B(n_132),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_178),
.A2(n_183),
.B(n_196),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_184),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_176),
.C(n_149),
.Y(n_219)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_186),
.B(n_190),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_195),
.B1(n_197),
.B2(n_202),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_6),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_6),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_15),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_166),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_147),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_165),
.B1(n_175),
.B2(n_159),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_163),
.B1(n_148),
.B2(n_152),
.Y(n_215)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_213),
.Y(n_226)
);

XOR2x2_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_161),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_208),
.B(n_212),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_156),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_216),
.B1(n_220),
.B2(n_199),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_169),
.B1(n_150),
.B2(n_146),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_201),
.B(n_172),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_203),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_219),
.B(n_223),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_150),
.B1(n_174),
.B2(n_154),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_177),
.C(n_162),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_224),
.C(n_182),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_148),
.C(n_170),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_198),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_188),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_236),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_231),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_185),
.B1(n_204),
.B2(n_184),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_213),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_233),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_234),
.A2(n_240),
.B(n_205),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_178),
.B(n_183),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_235),
.A2(n_218),
.B(n_234),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_206),
.B(n_166),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_239),
.C(n_241),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_192),
.Y(n_239)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_181),
.B(n_187),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_192),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_224),
.C(n_214),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_241),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_210),
.Y(n_255)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_210),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_235),
.A2(n_197),
.B1(n_195),
.B2(n_202),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_252),
.B1(n_254),
.B2(n_251),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_250),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_158),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_248),
.B1(n_242),
.B2(n_180),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_242),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_239),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_266),
.B(n_268),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_219),
.B(n_209),
.C(n_181),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_245),
.B1(n_253),
.B2(n_187),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_275),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_277),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_180),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_248),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_247),
.C(n_4),
.Y(n_285)
);

A2O1A1O1Ixp25_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_247),
.B(n_217),
.C(n_229),
.D(n_225),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_265),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_285),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_262),
.B(n_267),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_281),
.B(n_279),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_289),
.C(n_272),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_280),
.A2(n_276),
.B(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_273),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_287),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_293),
.Y(n_294)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_3),
.A3(n_5),
.B1(n_284),
.B2(n_292),
.C(n_293),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_3),
.Y(n_297)
);


endmodule