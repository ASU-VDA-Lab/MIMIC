module fake_ibex_1295_n_1403 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1403);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1403;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_262;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_291;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_485;
wire n_1315;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_326;
wire n_270;
wire n_1340;
wire n_259;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1374;
wire n_792;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g259 ( 
.A(n_164),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_53),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_16),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_209),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_L g265 ( 
.A(n_193),
.B(n_251),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_220),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_73),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_234),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_254),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_179),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_175),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_L g273 ( 
.A(n_139),
.B(n_190),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_32),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_163),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_107),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_2),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_18),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_98),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_116),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_2),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_194),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_118),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_151),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_198),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_0),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_96),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_130),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_221),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_225),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_205),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_94),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_25),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_42),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_236),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_233),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_10),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_22),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_157),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_200),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_17),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_74),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_44),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_78),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_136),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_162),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_155),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_214),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_114),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_100),
.B(n_189),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_186),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_166),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_102),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_207),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_156),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_97),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_93),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_140),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_77),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_132),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_174),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_258),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_244),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_56),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_222),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_101),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_108),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_51),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_142),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_228),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_64),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_145),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_23),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_181),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_182),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_7),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_226),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_248),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_253),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_224),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_148),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_26),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_159),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_229),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_201),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_238),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_57),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_143),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_243),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_37),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_147),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_144),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_231),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_170),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_69),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_252),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_223),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_196),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_111),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_150),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_138),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_216),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_79),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_230),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_137),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_87),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_83),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_203),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_199),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_68),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_213),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_89),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_255),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_34),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_168),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_239),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_218),
.B(n_217),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_232),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_23),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_152),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_6),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_73),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_135),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_46),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_184),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_59),
.Y(n_389)
);

CKINVDCx11_ASAP7_75t_R g390 ( 
.A(n_211),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_33),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_129),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_68),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_227),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_15),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_188),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_169),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_195),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_158),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_154),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_8),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_22),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_63),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_160),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_192),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_134),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_119),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_15),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_165),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_90),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_3),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_167),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_161),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_87),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_131),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_146),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_123),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_245),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_149),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_67),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_20),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_113),
.B(n_46),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_187),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_115),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_183),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_21),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_75),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_180),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_29),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_112),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_235),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_57),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_64),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_17),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_202),
.Y(n_435)
);

BUFx5_ASAP7_75t_L g436 ( 
.A(n_208),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_72),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_83),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_197),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_67),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_178),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_24),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_133),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_99),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_141),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_219),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_103),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_61),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_55),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_237),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_206),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_176),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_105),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_246),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_58),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_177),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_266),
.Y(n_457)
);

BUFx8_ASAP7_75t_SL g458 ( 
.A(n_353),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_314),
.B(n_1),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_318),
.B(n_1),
.Y(n_460)
);

BUFx12f_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_290),
.Y(n_462)
);

INVxp33_ASAP7_75t_SL g463 ( 
.A(n_263),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_266),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_266),
.Y(n_465)
);

OA21x2_ASAP7_75t_L g466 ( 
.A1(n_262),
.A2(n_104),
.B(n_95),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_290),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_R g468 ( 
.A1(n_261),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_468)
);

OA21x2_ASAP7_75t_L g469 ( 
.A1(n_262),
.A2(n_109),
.B(n_106),
.Y(n_469)
);

OA21x2_ASAP7_75t_L g470 ( 
.A1(n_335),
.A2(n_117),
.B(n_110),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_330),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_353),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_472)
);

CKINVDCx11_ASAP7_75t_R g473 ( 
.A(n_358),
.Y(n_473)
);

BUFx8_ASAP7_75t_SL g474 ( 
.A(n_358),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_384),
.B(n_7),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_427),
.B(n_9),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_456),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_327),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_296),
.Y(n_479)
);

CKINVDCx6p67_ASAP7_75t_R g480 ( 
.A(n_390),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_266),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_296),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_437),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_284),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_407),
.B(n_9),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g486 ( 
.A1(n_335),
.A2(n_357),
.B(n_346),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_437),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_296),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_296),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_346),
.A2(n_121),
.B(n_120),
.Y(n_490)
);

INVx6_ASAP7_75t_L g491 ( 
.A(n_308),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_308),
.Y(n_492)
);

BUFx8_ASAP7_75t_SL g493 ( 
.A(n_366),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_431),
.B(n_454),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_367),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_294),
.B(n_10),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_271),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_306),
.B(n_382),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_367),
.Y(n_499)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_308),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_294),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_275),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_336),
.Y(n_503)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_365),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_334),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_334),
.B(n_11),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_271),
.Y(n_507)
);

BUFx8_ASAP7_75t_SL g508 ( 
.A(n_366),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_414),
.B(n_11),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_344),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_271),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_296),
.B(n_12),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_296),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_292),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_296),
.B(n_14),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_452),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_292),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_292),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_448),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_292),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_412),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_357),
.B(n_19),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_448),
.B(n_20),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_267),
.Y(n_524)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_412),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_276),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_278),
.B(n_27),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_301),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_436),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_304),
.B(n_27),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_412),
.Y(n_531)
);

BUFx8_ASAP7_75t_L g532 ( 
.A(n_436),
.Y(n_532)
);

BUFx12f_ASAP7_75t_L g533 ( 
.A(n_264),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_305),
.B(n_28),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_410),
.Y(n_535)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_361),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_320),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_322),
.B(n_28),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_361),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_260),
.Y(n_540)
);

OA21x2_ASAP7_75t_L g541 ( 
.A1(n_372),
.A2(n_409),
.B(n_399),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_276),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_372),
.B(n_399),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_436),
.Y(n_544)
);

BUFx12f_ASAP7_75t_L g545 ( 
.A(n_268),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_345),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_338),
.B(n_30),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_409),
.A2(n_124),
.B(n_122),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_280),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_396),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_436),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_410),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_350),
.B(n_34),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_413),
.A2(n_126),
.B(n_125),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_396),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_269),
.Y(n_557)
);

BUFx8_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_338),
.B(n_35),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_361),
.Y(n_560)
);

OAI22x1_ASAP7_75t_SL g561 ( 
.A1(n_389),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_436),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_413),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_361),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_410),
.Y(n_565)
);

INVx8_ASAP7_75t_L g566 ( 
.A(n_500),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_496),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_L g568 ( 
.A(n_548),
.B(n_313),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_479),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_532),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_495),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_532),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_482),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_492),
.B(n_270),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_482),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_488),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_492),
.B(n_347),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_488),
.Y(n_579)
);

NOR2x1p5_ASAP7_75t_L g580 ( 
.A(n_480),
.B(n_370),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_489),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_489),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_513),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_478),
.B(n_347),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_513),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_496),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_506),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_506),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_457),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_486),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_463),
.A2(n_356),
.B1(n_378),
.B2(n_280),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_461),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_509),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_486),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_491),
.B(n_259),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_523),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_529),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_540),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_541),
.Y(n_599)
);

AO21x2_ASAP7_75t_L g600 ( 
.A1(n_555),
.A2(n_274),
.B(n_272),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_529),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_544),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_544),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_462),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_547),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_495),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_487),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_487),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_552),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_462),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_552),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_562),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_562),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_538),
.Y(n_614)
);

AOI21x1_ASAP7_75t_L g615 ( 
.A1(n_512),
.A2(n_451),
.B(n_277),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_457),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_457),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_521),
.B(n_283),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_464),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_462),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_464),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_558),
.Y(n_622)
);

AND3x2_ASAP7_75t_L g623 ( 
.A(n_503),
.B(n_395),
.C(n_391),
.Y(n_623)
);

AND3x2_ASAP7_75t_L g624 ( 
.A(n_502),
.B(n_411),
.C(n_402),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_465),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_465),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_465),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_481),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_531),
.B(n_279),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_499),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_462),
.Y(n_631)
);

INVxp33_ASAP7_75t_SL g632 ( 
.A(n_516),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_461),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_558),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_499),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_483),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_467),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_498),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_557),
.B(n_282),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_497),
.Y(n_640)
);

AO21x2_ASAP7_75t_L g641 ( 
.A1(n_515),
.A2(n_285),
.B(n_281),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_504),
.B(n_288),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_557),
.B(n_286),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_504),
.B(n_287),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_504),
.B(n_433),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_559),
.B(n_451),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_525),
.B(n_298),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_477),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_475),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_525),
.Y(n_650)
);

CKINVDCx6p67_ASAP7_75t_R g651 ( 
.A(n_533),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_525),
.B(n_302),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_471),
.B(n_463),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_563),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_497),
.Y(n_655)
);

BUFx6f_ASAP7_75t_SL g656 ( 
.A(n_551),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_494),
.B(n_295),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_507),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_556),
.Y(n_659)
);

AND3x2_ASAP7_75t_L g660 ( 
.A(n_468),
.B(n_442),
.C(n_438),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_516),
.B(n_524),
.Y(n_661)
);

NOR2x1p5_ASAP7_75t_L g662 ( 
.A(n_484),
.B(n_533),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_507),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_485),
.B(n_289),
.Y(n_664)
);

AOI21x1_ASAP7_75t_L g665 ( 
.A1(n_466),
.A2(n_315),
.B(n_309),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_507),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_563),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_511),
.Y(n_668)
);

INVxp33_ASAP7_75t_L g669 ( 
.A(n_459),
.Y(n_669)
);

AOI21x1_ASAP7_75t_L g670 ( 
.A1(n_466),
.A2(n_321),
.B(n_316),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_556),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_528),
.Y(n_672)
);

OAI22xp33_ASAP7_75t_SL g673 ( 
.A1(n_526),
.A2(n_307),
.B1(n_331),
.B2(n_300),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_458),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_537),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_535),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_546),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_545),
.B(n_323),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_501),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_511),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_545),
.B(n_332),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_505),
.B(n_455),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_514),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_514),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_519),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_527),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_543),
.B(n_291),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_514),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_514),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_535),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_530),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_534),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_553),
.Y(n_693)
);

AO22x2_ASAP7_75t_L g694 ( 
.A1(n_476),
.A2(n_342),
.B1(n_343),
.B2(n_341),
.Y(n_694)
);

AND3x2_ASAP7_75t_L g695 ( 
.A(n_459),
.B(n_354),
.C(n_348),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_510),
.A2(n_408),
.B1(n_434),
.B2(n_389),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_517),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_517),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_554),
.B(n_293),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_543),
.B(n_339),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_522),
.B(n_297),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_522),
.B(n_299),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_517),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_553),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_460),
.B(n_369),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_517),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_565),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_518),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_565),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_460),
.B(n_303),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_458),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_565),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_520),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_686),
.B(n_691),
.Y(n_714)
);

NAND2x1_ASAP7_75t_L g715 ( 
.A(n_567),
.B(n_466),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_692),
.B(n_469),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_571),
.B(n_310),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_672),
.B(n_469),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_653),
.A2(n_356),
.B1(n_383),
.B2(n_378),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_694),
.A2(n_426),
.B1(n_410),
.B2(n_388),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_571),
.B(n_311),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_672),
.B(n_584),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_584),
.B(n_469),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_641),
.B(n_470),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_638),
.B(n_432),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_675),
.A2(n_363),
.B(n_371),
.C(n_360),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_641),
.B(n_470),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_694),
.A2(n_550),
.B1(n_542),
.B2(n_388),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_641),
.B(n_470),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_607),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_598),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_677),
.B(n_490),
.Y(n_732)
);

NOR2xp67_ASAP7_75t_L g733 ( 
.A(n_592),
.B(n_536),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_573),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_608),
.Y(n_735)
);

INVx8_ASAP7_75t_L g736 ( 
.A(n_566),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_657),
.B(n_700),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_573),
.B(n_312),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_700),
.B(n_317),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_629),
.B(n_444),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_659),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_649),
.B(n_319),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_622),
.B(n_324),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_578),
.B(n_325),
.Y(n_744)
);

NOR3xp33_ASAP7_75t_L g745 ( 
.A(n_696),
.B(n_473),
.C(n_472),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_671),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_694),
.A2(n_426),
.B1(n_397),
.B2(n_419),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_639),
.B(n_326),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_587),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_633),
.B(n_561),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_669),
.B(n_328),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_669),
.B(n_329),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_614),
.B(n_333),
.Y(n_753)
);

INVxp33_ASAP7_75t_L g754 ( 
.A(n_591),
.Y(n_754)
);

INVxp33_ASAP7_75t_L g755 ( 
.A(n_661),
.Y(n_755)
);

AO221x1_ASAP7_75t_L g756 ( 
.A1(n_694),
.A2(n_473),
.B1(n_474),
.B2(n_493),
.C(n_508),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_622),
.B(n_337),
.Y(n_757)
);

AOI221xp5_ASAP7_75t_L g758 ( 
.A1(n_673),
.A2(n_440),
.B1(n_373),
.B2(n_375),
.C(n_377),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_596),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_572),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_586),
.B(n_340),
.Y(n_761)
);

AND2x2_ASAP7_75t_SL g762 ( 
.A(n_633),
.B(n_474),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_568),
.B(n_387),
.C(n_385),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_580),
.B(n_408),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_651),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_588),
.B(n_349),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_645),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_644),
.B(n_351),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_650),
.B(n_352),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_L g770 ( 
.A(n_592),
.B(n_536),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_593),
.B(n_355),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_596),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_572),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_650),
.B(n_359),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_710),
.B(n_362),
.Y(n_775)
);

BUFx5_ASAP7_75t_L g776 ( 
.A(n_597),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_637),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_595),
.B(n_364),
.Y(n_778)
);

INVxp33_ASAP7_75t_L g779 ( 
.A(n_705),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_606),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_606),
.B(n_368),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_575),
.B(n_374),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_630),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_590),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_643),
.B(n_376),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_642),
.B(n_381),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_630),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_647),
.B(n_652),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_568),
.B(n_386),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_594),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_597),
.B(n_490),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_566),
.B(n_400),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_635),
.B(n_405),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_634),
.B(n_393),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_687),
.B(n_415),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_701),
.B(n_416),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_674),
.B(n_403),
.C(n_401),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_676),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_SL g799 ( 
.A(n_656),
.B(n_383),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_651),
.B(n_420),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_678),
.B(n_423),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_646),
.A2(n_681),
.B1(n_699),
.B2(n_632),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_648),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_682),
.B(n_421),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_702),
.B(n_428),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_648),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_646),
.B(n_430),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_679),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_699),
.B(n_664),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_632),
.A2(n_419),
.B1(n_435),
.B2(n_397),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_636),
.B(n_441),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_685),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_654),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_667),
.Y(n_814)
);

BUFx6f_ASAP7_75t_SL g815 ( 
.A(n_711),
.Y(n_815)
);

BUFx5_ASAP7_75t_L g816 ( 
.A(n_602),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_603),
.B(n_429),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_603),
.B(n_490),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_599),
.B(n_549),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_690),
.Y(n_820)
);

CKINVDCx11_ASAP7_75t_R g821 ( 
.A(n_662),
.Y(n_821)
);

NOR2x1p5_ASAP7_75t_L g822 ( 
.A(n_660),
.B(n_493),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_656),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_618),
.B(n_379),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_624),
.B(n_449),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_615),
.B(n_392),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_574),
.B(n_394),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_574),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_576),
.B(n_398),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_695),
.B(n_404),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_576),
.B(n_406),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_604),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_601),
.B(n_418),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_704),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_656),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_605),
.B(n_424),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_605),
.B(n_425),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_610),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_704),
.B(n_38),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_623),
.B(n_434),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_609),
.B(n_439),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_620),
.Y(n_842)
);

OAI22xp33_ASAP7_75t_L g843 ( 
.A1(n_631),
.A2(n_435),
.B1(n_445),
.B2(n_426),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_631),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_693),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_611),
.B(n_443),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_612),
.B(n_446),
.Y(n_847)
);

NOR2xp67_ASAP7_75t_L g848 ( 
.A(n_693),
.B(n_39),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_612),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_613),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_724),
.A2(n_670),
.B(n_665),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_714),
.B(n_600),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_819),
.A2(n_600),
.B(n_577),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_819),
.A2(n_718),
.B(n_716),
.Y(n_854)
);

OAI21xp33_ASAP7_75t_L g855 ( 
.A1(n_779),
.A2(n_577),
.B(n_570),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_765),
.Y(n_856)
);

O2A1O1Ixp5_ASAP7_75t_L g857 ( 
.A1(n_715),
.A2(n_670),
.B(n_665),
.C(n_579),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_722),
.B(n_600),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_716),
.A2(n_582),
.B(n_581),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_731),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_723),
.A2(n_582),
.B(n_581),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_722),
.B(n_737),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_723),
.A2(n_585),
.B(n_583),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_804),
.B(n_426),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_720),
.A2(n_828),
.B1(n_747),
.B2(n_843),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_725),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_732),
.A2(n_713),
.B(n_450),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_736),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_732),
.A2(n_713),
.B(n_453),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_755),
.B(n_508),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_808),
.B(n_812),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_724),
.A2(n_447),
.B(n_707),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_749),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_727),
.A2(n_273),
.B(n_265),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_729),
.A2(n_380),
.B(n_422),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_791),
.A2(n_712),
.B(n_709),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_759),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_751),
.B(n_417),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_752),
.B(n_40),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_791),
.A2(n_712),
.B(n_617),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_772),
.Y(n_881)
);

NOR2x2_ASAP7_75t_L g882 ( 
.A(n_764),
.B(n_41),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_736),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_818),
.A2(n_617),
.B(n_616),
.Y(n_884)
);

OR2x2_ASAP7_75t_SL g885 ( 
.A(n_762),
.B(n_42),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_818),
.A2(n_619),
.B(n_616),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_813),
.A2(n_520),
.B(n_539),
.C(n_560),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_754),
.B(n_43),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_767),
.B(n_45),
.Y(n_889)
);

AO21x1_ASAP7_75t_L g890 ( 
.A1(n_826),
.A2(n_626),
.B(n_625),
.Y(n_890)
);

NOR2x1_ASAP7_75t_L g891 ( 
.A(n_763),
.B(n_800),
.Y(n_891)
);

AND2x2_ASAP7_75t_SL g892 ( 
.A(n_799),
.B(n_47),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_742),
.B(n_48),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_740),
.B(n_48),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_739),
.B(n_49),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_730),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_809),
.A2(n_628),
.B(n_627),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_817),
.B(n_50),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_734),
.B(n_50),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_776),
.B(n_52),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_735),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_816),
.B(n_52),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_816),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_726),
.A2(n_849),
.B(n_850),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_802),
.B(n_794),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_827),
.A2(n_831),
.B(n_829),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_816),
.B(n_54),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_788),
.B(n_55),
.Y(n_908)
);

BUFx4f_ASAP7_75t_L g909 ( 
.A(n_750),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_810),
.Y(n_910)
);

CKINVDCx8_ASAP7_75t_R g911 ( 
.A(n_750),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_814),
.A2(n_539),
.B(n_560),
.C(n_564),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_801),
.B(n_56),
.Y(n_913)
);

BUFx12f_ASAP7_75t_L g914 ( 
.A(n_821),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_777),
.B(n_59),
.Y(n_915)
);

AO21x1_ASAP7_75t_L g916 ( 
.A1(n_829),
.A2(n_655),
.B(n_640),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_717),
.B(n_60),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_764),
.B(n_60),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_721),
.B(n_61),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_764),
.B(n_62),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_784),
.A2(n_658),
.B(n_655),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_790),
.A2(n_666),
.B(n_663),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_789),
.B(n_748),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_833),
.A2(n_668),
.B(n_666),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_790),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_811),
.B(n_753),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_743),
.B(n_757),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_L g928 ( 
.A(n_790),
.B(n_569),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_823),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_741),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_761),
.B(n_63),
.Y(n_931)
);

OAI21xp33_ASAP7_75t_L g932 ( 
.A1(n_728),
.A2(n_684),
.B(n_683),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_758),
.A2(n_689),
.B1(n_706),
.B2(n_703),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_745),
.A2(n_688),
.B(n_689),
.C(n_697),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_768),
.B(n_65),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_807),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_936)
);

BUFx4f_ASAP7_75t_L g937 ( 
.A(n_750),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_744),
.B(n_569),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_775),
.B(n_66),
.Y(n_939)
);

AOI21xp33_ASAP7_75t_L g940 ( 
.A1(n_796),
.A2(n_70),
.B(n_71),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_792),
.B(n_589),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_835),
.B(n_71),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_766),
.B(n_771),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_832),
.A2(n_708),
.B(n_698),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_836),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_746),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_760),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_781),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_805),
.B(n_76),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_773),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_795),
.B(n_77),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_836),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_837),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_953)
);

OAI21xp33_ASAP7_75t_L g954 ( 
.A1(n_837),
.A2(n_708),
.B(n_698),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_733),
.B(n_81),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_785),
.B(n_84),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_838),
.A2(n_708),
.B(n_698),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_844),
.A2(n_680),
.B(n_621),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_841),
.B(n_85),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_803),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_806),
.Y(n_961)
);

NOR3xp33_ASAP7_75t_L g962 ( 
.A(n_840),
.B(n_86),
.C(n_88),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_847),
.B(n_89),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_847),
.A2(n_680),
.B1(n_621),
.B2(n_589),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_830),
.B(n_90),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_845),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_782),
.B(n_91),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_825),
.Y(n_968)
);

AO21x2_ASAP7_75t_L g969 ( 
.A1(n_848),
.A2(n_839),
.B(n_846),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_780),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_842),
.A2(n_820),
.B(n_798),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_797),
.B(n_91),
.Y(n_972)
);

CKINVDCx10_ASAP7_75t_R g973 ( 
.A(n_815),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_738),
.B(n_92),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_783),
.Y(n_975)
);

NOR2x1_ASAP7_75t_L g976 ( 
.A(n_868),
.B(n_822),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_854),
.A2(n_834),
.B(n_787),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_868),
.B(n_770),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_SL g979 ( 
.A1(n_862),
.A2(n_778),
.B(n_786),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_901),
.Y(n_980)
);

AND3x4_ASAP7_75t_L g981 ( 
.A(n_973),
.B(n_756),
.C(n_815),
.Y(n_981)
);

NOR2x1_ASAP7_75t_L g982 ( 
.A(n_929),
.B(n_793),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_906),
.A2(n_769),
.B1(n_774),
.B2(n_824),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_883),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_851),
.A2(n_127),
.B(n_128),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_871),
.Y(n_986)
);

AND3x4_ASAP7_75t_L g987 ( 
.A(n_962),
.B(n_911),
.C(n_909),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_966),
.Y(n_988)
);

AOI21xp33_ASAP7_75t_L g989 ( 
.A1(n_879),
.A2(n_894),
.B(n_865),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_860),
.B(n_153),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_909),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_892),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_910),
.B(n_204),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_861),
.A2(n_212),
.B(n_215),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_876),
.A2(n_859),
.B(n_863),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_864),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_915),
.Y(n_997)
);

AO31x2_ASAP7_75t_L g998 ( 
.A1(n_890),
.A2(n_240),
.A3(n_241),
.B(n_242),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_891),
.B(n_247),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_968),
.B(n_256),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_867),
.A2(n_869),
.B(n_872),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_927),
.B(n_899),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_899),
.B(n_943),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_880),
.A2(n_886),
.B(n_884),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_964),
.A2(n_875),
.B(n_938),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_856),
.B(n_914),
.Y(n_1006)
);

AO21x1_ASAP7_75t_L g1007 ( 
.A1(n_964),
.A2(n_902),
.B(n_900),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_944),
.A2(n_958),
.B(n_957),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_942),
.B(n_908),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_932),
.A2(n_904),
.B(n_959),
.C(n_963),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_942),
.B(n_895),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_928),
.A2(n_971),
.B(n_878),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_918),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_SL g1014 ( 
.A1(n_925),
.A2(n_907),
.B(n_903),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_924),
.A2(n_897),
.B(n_941),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_SL g1016 ( 
.A1(n_904),
.A2(n_893),
.B(n_898),
.Y(n_1016)
);

AOI21xp33_ASAP7_75t_L g1017 ( 
.A1(n_935),
.A2(n_951),
.B(n_949),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_870),
.B(n_948),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_955),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_921),
.A2(n_922),
.B(n_954),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_972),
.B(n_873),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_889),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_877),
.B(n_881),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_920),
.B(n_937),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_960),
.A2(n_961),
.B(n_950),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_SL g1026 ( 
.A1(n_974),
.A2(n_939),
.B(n_967),
.Y(n_1026)
);

OA21x2_ASAP7_75t_L g1027 ( 
.A1(n_887),
.A2(n_912),
.B(n_956),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_945),
.Y(n_1028)
);

AO31x2_ASAP7_75t_L g1029 ( 
.A1(n_952),
.A2(n_953),
.A3(n_936),
.B(n_913),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_882),
.Y(n_1030)
);

AO31x2_ASAP7_75t_L g1031 ( 
.A1(n_931),
.A2(n_919),
.A3(n_917),
.B(n_946),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_965),
.B(n_855),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_930),
.A2(n_933),
.B(n_940),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_947),
.B(n_970),
.Y(n_1034)
);

AND3x1_ASAP7_75t_SL g1035 ( 
.A(n_885),
.B(n_969),
.C(n_947),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_970),
.B(n_975),
.Y(n_1036)
);

OR2x6_ASAP7_75t_L g1037 ( 
.A(n_970),
.B(n_975),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_906),
.A2(n_923),
.B(n_926),
.C(n_905),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_883),
.B(n_868),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_910),
.A2(n_754),
.B1(n_745),
.B2(n_728),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_854),
.A2(n_819),
.B(n_718),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_854),
.A2(n_819),
.B(n_718),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_854),
.A2(n_819),
.B(n_718),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_862),
.B(n_714),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_854),
.A2(n_819),
.B(n_718),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_866),
.B(n_754),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_862),
.B(n_714),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_875),
.B(n_874),
.C(n_888),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_SL g1049 ( 
.A1(n_906),
.A2(n_868),
.B(n_871),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_854),
.A2(n_819),
.B(n_718),
.Y(n_1050)
);

OAI21xp33_ASAP7_75t_L g1051 ( 
.A1(n_862),
.A2(n_755),
.B(n_669),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_854),
.A2(n_853),
.B(n_852),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_862),
.B(n_714),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_866),
.B(n_779),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_862),
.B(n_714),
.Y(n_1055)
);

BUFx4f_ASAP7_75t_L g1056 ( 
.A(n_883),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_866),
.B(n_779),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_SL g1058 ( 
.A1(n_906),
.A2(n_868),
.B(n_871),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_866),
.B(n_754),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_860),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_854),
.A2(n_853),
.B(n_852),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_860),
.Y(n_1062)
);

AOI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_866),
.A2(n_755),
.B(n_779),
.Y(n_1063)
);

CKINVDCx6p67_ASAP7_75t_R g1064 ( 
.A(n_973),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_883),
.B(n_868),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_854),
.A2(n_853),
.B(n_852),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_866),
.B(n_779),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_906),
.A2(n_923),
.B(n_926),
.C(n_905),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_SL g1069 ( 
.A1(n_906),
.A2(n_868),
.B(n_871),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_896),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_862),
.B(n_714),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_862),
.B(n_714),
.Y(n_1072)
);

AND3x2_ASAP7_75t_L g1073 ( 
.A(n_860),
.B(n_674),
.C(n_799),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_868),
.B(n_714),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_883),
.B(n_868),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_860),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_883),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_866),
.B(n_779),
.Y(n_1078)
);

AO21x1_ASAP7_75t_L g1079 ( 
.A1(n_858),
.A2(n_874),
.B(n_852),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_896),
.Y(n_1080)
);

AOI21xp33_ASAP7_75t_L g1081 ( 
.A1(n_934),
.A2(n_879),
.B(n_858),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_862),
.B(n_714),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_854),
.A2(n_819),
.B(n_718),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_866),
.B(n_779),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_862),
.B(n_714),
.Y(n_1085)
);

AOI21xp33_ASAP7_75t_L g1086 ( 
.A1(n_934),
.A2(n_879),
.B(n_858),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_866),
.B(n_754),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_862),
.B(n_714),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_862),
.B(n_714),
.Y(n_1089)
);

OA22x2_ASAP7_75t_L g1090 ( 
.A1(n_910),
.A2(n_810),
.B1(n_591),
.B2(n_719),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_866),
.B(n_779),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_862),
.B(n_714),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_866),
.B(n_779),
.Y(n_1093)
);

OA21x2_ASAP7_75t_L g1094 ( 
.A1(n_851),
.A2(n_853),
.B(n_857),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_862),
.B(n_714),
.Y(n_1095)
);

AND3x4_ASAP7_75t_L g1096 ( 
.A(n_973),
.B(n_745),
.C(n_765),
.Y(n_1096)
);

NAND2x1p5_ASAP7_75t_L g1097 ( 
.A(n_868),
.B(n_883),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1090),
.A2(n_1040),
.B1(n_1028),
.B2(n_1030),
.Y(n_1098)
);

INVxp67_ASAP7_75t_SL g1099 ( 
.A(n_1052),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1044),
.B(n_1047),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_1062),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1038),
.A2(n_1068),
.B(n_1061),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1053),
.B(n_1055),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1071),
.Y(n_1104)
);

AO21x2_ASAP7_75t_L g1105 ( 
.A1(n_1066),
.A2(n_1007),
.B(n_1016),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1048),
.A2(n_987),
.B1(n_986),
.B2(n_1051),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1072),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1082),
.A2(n_1085),
.B1(n_1089),
.B2(n_1088),
.Y(n_1108)
);

OR2x6_ASAP7_75t_L g1109 ( 
.A(n_1092),
.B(n_1095),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_980),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1041),
.A2(n_1043),
.B(n_1042),
.Y(n_1111)
);

OAI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_992),
.A2(n_1019),
.B1(n_1009),
.B2(n_1011),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_1069),
.A2(n_1086),
.B(n_1081),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_1054),
.B(n_1057),
.Y(n_1114)
);

BUFx8_ASAP7_75t_SL g1115 ( 
.A(n_1006),
.Y(n_1115)
);

BUFx10_ASAP7_75t_L g1116 ( 
.A(n_1006),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1020),
.A2(n_1004),
.B(n_995),
.Y(n_1117)
);

CKINVDCx6p67_ASAP7_75t_R g1118 ( 
.A(n_1064),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1004),
.A2(n_1008),
.B(n_1015),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_1056),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_1076),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_991),
.B(n_976),
.Y(n_1122)
);

AO21x2_ASAP7_75t_L g1123 ( 
.A1(n_1048),
.A2(n_989),
.B(n_1005),
.Y(n_1123)
);

OAI22x1_ASAP7_75t_L g1124 ( 
.A1(n_981),
.A2(n_992),
.B1(n_1096),
.B2(n_991),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_984),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1045),
.A2(n_1083),
.B(n_1050),
.Y(n_1126)
);

NAND2x1p5_ASAP7_75t_L g1127 ( 
.A(n_1056),
.B(n_1077),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_SL g1128 ( 
.A1(n_985),
.A2(n_1026),
.B(n_994),
.Y(n_1128)
);

BUFx2_ASAP7_75t_SL g1129 ( 
.A(n_1077),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1046),
.A2(n_1059),
.B1(n_1087),
.B2(n_1051),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1097),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1067),
.B(n_1078),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1017),
.A2(n_1001),
.B(n_1012),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_1097),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1070),
.B(n_1080),
.Y(n_1135)
);

AO21x2_ASAP7_75t_L g1136 ( 
.A1(n_1017),
.A2(n_1033),
.B(n_1001),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1094),
.A2(n_1032),
.B(n_1033),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1025),
.A2(n_977),
.B(n_1014),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_988),
.Y(n_1139)
);

AOI21x1_ASAP7_75t_L g1140 ( 
.A1(n_999),
.A2(n_1034),
.B(n_1027),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_1006),
.Y(n_1141)
);

BUFx2_ASAP7_75t_R g1142 ( 
.A(n_1003),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1023),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1021),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_979),
.B(n_997),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_979),
.A2(n_983),
.B(n_996),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1022),
.B(n_1002),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1060),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_978),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_993),
.A2(n_1036),
.B(n_1000),
.Y(n_1150)
);

INVx5_ASAP7_75t_L g1151 ( 
.A(n_1037),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1029),
.B(n_1031),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_990),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1039),
.A2(n_1065),
.B(n_1075),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1084),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1013),
.B(n_1063),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1091),
.B(n_1093),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_998),
.A2(n_982),
.B(n_1035),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_978),
.A2(n_1018),
.B1(n_1024),
.B2(n_1029),
.Y(n_1159)
);

OA21x2_ASAP7_75t_L g1160 ( 
.A1(n_1031),
.A2(n_1029),
.B(n_1073),
.Y(n_1160)
);

OR3x4_ASAP7_75t_SL g1161 ( 
.A(n_1031),
.B(n_981),
.C(n_973),
.Y(n_1161)
);

INVx5_ASAP7_75t_L g1162 ( 
.A(n_984),
.Y(n_1162)
);

INVx3_ASAP7_75t_SL g1163 ( 
.A(n_1064),
.Y(n_1163)
);

BUFx8_ASAP7_75t_L g1164 ( 
.A(n_1030),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1038),
.B(n_1068),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_1056),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1044),
.B(n_1047),
.Y(n_1167)
);

INVx8_ASAP7_75t_L g1168 ( 
.A(n_1074),
.Y(n_1168)
);

BUFx2_ASAP7_75t_SL g1169 ( 
.A(n_991),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1038),
.B(n_1068),
.Y(n_1170)
);

BUFx4f_ASAP7_75t_SL g1171 ( 
.A(n_1064),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_1064),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1038),
.B(n_1068),
.Y(n_1173)
);

NAND2x1p5_ASAP7_75t_L g1174 ( 
.A(n_1056),
.B(n_868),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1074),
.B(n_1044),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1044),
.B(n_1047),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_1064),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1038),
.B(n_1068),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1044),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_SL g1180 ( 
.A1(n_1049),
.A2(n_1069),
.B(n_1058),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1074),
.B(n_1044),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1079),
.A2(n_1007),
.A3(n_1010),
.B(n_916),
.Y(n_1182)
);

AO21x2_ASAP7_75t_L g1183 ( 
.A1(n_1052),
.A2(n_1066),
.B(n_1061),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1044),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1044),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1109),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1175),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_1100),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1100),
.B(n_1103),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1104),
.Y(n_1190)
);

BUFx4f_ASAP7_75t_L g1191 ( 
.A(n_1168),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1103),
.B(n_1167),
.Y(n_1192)
);

OAI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1108),
.A2(n_1168),
.B1(n_1145),
.B2(n_1185),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1148),
.Y(n_1194)
);

AO21x1_ASAP7_75t_L g1195 ( 
.A1(n_1112),
.A2(n_1133),
.B(n_1152),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1107),
.Y(n_1196)
);

BUFx2_ASAP7_75t_R g1197 ( 
.A(n_1115),
.Y(n_1197)
);

NAND2x1p5_ASAP7_75t_L g1198 ( 
.A(n_1120),
.B(n_1166),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1135),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1135),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1108),
.A2(n_1145),
.B1(n_1181),
.B2(n_1106),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1184),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1168),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1159),
.A2(n_1181),
.B1(n_1128),
.B2(n_1149),
.Y(n_1204)
);

BUFx4f_ASAP7_75t_SL g1205 ( 
.A(n_1172),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1179),
.Y(n_1206)
);

BUFx4f_ASAP7_75t_SL g1207 ( 
.A(n_1172),
.Y(n_1207)
);

OR2x6_ASAP7_75t_L g1208 ( 
.A(n_1180),
.B(n_1129),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1117),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1138),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1176),
.B(n_1144),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1101),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1143),
.B(n_1157),
.Y(n_1213)
);

INVxp67_ASAP7_75t_L g1214 ( 
.A(n_1157),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1146),
.B(n_1139),
.Y(n_1215)
);

NAND2x1p5_ASAP7_75t_L g1216 ( 
.A(n_1120),
.B(n_1166),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1183),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1119),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_1162),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1174),
.Y(n_1220)
);

NOR2x1_ASAP7_75t_L g1221 ( 
.A(n_1169),
.B(n_1134),
.Y(n_1221)
);

AOI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1111),
.A2(n_1137),
.B(n_1140),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1155),
.B(n_1132),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1110),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1106),
.A2(n_1098),
.B1(n_1130),
.B2(n_1112),
.Y(n_1225)
);

CKINVDCx12_ASAP7_75t_R g1226 ( 
.A(n_1171),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1147),
.B(n_1156),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1121),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1127),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1136),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1098),
.A2(n_1150),
.B1(n_1146),
.B2(n_1142),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1124),
.A2(n_1159),
.B1(n_1178),
.B2(n_1170),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1139),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1121),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1125),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1114),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1193),
.A2(n_1173),
.B1(n_1178),
.B2(n_1165),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1219),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1208),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1215),
.B(n_1099),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1215),
.B(n_1099),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1190),
.B(n_1102),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1196),
.B(n_1102),
.Y(n_1243)
);

INVx2_ASAP7_75t_SL g1244 ( 
.A(n_1208),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1208),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1208),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1233),
.B(n_1192),
.Y(n_1247)
);

NOR2x1_ASAP7_75t_SL g1248 ( 
.A(n_1201),
.B(n_1151),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1232),
.B(n_1105),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1232),
.B(n_1160),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1202),
.B(n_1123),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1217),
.B(n_1158),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1228),
.B(n_1123),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1235),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1227),
.B(n_1113),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1227),
.B(n_1182),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1235),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1230),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1199),
.B(n_1182),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1210),
.B(n_1126),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1200),
.B(n_1182),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1230),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1224),
.B(n_1182),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1234),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1225),
.B(n_1173),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1212),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1256),
.A2(n_1231),
.B1(n_1204),
.B2(n_1214),
.Y(n_1267)
);

AND2x4_ASAP7_75t_SL g1268 ( 
.A(n_1244),
.B(n_1187),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1262),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1257),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1240),
.B(n_1195),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1253),
.B(n_1236),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1241),
.B(n_1209),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1239),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1239),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1251),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1257),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1237),
.A2(n_1189),
.B1(n_1188),
.B2(n_1191),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1251),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1255),
.B(n_1218),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1259),
.B(n_1186),
.Y(n_1281)
);

OR2x6_ASAP7_75t_SL g1282 ( 
.A(n_1237),
.B(n_1149),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1258),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1252),
.Y(n_1284)
);

NOR2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1250),
.B(n_1220),
.Y(n_1285)
);

INVxp67_ASAP7_75t_L g1286 ( 
.A(n_1254),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1255),
.B(n_1218),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1253),
.B(n_1223),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1254),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1261),
.B(n_1222),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1245),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1283),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1278),
.B(n_1244),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1280),
.B(n_1249),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1283),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1288),
.B(n_1242),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1287),
.B(n_1271),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1288),
.B(n_1242),
.Y(n_1298)
);

AND2x4_ASAP7_75t_SL g1299 ( 
.A(n_1289),
.B(n_1246),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1272),
.B(n_1243),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1272),
.B(n_1243),
.Y(n_1301)
);

AND2x4_ASAP7_75t_SL g1302 ( 
.A(n_1270),
.B(n_1246),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1268),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1271),
.B(n_1260),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1290),
.B(n_1260),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1277),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1269),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1276),
.B(n_1263),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1292),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1307),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1305),
.B(n_1284),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1306),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1296),
.B(n_1276),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1292),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1297),
.B(n_1290),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1297),
.B(n_1279),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1293),
.B(n_1264),
.C(n_1266),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1308),
.B(n_1279),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1305),
.B(n_1273),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1295),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1302),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1302),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1302),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1298),
.B(n_1264),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1299),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1304),
.B(n_1273),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1312),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1309),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1324),
.B(n_1300),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1315),
.B(n_1304),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1310),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1309),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1313),
.B(n_1318),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1316),
.B(n_1315),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1316),
.B(n_1294),
.Y(n_1335)
);

AOI21xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1325),
.A2(n_1163),
.B(n_1303),
.Y(n_1336)
);

AOI32xp33_ASAP7_75t_L g1337 ( 
.A1(n_1321),
.A2(n_1299),
.A3(n_1267),
.B1(n_1303),
.B2(n_1245),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1314),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1310),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1314),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1317),
.A2(n_1282),
.B1(n_1278),
.B2(n_1246),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1319),
.B(n_1294),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1320),
.Y(n_1343)
);

AOI32xp33_ASAP7_75t_L g1344 ( 
.A1(n_1321),
.A2(n_1299),
.A3(n_1275),
.B1(n_1291),
.B2(n_1274),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1331),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1341),
.A2(n_1317),
.B(n_1325),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1333),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1341),
.A2(n_1311),
.B1(n_1323),
.B2(n_1322),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1336),
.A2(n_1322),
.B(n_1323),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1328),
.Y(n_1350)
);

OAI21xp33_ASAP7_75t_L g1351 ( 
.A1(n_1337),
.A2(n_1318),
.B(n_1313),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1330),
.B(n_1319),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1330),
.B(n_1326),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1327),
.A2(n_1194),
.B(n_1163),
.C(n_1141),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_SL g1355 ( 
.A(n_1346),
.B(n_1344),
.C(n_1177),
.Y(n_1355)
);

NAND2x1_ASAP7_75t_L g1356 ( 
.A(n_1349),
.B(n_1342),
.Y(n_1356)
);

AOI221xp5_ASAP7_75t_L g1357 ( 
.A1(n_1351),
.A2(n_1348),
.B1(n_1354),
.B2(n_1347),
.C(n_1350),
.Y(n_1357)
);

OAI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1345),
.A2(n_1282),
.B1(n_1329),
.B2(n_1334),
.Y(n_1358)
);

NAND3xp33_ASAP7_75t_L g1359 ( 
.A(n_1345),
.B(n_1338),
.C(n_1332),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1352),
.A2(n_1248),
.B(n_1340),
.Y(n_1360)
);

AOI211xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1352),
.A2(n_1171),
.B(n_1207),
.C(n_1205),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1353),
.B(n_1205),
.Y(n_1362)
);

AND4x1_ASAP7_75t_L g1363 ( 
.A(n_1353),
.B(n_1226),
.C(n_1197),
.D(n_1115),
.Y(n_1363)
);

OAI322xp33_ASAP7_75t_L g1364 ( 
.A1(n_1348),
.A2(n_1335),
.A3(n_1343),
.B1(n_1286),
.B2(n_1301),
.C1(n_1339),
.C2(n_1331),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1347),
.Y(n_1365)
);

OAI31xp33_ASAP7_75t_L g1366 ( 
.A1(n_1346),
.A2(n_1342),
.A3(n_1285),
.B(n_1311),
.Y(n_1366)
);

NAND3xp33_ASAP7_75t_L g1367 ( 
.A(n_1357),
.B(n_1164),
.C(n_1156),
.Y(n_1367)
);

NOR3xp33_ASAP7_75t_L g1368 ( 
.A(n_1355),
.B(n_1226),
.C(n_1221),
.Y(n_1368)
);

AOI321xp33_ASAP7_75t_L g1369 ( 
.A1(n_1358),
.A2(n_1265),
.A3(n_1311),
.B1(n_1213),
.B2(n_1247),
.C(n_1281),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1365),
.B(n_1326),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1356),
.A2(n_1177),
.B(n_1191),
.Y(n_1371)
);

NOR3xp33_ASAP7_75t_L g1372 ( 
.A(n_1364),
.B(n_1118),
.C(n_1122),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1359),
.Y(n_1373)
);

NAND4xp25_ASAP7_75t_L g1374 ( 
.A(n_1361),
.B(n_1161),
.C(n_1265),
.D(n_1211),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1373),
.B(n_1362),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1367),
.B(n_1363),
.Y(n_1376)
);

NOR2x1_ASAP7_75t_L g1377 ( 
.A(n_1371),
.B(n_1148),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1372),
.B(n_1366),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1370),
.B(n_1360),
.Y(n_1379)
);

NAND3xp33_ASAP7_75t_SL g1380 ( 
.A(n_1368),
.B(n_1216),
.C(n_1198),
.Y(n_1380)
);

NAND3xp33_ASAP7_75t_L g1381 ( 
.A(n_1369),
.B(n_1164),
.C(n_1339),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1374),
.Y(n_1382)
);

NAND4xp75_ASAP7_75t_L g1383 ( 
.A(n_1378),
.B(n_1207),
.C(n_1116),
.D(n_1161),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1382),
.B(n_1311),
.Y(n_1384)
);

NOR2x1_ASAP7_75t_L g1385 ( 
.A(n_1376),
.B(n_1220),
.Y(n_1385)
);

NAND3xp33_ASAP7_75t_L g1386 ( 
.A(n_1375),
.B(n_1162),
.C(n_1153),
.Y(n_1386)
);

NAND4xp75_ASAP7_75t_L g1387 ( 
.A(n_1377),
.B(n_1116),
.C(n_1203),
.D(n_1150),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1381),
.B(n_1320),
.Y(n_1388)
);

AO22x1_ASAP7_75t_L g1389 ( 
.A1(n_1379),
.A2(n_1203),
.B1(n_1229),
.B2(n_1238),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1385),
.B(n_1386),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1388),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1384),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1387),
.A2(n_1380),
.B1(n_1285),
.B2(n_1206),
.Y(n_1393)
);

XNOR2xp5_ASAP7_75t_L g1394 ( 
.A(n_1392),
.B(n_1383),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1390),
.B(n_1389),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1394),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1396),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1397),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1398),
.A2(n_1395),
.B(n_1391),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1399),
.A2(n_1395),
.B(n_1393),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1400),
.A2(n_1154),
.B(n_1131),
.Y(n_1401)
);

OR2x6_ASAP7_75t_L g1402 ( 
.A(n_1401),
.B(n_1198),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1402),
.A2(n_1174),
.B(n_1216),
.C(n_1127),
.Y(n_1403)
);


endmodule