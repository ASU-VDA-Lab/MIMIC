module real_jpeg_6426_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_0),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_0),
.A2(n_36),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_2),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_2),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_2),
.A2(n_110),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_2),
.A2(n_110),
.B1(n_305),
.B2(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_2),
.A2(n_110),
.B1(n_362),
.B2(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_3),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_3),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_124),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_124),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_3),
.A2(n_124),
.B1(n_369),
.B2(n_394),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_4),
.B(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_4),
.B(n_271),
.C(n_273),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_4),
.A2(n_276),
.B1(n_277),
.B2(n_279),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_4),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_4),
.B(n_144),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_4),
.A2(n_24),
.B1(n_43),
.B2(n_322),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_4),
.B(n_203),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_4),
.A2(n_233),
.B(n_410),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_5),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_5),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_5),
.A2(n_253),
.B1(n_279),
.B2(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_5),
.A2(n_253),
.B1(n_311),
.B2(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_5),
.A2(n_215),
.B1(n_253),
.B2(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_7),
.A2(n_56),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_7),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_7),
.A2(n_82),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_7),
.A2(n_82),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_8),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_8),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_8),
.A2(n_115),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_8),
.A2(n_115),
.B1(n_299),
.B2(n_302),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_8),
.A2(n_115),
.B1(n_279),
.B2(n_365),
.Y(n_364)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_10),
.Y(n_157)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_10),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_10),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g383 ( 
.A(n_10),
.Y(n_383)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_13),
.Y(n_109)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_13),
.Y(n_112)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_13),
.Y(n_116)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_13),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_14),
.A2(n_48),
.B1(n_75),
.B2(n_78),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_48),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_260),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_258),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_207),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_19),
.B(n_207),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_152),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_87),
.C(n_118),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_22),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_23),
.B(n_52),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_32),
.B(n_41),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_24),
.A2(n_156),
.B(n_158),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_24),
.B(n_46),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_24),
.A2(n_32),
.B1(n_237),
.B2(n_245),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_24),
.A2(n_179),
.B(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_24),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_24),
.A2(n_43),
.B1(n_310),
.B2(n_322),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_24),
.A2(n_41),
.B(n_158),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_27),
.Y(n_244)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_27),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_27),
.Y(n_311)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_31),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_31),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_33),
.Y(n_273)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_37),
.Y(n_159)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_40),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_73),
.B1(n_81),
.B2(n_85),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_53),
.A2(n_166),
.B(n_172),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_53),
.A2(n_390),
.B(n_391),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_53),
.A2(n_172),
.B(n_393),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_54),
.A2(n_86),
.B1(n_167),
.B2(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_54),
.A2(n_86),
.B1(n_275),
.B2(n_282),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_54),
.A2(n_86),
.B1(n_282),
.B2(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_54),
.A2(n_86),
.B1(n_292),
.B2(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_67),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_58),
.B1(n_61),
.B2(n_65),
.Y(n_55)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_56),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_57),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_57),
.Y(n_278)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_57),
.Y(n_356)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_64),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_65),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_66),
.Y(n_281)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_66),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_66),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_66),
.Y(n_369)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_70),
.Y(n_241)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_74),
.B(n_86),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_80),
.B1(n_130),
.B2(n_133),
.Y(n_129)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_77),
.Y(n_168)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_85),
.B(n_276),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_85),
.B(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_87),
.A2(n_88),
.B1(n_118),
.B2(n_119),
.Y(n_209)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_107),
.B1(n_113),
.B2(n_117),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_89),
.A2(n_113),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_89),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_89),
.A2(n_117),
.B1(n_409),
.B2(n_411),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_99),
.Y(n_362)
);

INVx6_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_106),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_107),
.Y(n_257)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_108),
.A2(n_224),
.A3(n_226),
.B1(n_228),
.B2(n_232),
.Y(n_223)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_114),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_117),
.Y(n_203)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_127),
.B(n_143),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_120),
.B(n_129),
.Y(n_221)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_123),
.Y(n_229)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_123),
.Y(n_379)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_125),
.Y(n_216)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_127),
.A2(n_129),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_127),
.A2(n_129),
.B1(n_378),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_128),
.B(n_145),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_128),
.A2(n_214),
.B(n_221),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_128),
.A2(n_144),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_129),
.A2(n_188),
.B(n_194),
.Y(n_187)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_131),
.Y(n_353)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_134)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_138),
.Y(n_349)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_148),
.B(n_276),
.Y(n_350)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_174),
.B1(n_205),
.B2(n_206),
.Y(n_152)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_165),
.B2(n_173),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_163),
.Y(n_324)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_164),
.Y(n_301)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_164),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_186),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_183),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_176),
.A2(n_183),
.B1(n_184),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_178),
.A2(n_238),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_195),
.B1(n_196),
.B2(n_204),
.Y(n_186)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_189),
.A2(n_344),
.A3(n_347),
.B1(n_350),
.B2(n_351),
.Y(n_343)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_SL g360 ( 
.A1(n_190),
.A2(n_276),
.B(n_350),
.Y(n_360)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_203),
.A2(n_250),
.B1(n_256),
.B2(n_257),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_212),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_208),
.B(n_210),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_212),
.B(n_421),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_222),
.C(n_249),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_213),
.B(n_249),
.Y(n_417)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_214),
.Y(n_406)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_222),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_236),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_223),
.B(n_236),
.Y(n_402)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_250),
.Y(n_411)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_251),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_413),
.B(n_426),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_398),
.B(n_412),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_371),
.B(n_397),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_339),
.B(n_370),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_306),
.B(n_338),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_287),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_267),
.B(n_287),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_274),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_268),
.B(n_274),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_276),
.B(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_297),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_296),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_289),
.B(n_296),
.C(n_297),
.Y(n_340)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_291),
.Y(n_296)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_318),
.B(n_337),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_317),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_325),
.B(n_336),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_320),
.B(n_321),
.Y(n_336)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_SL g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_341),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_358),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_359),
.C(n_363),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_357),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_357),
.Y(n_388)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx11_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_363),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_361),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_372),
.B(n_373),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_374),
.A2(n_375),
.B1(n_386),
.B2(n_387),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_389),
.C(n_395),
.Y(n_399)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_380),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_381),
.C(n_385),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_384),
.B2(n_385),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_384),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_395),
.B2(n_396),
.Y(n_387)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_388),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_389),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_400),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_403),
.C(n_404),
.Y(n_423)
);

BUFx24_ASAP7_75t_SL g430 ( 
.A(n_404),
.Y(n_430)
);

FAx1_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_407),
.CI(n_408),
.CON(n_404),
.SN(n_404)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_407),
.C(n_408),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_422),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_414),
.A2(n_427),
.B(n_428),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_420),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_420),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.C(n_419),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_416),
.B(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_419),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_423),
.B(n_424),
.Y(n_427)
);


endmodule