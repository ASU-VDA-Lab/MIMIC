module fake_jpeg_24843_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_32),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_1),
.Y(n_32)
);

NOR3xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_2),
.C(n_4),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_25),
.B1(n_21),
.B2(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_36),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_5),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_25),
.B1(n_13),
.B2(n_16),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_16),
.B1(n_13),
.B2(n_21),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_47),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_13),
.C(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_25),
.B1(n_16),
.B2(n_13),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_67),
.B(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_64),
.Y(n_70)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_24),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_46),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_50),
.B1(n_27),
.B2(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_19),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_42),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_29),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_39),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_59),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_29),
.B(n_49),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_81),
.B(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_65),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_35),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_78),
.C(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_77),
.Y(n_86)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_18),
.A3(n_20),
.B1(n_14),
.B2(n_19),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_50),
.C(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_82),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_14),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_57),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_84),
.Y(n_102)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_92),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_58),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_71),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_55),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_96),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_68),
.Y(n_97)
);

AOI221xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_67),
.B1(n_84),
.B2(n_15),
.C(n_26),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_101),
.C(n_95),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_69),
.B(n_58),
.C(n_71),
.D(n_57),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_78),
.B1(n_62),
.B2(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_83),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_87),
.A3(n_89),
.B1(n_92),
.B2(n_96),
.C1(n_95),
.C2(n_73),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_110),
.B1(n_67),
.B2(n_51),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_112),
.B(n_115),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_81),
.C(n_60),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_113),
.Y(n_117)
);

XNOR2x1_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_85),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_60),
.C(n_80),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_107),
.C(n_103),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_116),
.B(n_27),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_106),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_102),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_35),
.A3(n_46),
.B1(n_31),
.B2(n_11),
.C1(n_12),
.C2(n_10),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_102),
.B1(n_104),
.B2(n_99),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_15),
.B1(n_20),
.B2(n_14),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_122),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_67),
.Y(n_124)
);

OAI21x1_ASAP7_75t_SL g130 ( 
.A1(n_124),
.A2(n_35),
.B(n_6),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_127),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_51),
.C(n_31),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_121),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_130),
.A3(n_123),
.B1(n_127),
.B2(n_7),
.C1(n_8),
.C2(n_5),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_9),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_35),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_6),
.B(n_8),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);


endmodule