module fake_jpeg_26367_n_80 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_80);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_7),
.B(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_33),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_3),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_52),
.B(n_37),
.C(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_3),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_54),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_35),
.B1(n_43),
.B2(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_5),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_61),
.B(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_57),
.B1(n_9),
.B2(n_11),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_67),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_68),
.C(n_71),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_57),
.C(n_13),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_6),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_17),
.Y(n_77)
);

OAI321xp33_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_18),
.A3(n_19),
.B1(n_21),
.B2(n_23),
.C(n_24),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_25),
.B(n_26),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_28),
.B(n_29),
.Y(n_80)
);


endmodule