module fake_jpeg_29111_n_531 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_531);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_531;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_52),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_53),
.Y(n_150)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_76),
.Y(n_110)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_7),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_50),
.Y(n_107)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_38),
.Y(n_72)
);

INVx5_ASAP7_75t_SL g116 ( 
.A(n_72),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_38),
.Y(n_73)
);

INVx5_ASAP7_75t_SL g131 ( 
.A(n_73),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_17),
.B(n_7),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_17),
.B(n_7),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_99),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_16),
.B(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_37),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_104),
.B(n_107),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_44),
.B1(n_19),
.B2(n_20),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_106),
.A2(n_108),
.B1(n_144),
.B2(n_152),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_44),
.B1(n_19),
.B2(n_20),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_68),
.B(n_50),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_119),
.B(n_125),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_19),
.B1(n_44),
.B2(n_32),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_122),
.A2(n_30),
.B1(n_48),
.B2(n_97),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_124),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_16),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_55),
.A2(n_25),
.B1(n_30),
.B2(n_48),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_130),
.A2(n_25),
.B1(n_35),
.B2(n_42),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_32),
.C(n_47),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_37),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_100),
.A2(n_27),
.B1(n_16),
.B2(n_45),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_20),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_60),
.A2(n_27),
.B1(n_45),
.B2(n_47),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_74),
.B(n_27),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_74),
.B(n_45),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_30),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_177),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_116),
.A2(n_52),
.B1(n_57),
.B2(n_88),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_162),
.Y(n_217)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_166),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_SL g168 ( 
.A1(n_109),
.A2(n_37),
.B(n_89),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_168),
.B(n_169),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_132),
.A2(n_35),
.B1(n_21),
.B2(n_47),
.Y(n_169)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_174),
.A2(n_180),
.B1(n_196),
.B2(n_198),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_48),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_122),
.A2(n_92),
.B1(n_91),
.B2(n_86),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_130),
.A2(n_85),
.B1(n_61),
.B2(n_62),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_181),
.A2(n_189),
.B1(n_102),
.B2(n_156),
.Y(n_247)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_110),
.B(n_21),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_200),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_209),
.B1(n_28),
.B2(n_127),
.Y(n_219)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_103),
.Y(n_186)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_190),
.Y(n_230)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_117),
.A2(n_82),
.B1(n_78),
.B2(n_135),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_144),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_205),
.Y(n_236)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_197),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_108),
.A2(n_42),
.B1(n_41),
.B2(n_26),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_117),
.A2(n_42),
.B1(n_41),
.B2(n_26),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_116),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_128),
.B(n_41),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_114),
.A2(n_32),
.B1(n_35),
.B2(n_26),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_115),
.B(n_139),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_103),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_204),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_129),
.B(n_28),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_23),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_160),
.A2(n_28),
.B1(n_25),
.B2(n_12),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_114),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_210),
.B(n_155),
.Y(n_223)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_150),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_215),
.B(n_221),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_219),
.A2(n_225),
.B1(n_234),
.B2(n_239),
.Y(n_256)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_155),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_223),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_127),
.B1(n_115),
.B2(n_135),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_226),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_207),
.B(n_156),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_228),
.B(n_249),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_194),
.A2(n_161),
.B1(n_177),
.B2(n_167),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_180),
.A2(n_118),
.B1(n_147),
.B2(n_101),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_209),
.B1(n_210),
.B2(n_169),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_243),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_191),
.A2(n_147),
.B1(n_118),
.B2(n_101),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_208),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_247),
.A2(n_204),
.B1(n_203),
.B2(n_111),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_207),
.B(n_37),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_253),
.A2(n_268),
.B1(n_269),
.B2(n_274),
.Y(n_292)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_191),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_248),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_257),
.B(n_276),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_206),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_263),
.Y(n_301)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_213),
.Y(n_261)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_183),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_176),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_273),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_176),
.C(n_164),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_224),
.C(n_242),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_221),
.A2(n_164),
.B1(n_192),
.B2(n_188),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_266),
.A2(n_237),
.B1(n_217),
.B2(n_236),
.Y(n_294)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_220),
.A2(n_170),
.B1(n_193),
.B2(n_186),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_220),
.A2(n_178),
.B1(n_171),
.B2(n_179),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_197),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_282),
.Y(n_290)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_272),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_165),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_218),
.A2(n_163),
.B1(n_173),
.B2(n_182),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_238),
.B(n_172),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_230),
.A2(n_102),
.B1(n_205),
.B2(n_105),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_278),
.B1(n_217),
.B2(n_221),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g278 ( 
.A1(n_215),
.A2(n_136),
.B1(n_195),
.B2(n_159),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_214),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_280),
.B(n_281),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_228),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_215),
.B(n_23),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_224),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_284),
.A2(n_240),
.B1(n_216),
.B2(n_229),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_245),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_285),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_316),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_281),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_288),
.B(n_263),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_294),
.A2(n_304),
.B1(n_311),
.B2(n_231),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_295),
.A2(n_261),
.B1(n_254),
.B2(n_251),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_268),
.A2(n_269),
.B1(n_253),
.B2(n_252),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_296),
.A2(n_313),
.B1(n_285),
.B2(n_276),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_259),
.A2(n_226),
.B(n_227),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_299),
.A2(n_306),
.B(n_262),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_227),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_317),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_256),
.A2(n_227),
.B1(n_236),
.B2(n_219),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_252),
.A2(n_236),
.B(n_239),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_310),
.C(n_312),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_255),
.B(n_242),
.C(n_214),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_256),
.A2(n_240),
.B1(n_246),
.B2(n_139),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_255),
.B(n_222),
.C(n_229),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_270),
.A2(n_245),
.B1(n_240),
.B2(n_246),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g314 ( 
.A(n_282),
.B(n_216),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_314),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_262),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_258),
.B(n_245),
.Y(n_317)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_319),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_280),
.Y(n_320)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

AO22x1_ASAP7_75t_L g321 ( 
.A1(n_306),
.A2(n_259),
.B1(n_266),
.B2(n_271),
.Y(n_321)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_321),
.A2(n_354),
.B(n_336),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_271),
.Y(n_322)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_257),
.Y(n_324)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_325),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_286),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_327),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_258),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_329),
.B(n_335),
.C(n_347),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_264),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_331),
.B(n_338),
.Y(n_380)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_265),
.C(n_260),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_343),
.Y(n_360)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_303),
.Y(n_334)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_334),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_290),
.B(n_273),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_336),
.A2(n_349),
.B1(n_294),
.B2(n_314),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_318),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_339),
.A2(n_231),
.B(n_241),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_340),
.A2(n_296),
.B1(n_292),
.B2(n_313),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_274),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_341),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_315),
.B(n_279),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_342),
.B(n_348),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_302),
.B(n_277),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_212),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_346),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_289),
.B(n_275),
.C(n_272),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_298),
.B(n_267),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_298),
.B(n_250),
.Y(n_350)
);

NAND3xp33_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_305),
.C(n_300),
.Y(n_369)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_353),
.A2(n_311),
.B1(n_309),
.B2(n_300),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_212),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_355),
.B(n_310),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_356),
.A2(n_343),
.B1(n_345),
.B2(n_344),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_328),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_358),
.B(n_362),
.Y(n_398)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_328),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_353),
.A2(n_292),
.B1(n_295),
.B2(n_299),
.Y(n_366)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_366),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_321),
.A2(n_314),
.B1(n_308),
.B2(n_305),
.Y(n_367)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_379),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_329),
.B(n_309),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_377),
.B(n_326),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_337),
.B(n_312),
.Y(n_379)
);

XNOR2x1_ASAP7_75t_L g382 ( 
.A(n_337),
.B(n_289),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_23),
.Y(n_417)
);

INVxp33_ASAP7_75t_L g383 ( 
.A(n_321),
.Y(n_383)
);

INVx13_ASAP7_75t_L g409 ( 
.A(n_383),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_384),
.A2(n_387),
.B1(n_388),
.B2(n_334),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_385),
.A2(n_386),
.B(n_339),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_347),
.A2(n_222),
.B1(n_241),
.B2(n_184),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_330),
.A2(n_113),
.B1(n_138),
.B2(n_121),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_351),
.Y(n_389)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_389),
.Y(n_394)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_357),
.Y(n_390)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_390),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_335),
.C(n_333),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_392),
.C(n_403),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_355),
.C(n_326),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_395),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_397),
.B(n_401),
.Y(n_423)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_368),
.Y(n_399)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_399),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_400),
.A2(n_356),
.B1(n_385),
.B2(n_373),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_380),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_402),
.A2(n_407),
.B1(n_414),
.B2(n_419),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_332),
.C(n_325),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_404),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_376),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_405),
.A2(n_412),
.B1(n_374),
.B2(n_364),
.Y(n_431)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_385),
.A2(n_352),
.B(n_323),
.Y(n_406)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_406),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_384),
.A2(n_323),
.B1(n_113),
.B2(n_134),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_166),
.C(n_212),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_396),
.C(n_392),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_175),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_375),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_387),
.A2(n_137),
.B1(n_1),
.B2(n_2),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_370),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_415),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_372),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_381),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_418),
.A2(n_11),
.B(n_15),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_359),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_433),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_424),
.B(n_439),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_360),
.C(n_371),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_425),
.B(n_429),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_393),
.A2(n_374),
.B1(n_370),
.B2(n_388),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_426),
.A2(n_435),
.B1(n_414),
.B2(n_402),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_360),
.C(n_364),
.Y(n_429)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_431),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_391),
.B(n_389),
.C(n_372),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_432),
.B(n_434),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_365),
.C(n_363),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_408),
.A2(n_365),
.B1(n_363),
.B2(n_383),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_400),
.C(n_395),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_440),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_23),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_398),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_390),
.B(n_23),
.C(n_34),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_37),
.Y(n_463)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_443),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_437),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_447),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_416),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_418),
.Y(n_449)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_449),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_411),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_454),
.Y(n_471)
);

BUFx24_ASAP7_75t_SL g455 ( 
.A(n_423),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_462),
.Y(n_474)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_436),
.Y(n_457)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_457),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_444),
.A2(n_411),
.B1(n_394),
.B2(n_409),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_458),
.A2(n_459),
.B1(n_441),
.B2(n_407),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_420),
.A2(n_394),
.B1(n_409),
.B2(n_415),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_427),
.A2(n_404),
.B(n_399),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_461),
.A2(n_464),
.B(n_419),
.Y(n_477)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_428),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_463),
.B(n_433),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_427),
.A2(n_441),
.B(n_421),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_470),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_422),
.C(n_424),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_458),
.C(n_449),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_469),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_434),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_425),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_438),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_473),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_452),
.A2(n_422),
.B1(n_439),
.B2(n_442),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_446),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_479),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_477),
.Y(n_486)
);

MAJx2_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_11),
.C(n_15),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_9),
.Y(n_480)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_480),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_464),
.B(n_6),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_481),
.B(n_445),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_459),
.A2(n_6),
.B1(n_14),
.B2(n_4),
.Y(n_482)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_482),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_446),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_487),
.B(n_489),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_474),
.B(n_448),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_465),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_491),
.B(n_492),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_498),
.Y(n_507)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_478),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_495),
.B(n_0),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_475),
.A2(n_473),
.B(n_445),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_496),
.A2(n_493),
.B(n_484),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_23),
.C(n_37),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_471),
.C(n_479),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_476),
.A2(n_5),
.B1(n_14),
.B2(n_13),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_486),
.A2(n_471),
.B1(n_470),
.B2(n_481),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_505),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_504),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_483),
.A2(n_4),
.B(n_5),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_503),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_34),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_506),
.B(n_509),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_483),
.A2(n_0),
.B(n_1),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_508),
.A2(n_507),
.B1(n_490),
.B2(n_509),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_484),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_510),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_488),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_501),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_517),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_485),
.C(n_497),
.Y(n_517)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_519),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_514),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_515),
.C(n_518),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_516),
.A2(n_507),
.B(n_504),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_511),
.B(n_516),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_523),
.A2(n_524),
.B(n_521),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_525),
.B1(n_518),
.B2(n_498),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_527),
.B(n_2),
.Y(n_528)
);

AO21x1_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_3),
.B(n_39),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_3),
.B1(n_39),
.B2(n_199),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_39),
.Y(n_531)
);


endmodule