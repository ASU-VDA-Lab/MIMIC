module fake_jpeg_2125_n_692 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_692);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_692;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_540;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_SL g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_10),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_60),
.B(n_69),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_61),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_62),
.B(n_77),
.Y(n_185)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_64),
.Y(n_168)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g194 ( 
.A(n_67),
.Y(n_194)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_68),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_70),
.Y(n_171)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_72),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_76),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_35),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_78),
.Y(n_218)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_87),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_10),
.B1(n_18),
.B2(n_17),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_85),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_86),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_28),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_91),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_92),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

HAxp5_ASAP7_75t_SL g95 ( 
.A(n_28),
.B(n_0),
.CON(n_95),
.SN(n_95)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_95),
.B(n_97),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_96),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_26),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

INVx5_ASAP7_75t_SL g101 ( 
.A(n_28),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_122),
.Y(n_146)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_111),
.Y(n_222)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_33),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_121),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_10),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_125),
.Y(n_214)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_22),
.Y(n_126)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_20),
.B(n_8),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_127),
.B(n_16),
.Y(n_186)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_21),
.Y(n_128)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_33),
.Y(n_129)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_21),
.Y(n_130)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_33),
.Y(n_131)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_23),
.Y(n_132)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_132),
.Y(n_209)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_22),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_22),
.B1(n_57),
.B2(n_34),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g302 ( 
.A1(n_141),
.A2(n_161),
.B1(n_163),
.B2(n_201),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_60),
.B(n_122),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_145),
.B(n_197),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_87),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_151),
.B(n_167),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_75),
.A2(n_40),
.B1(n_57),
.B2(n_23),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_152),
.A2(n_178),
.B1(n_215),
.B2(n_201),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_82),
.A2(n_23),
.B1(n_57),
.B2(n_34),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_95),
.A2(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_96),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_76),
.A2(n_58),
.B1(n_35),
.B2(n_47),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_177),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_78),
.A2(n_40),
.B1(n_29),
.B2(n_31),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_188),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_100),
.B(n_32),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_103),
.B(n_27),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_198),
.A2(n_101),
.B1(n_1),
.B2(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_200),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_86),
.A2(n_27),
.B1(n_38),
.B2(n_47),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_202),
.Y(n_280)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_204),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_61),
.B(n_46),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_206),
.B(n_211),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_64),
.B(n_46),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_91),
.B(n_58),
.C(n_20),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_48),
.C(n_39),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_73),
.A2(n_44),
.B1(n_38),
.B2(n_32),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_113),
.B(n_25),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_217),
.B(n_14),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_118),
.B(n_25),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_0),
.Y(n_271)
);

AO22x1_ASAP7_75t_SL g225 ( 
.A1(n_93),
.A2(n_48),
.B1(n_39),
.B2(n_33),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_0),
.Y(n_241)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_119),
.Y(n_226)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_226),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_121),
.B(n_44),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_228),
.B(n_12),
.Y(n_265)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_124),
.Y(n_229)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_229),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_125),
.Y(n_231)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_231),
.Y(n_314)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_131),
.Y(n_232)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_136),
.A2(n_85),
.B1(n_129),
.B2(n_116),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_233),
.A2(n_244),
.B1(n_260),
.B2(n_274),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_153),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_236),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_239),
.A2(n_289),
.B1(n_293),
.B2(n_297),
.Y(n_373)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_157),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_240),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_241),
.B(n_255),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_196),
.A2(n_48),
.B1(n_39),
.B2(n_11),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_245),
.Y(n_329)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_164),
.Y(n_246)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_246),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_196),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_247),
.B(n_265),
.Y(n_318)
);

BUFx6f_ASAP7_75t_SL g248 ( 
.A(n_181),
.Y(n_248)
);

BUFx2_ASAP7_75t_SL g340 ( 
.A(n_248),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_164),
.Y(n_249)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_249),
.Y(n_365)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_142),
.Y(n_250)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_250),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_185),
.B(n_11),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_252),
.B(n_257),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_168),
.Y(n_253)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_253),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_135),
.Y(n_254)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_254),
.Y(n_378)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_217),
.B(n_0),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_146),
.A2(n_48),
.B(n_39),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_256),
.A2(n_276),
.B(n_161),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_148),
.B(n_150),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_166),
.Y(n_258)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_258),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_168),
.Y(n_259)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_259),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_160),
.A2(n_48),
.B1(n_39),
.B2(n_12),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_176),
.Y(n_261)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_261),
.Y(n_350)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_165),
.Y(n_263)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_263),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_136),
.B(n_12),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_266),
.B(n_267),
.Y(n_326)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_268),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_144),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_269),
.B(n_271),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_172),
.Y(n_270)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_270),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_144),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_273),
.B(n_277),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_146),
.A2(n_8),
.B1(n_18),
.B2(n_3),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_189),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_275),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_163),
.A2(n_8),
.B(n_17),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_231),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_278),
.Y(n_369)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_190),
.Y(n_279)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_281),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_197),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_282),
.B(n_285),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_220),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_283),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_284),
.A2(n_155),
.B1(n_137),
.B2(n_139),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_222),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_209),
.Y(n_286)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_193),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_287),
.B(n_292),
.Y(n_337)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_142),
.Y(n_288)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_290),
.Y(n_346)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_199),
.Y(n_291)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_291),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_186),
.B(n_7),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_192),
.A2(n_14),
.B1(n_17),
.B2(n_4),
.Y(n_293)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_199),
.Y(n_296)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_296),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_215),
.A2(n_6),
.B1(n_16),
.B2(n_4),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_298),
.Y(n_380)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_143),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_301),
.Y(n_349)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_158),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_145),
.B(n_5),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_304),
.Y(n_351)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_213),
.Y(n_304)
);

AO22x1_ASAP7_75t_L g305 ( 
.A1(n_223),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_311),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_227),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_306),
.B(n_307),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_177),
.B(n_19),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_159),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_308),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_140),
.B(n_14),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_309),
.Y(n_343)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_227),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_310),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_172),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_312),
.Y(n_361)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_230),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_313),
.Y(n_379)
);

INVx13_ASAP7_75t_L g315 ( 
.A(n_187),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_316),
.Y(n_334)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_134),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_203),
.B(n_15),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_195),
.C(n_138),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_237),
.B(n_180),
.C(n_169),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_325),
.B(n_332),
.C(n_368),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_327),
.A2(n_244),
.B1(n_239),
.B2(n_308),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_237),
.B(n_170),
.C(n_154),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_241),
.A2(n_152),
.B1(n_178),
.B2(n_171),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_341),
.A2(n_377),
.B1(n_305),
.B2(n_310),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_342),
.A2(n_263),
.B(n_261),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_264),
.B(n_225),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_352),
.B(n_366),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_274),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_248),
.A2(n_194),
.B1(n_182),
.B2(n_218),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_359),
.A2(n_367),
.B1(n_283),
.B2(n_278),
.Y(n_407)
);

OAI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_256),
.A2(n_141),
.B1(n_174),
.B2(n_147),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_363),
.A2(n_302),
.B1(n_286),
.B2(n_250),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_251),
.B(n_214),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_276),
.A2(n_194),
.B1(n_218),
.B2(n_175),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_267),
.B(n_156),
.C(n_221),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_255),
.B(n_224),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_317),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_242),
.B(n_138),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_374),
.C(n_272),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_233),
.B(n_311),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_241),
.A2(n_171),
.B1(n_179),
.B2(n_205),
.Y(n_377)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_336),
.Y(n_382)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_382),
.Y(n_439)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_323),
.Y(n_383)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_383),
.Y(n_440)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_385),
.A2(n_399),
.B1(n_407),
.B2(n_412),
.Y(n_431)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_387),
.Y(n_448)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_388),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_389),
.B(n_391),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_390),
.A2(n_411),
.B1(n_426),
.B2(n_361),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_333),
.B(n_238),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_393),
.B(n_395),
.Y(n_437)
);

OAI32xp33_ASAP7_75t_L g394 ( 
.A1(n_352),
.A2(n_302),
.A3(n_280),
.B1(n_262),
.B2(n_299),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_394),
.B(n_398),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_321),
.B(n_234),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_396),
.A2(n_419),
.B(n_423),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_365),
.Y(n_397)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_397),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_302),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_376),
.A2(n_314),
.B1(n_295),
.B2(n_294),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_378),
.Y(n_400)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_374),
.A2(n_235),
.B1(n_243),
.B2(n_298),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_401),
.A2(n_420),
.B1(n_421),
.B2(n_424),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_343),
.B(n_258),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_402),
.B(n_410),
.Y(n_463)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_346),
.Y(n_403)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_403),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_326),
.B(n_235),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_404),
.B(n_405),
.Y(n_462)
);

AO22x2_ASAP7_75t_L g405 ( 
.A1(n_341),
.A2(n_296),
.B1(n_291),
.B2(n_288),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_349),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_406),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_342),
.A2(n_260),
.B(n_293),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_408),
.A2(n_379),
.B(n_347),
.Y(n_438)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_380),
.Y(n_409)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_409),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_330),
.B(n_290),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_355),
.A2(n_175),
.B1(n_205),
.B2(n_230),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_373),
.A2(n_240),
.B1(n_268),
.B2(n_275),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_330),
.B(n_281),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_413),
.B(n_416),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_348),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_414),
.Y(n_453)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_380),
.Y(n_415)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

AND2x2_ASAP7_75t_SL g417 ( 
.A(n_358),
.B(n_236),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_417),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_378),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_418),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_377),
.A2(n_304),
.B1(n_312),
.B2(n_270),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_358),
.A2(n_253),
.B1(n_259),
.B2(n_249),
.Y(n_421)
);

BUFx24_ASAP7_75t_L g422 ( 
.A(n_340),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_422),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_334),
.Y(n_423)
);

AO21x2_ASAP7_75t_L g424 ( 
.A1(n_334),
.A2(n_313),
.B(n_246),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_358),
.A2(n_245),
.B1(n_279),
.B2(n_149),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_425),
.A2(n_430),
.B1(n_362),
.B2(n_322),
.Y(n_468)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_344),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_427),
.A2(n_428),
.B(n_429),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_318),
.B(n_254),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_375),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_371),
.A2(n_210),
.B1(n_315),
.B2(n_15),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_432),
.A2(n_435),
.B1(n_436),
.B2(n_446),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_398),
.A2(n_343),
.B1(n_337),
.B2(n_370),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_386),
.A2(n_360),
.B1(n_368),
.B2(n_356),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_438),
.A2(n_469),
.B(n_405),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_386),
.A2(n_351),
.B1(n_379),
.B2(n_361),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_392),
.B(n_416),
.C(n_404),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_417),
.C(n_393),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_390),
.A2(n_347),
.B1(n_375),
.B2(n_320),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_450),
.A2(n_458),
.B1(n_468),
.B2(n_470),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_385),
.A2(n_332),
.B1(n_325),
.B2(n_320),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_451),
.A2(n_459),
.B1(n_460),
.B2(n_424),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_396),
.A2(n_328),
.B1(n_339),
.B2(n_357),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_423),
.A2(n_357),
.B1(n_339),
.B2(n_328),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_408),
.A2(n_345),
.B1(n_372),
.B2(n_338),
.Y(n_460)
);

OAI32xp33_ASAP7_75t_L g466 ( 
.A1(n_410),
.A2(n_319),
.A3(n_362),
.B1(n_354),
.B2(n_353),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_405),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_419),
.A2(n_335),
.B(n_344),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_394),
.A2(n_338),
.B1(n_372),
.B2(n_365),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_424),
.A2(n_335),
.B1(n_319),
.B2(n_353),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_471),
.A2(n_424),
.B1(n_421),
.B2(n_420),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_406),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g538 ( 
.A(n_473),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_457),
.B(n_392),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_474),
.B(n_494),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_475),
.A2(n_479),
.B1(n_485),
.B2(n_487),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_472),
.A2(n_414),
.B1(n_411),
.B2(n_413),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_476),
.A2(n_496),
.B(n_497),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_477),
.B(n_480),
.Y(n_539)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_436),
.B(n_449),
.CI(n_435),
.CON(n_478),
.SN(n_478)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_478),
.B(n_492),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_456),
.A2(n_424),
.B1(n_401),
.B2(n_417),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_381),
.Y(n_481)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_481),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_482),
.B(n_488),
.C(n_502),
.Y(n_524)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_433),
.Y(n_484)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_484),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_462),
.A2(n_405),
.B1(n_430),
.B2(n_425),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_469),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_491),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_456),
.A2(n_405),
.B1(n_382),
.B2(n_429),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_449),
.B(n_403),
.C(n_383),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_433),
.Y(n_489)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_489),
.Y(n_522)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_439),
.Y(n_490)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_490),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_453),
.B(n_415),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_445),
.B(n_409),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_463),
.B(n_384),
.Y(n_493)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_493),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_457),
.B(n_388),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_427),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_499),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_434),
.A2(n_418),
.B(n_400),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_437),
.B(n_387),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_498),
.B(n_501),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_448),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_462),
.A2(n_397),
.B1(n_426),
.B2(n_354),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_500),
.A2(n_510),
.B1(n_441),
.B2(n_471),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_465),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_457),
.B(n_364),
.C(n_350),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_503),
.B(n_504),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_448),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_465),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_505),
.B(n_507),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_459),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_446),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_508),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_461),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_509),
.Y(n_528)
);

OA21x2_ASAP7_75t_L g510 ( 
.A1(n_438),
.A2(n_331),
.B(n_350),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_455),
.B(n_331),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_511),
.B(n_455),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_481),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_513),
.B(n_518),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_508),
.A2(n_432),
.B1(n_431),
.B2(n_438),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_514),
.B(n_546),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_474),
.B(n_451),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_516),
.B(n_517),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_482),
.B(n_488),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_491),
.Y(n_518)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_520),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_502),
.B(n_472),
.C(n_437),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_525),
.B(n_547),
.C(n_548),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_529),
.A2(n_530),
.B1(n_531),
.B2(n_537),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_487),
.A2(n_470),
.B1(n_450),
.B2(n_441),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_480),
.A2(n_477),
.B1(n_479),
.B2(n_505),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_494),
.B(n_461),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_SL g561 ( 
.A(n_533),
.B(n_543),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_492),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_535),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_507),
.A2(n_458),
.B1(n_468),
.B2(n_460),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_SL g543 ( 
.A(n_478),
.B(n_434),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_473),
.B(n_493),
.Y(n_544)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_544),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_495),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_545),
.A2(n_526),
.B1(n_538),
.B2(n_515),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_483),
.A2(n_431),
.B1(n_443),
.B2(n_464),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_478),
.B(n_447),
.C(n_440),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_483),
.B(n_466),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_536),
.Y(n_550)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_550),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_527),
.A2(n_501),
.B1(n_506),
.B2(n_486),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_555),
.A2(n_559),
.B1(n_560),
.B2(n_564),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_517),
.B(n_497),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_556),
.B(n_565),
.Y(n_586)
);

A2O1A1Ixp33_ASAP7_75t_L g558 ( 
.A1(n_541),
.A2(n_496),
.B(n_486),
.C(n_510),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_558),
.B(n_571),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_527),
.A2(n_506),
.B1(n_476),
.B2(n_485),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_531),
.A2(n_510),
.B1(n_499),
.B2(n_504),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_524),
.B(n_447),
.C(n_511),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_562),
.B(n_578),
.C(n_570),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_512),
.B(n_510),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g594 ( 
.A(n_563),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_530),
.A2(n_503),
.B1(n_489),
.B2(n_484),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_524),
.B(n_498),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_525),
.B(n_500),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_568),
.B(n_581),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_540),
.A2(n_475),
.B(n_467),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_569),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_539),
.A2(n_490),
.B1(n_442),
.B2(n_443),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_528),
.Y(n_572)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_572),
.Y(n_597)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_573),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_512),
.B(n_440),
.Y(n_574)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_574),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_548),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_575),
.B(n_576),
.Y(n_598)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_521),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_521),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_577),
.B(n_579),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_516),
.B(n_454),
.C(n_452),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_536),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_515),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_580),
.B(n_582),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_543),
.B(n_454),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_522),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_583),
.B(n_591),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_562),
.B(n_547),
.C(n_549),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_584),
.B(n_588),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_567),
.B(n_519),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_570),
.B(n_532),
.C(n_540),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_589),
.B(n_590),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_557),
.B(n_578),
.C(n_565),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_557),
.B(n_532),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_556),
.B(n_541),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_592),
.B(n_596),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_568),
.B(n_546),
.C(n_514),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_593),
.B(n_599),
.C(n_605),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_581),
.B(n_534),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_561),
.B(n_533),
.C(n_539),
.Y(n_599)
);

MAJx2_ASAP7_75t_L g600 ( 
.A(n_561),
.B(n_539),
.C(n_526),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_SL g621 ( 
.A(n_600),
.B(n_563),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_555),
.B(n_523),
.C(n_529),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_569),
.B(n_537),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_606),
.B(n_571),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_590),
.B(n_558),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_611),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_602),
.A2(n_553),
.B1(n_559),
.B2(n_554),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g639 ( 
.A1(n_613),
.A2(n_614),
.B1(n_628),
.B2(n_444),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_604),
.A2(n_554),
.B1(n_560),
.B2(n_550),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_608),
.A2(n_552),
.B1(n_566),
.B2(n_551),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_615),
.A2(n_618),
.B1(n_364),
.B2(n_329),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_585),
.Y(n_616)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_616),
.Y(n_636)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_607),
.Y(n_617)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_617),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_605),
.A2(n_574),
.B1(n_563),
.B2(n_522),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_597),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_619),
.B(n_630),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_620),
.B(n_621),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_603),
.A2(n_595),
.B1(n_601),
.B2(n_594),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_623),
.A2(n_329),
.B1(n_322),
.B2(n_324),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_584),
.B(n_564),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_624),
.B(n_626),
.Y(n_635)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_598),
.Y(n_625)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_625),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_583),
.B(n_444),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_600),
.Y(n_627)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_627),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_606),
.A2(n_523),
.B1(n_542),
.B2(n_467),
.Y(n_628)
);

FAx1_ASAP7_75t_SL g630 ( 
.A(n_599),
.B(n_464),
.CI(n_442),
.CON(n_630),
.SN(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_611),
.B(n_593),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_631),
.B(n_632),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_622),
.B(n_586),
.C(n_592),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_623),
.A2(n_596),
.B(n_586),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_633),
.A2(n_646),
.B(n_649),
.Y(n_660)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_639),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_622),
.B(n_587),
.C(n_591),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_640),
.B(n_643),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_616),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_609),
.B(n_587),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_645),
.B(n_609),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_614),
.A2(n_589),
.B(n_452),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_647),
.A2(n_369),
.B1(n_422),
.B2(n_15),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_SL g651 ( 
.A1(n_648),
.A2(n_643),
.B1(n_636),
.B2(n_638),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_628),
.A2(n_613),
.B(n_620),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_650),
.B(n_654),
.Y(n_671)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_651),
.Y(n_668)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_640),
.B(n_610),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_652),
.B(n_656),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_635),
.B(n_612),
.Y(n_653)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_653),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_632),
.B(n_629),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_634),
.B(n_610),
.Y(n_656)
);

AOI21x1_ASAP7_75t_L g657 ( 
.A1(n_633),
.A2(n_630),
.B(n_621),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_657),
.A2(n_662),
.B(n_637),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_644),
.A2(n_630),
.B1(n_369),
.B2(n_422),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_658),
.B(n_655),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_636),
.Y(n_659)
);

INVxp33_ASAP7_75t_L g667 ( 
.A(n_659),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_661),
.B(n_638),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_SL g662 ( 
.A1(n_641),
.A2(n_422),
.B(n_634),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_SL g666 ( 
.A(n_660),
.B(n_646),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_666),
.Y(n_682)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_654),
.B(n_641),
.C(n_645),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_669),
.B(n_670),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g670 ( 
.A(n_664),
.B(n_649),
.C(n_639),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_673),
.B(n_659),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_674),
.B(n_675),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_672),
.B(n_653),
.C(n_663),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_676),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_665),
.A2(n_650),
.B(n_637),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_SL g685 ( 
.A1(n_678),
.A2(n_667),
.B(n_671),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_679),
.A2(n_681),
.B(n_671),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_667),
.B(n_635),
.Y(n_681)
);

XNOR2xp5_ASAP7_75t_L g687 ( 
.A(n_684),
.B(n_685),
.Y(n_687)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g686 ( 
.A1(n_682),
.A2(n_680),
.B(n_666),
.C(n_668),
.D(n_642),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_SL g688 ( 
.A1(n_686),
.A2(n_680),
.B(n_677),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_688),
.B(n_683),
.Y(n_689)
);

BUFx24_ASAP7_75t_SL g690 ( 
.A(n_689),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_690),
.A2(n_687),
.B(n_642),
.Y(n_691)
);

XNOR2xp5_ASAP7_75t_L g692 ( 
.A(n_691),
.B(n_648),
.Y(n_692)
);


endmodule