module fake_netlist_6_3444_n_774 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_774);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_774;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_608;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_65),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_1),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_71),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_70),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_106),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_102),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_116),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_42),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_60),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_99),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_19),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_74),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_83),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_39),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_127),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_113),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_11),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_51),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_57),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_134),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_50),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_91),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_45),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_33),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_89),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_58),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_48),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_22),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_76),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_8),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_40),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_59),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_135),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_3),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_120),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_1),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_84),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_87),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_17),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_27),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_140),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_154),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_157),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_L g217 ( 
.A(n_159),
.B(n_0),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_160),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_0),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_154),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_155),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_156),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_161),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_R g228 ( 
.A(n_164),
.B(n_21),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_162),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_2),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_163),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_159),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_165),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_179),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_167),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_215),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_185),
.B1(n_197),
.B2(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_209),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_190),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_213),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_217),
.B(n_174),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_190),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_218),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_219),
.B(n_174),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_219),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_211),
.B(n_205),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

BUFx8_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

OA21x2_ASAP7_75t_L g281 ( 
.A1(n_220),
.A2(n_206),
.B(n_198),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_236),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_243),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_230),
.B(n_195),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_242),
.B(n_168),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_242),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_171),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_244),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_215),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_222),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_252),
.B(n_172),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_173),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_281),
.B(n_291),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_268),
.Y(n_305)
);

AND2x6_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_174),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_258),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_250),
.B(n_175),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_281),
.B1(n_289),
.B2(n_259),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_254),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_176),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_180),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_258),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_254),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_269),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_285),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

AO21x2_ASAP7_75t_L g323 ( 
.A1(n_257),
.A2(n_194),
.B(n_193),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

NAND3x1_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_3),
.C(n_4),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_277),
.B(n_222),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_282),
.A2(n_187),
.B1(n_184),
.B2(n_182),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_248),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_174),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_SL g331 ( 
.A(n_283),
.B(n_210),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_271),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_251),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_284),
.B(n_210),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_271),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_260),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_260),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_273),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_L g340 ( 
.A(n_279),
.B(n_4),
.C(n_5),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_251),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_284),
.B(n_286),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_249),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_264),
.B(n_5),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_253),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_270),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_266),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_275),
.B(n_23),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_280),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_267),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_270),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_255),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_263),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_255),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_296),
.B(n_288),
.Y(n_357)
);

OAI221xp5_ASAP7_75t_L g358 ( 
.A1(n_312),
.A2(n_267),
.B1(n_256),
.B2(n_257),
.C(n_281),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_350),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_355),
.Y(n_361)
);

NAND2x1p5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_263),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_343),
.A2(n_310),
.B1(n_302),
.B2(n_297),
.Y(n_363)
);

AO22x2_ASAP7_75t_L g364 ( 
.A1(n_309),
.A2(n_288),
.B1(n_293),
.B2(n_292),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_256),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_355),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_326),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_297),
.B(n_263),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_280),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_348),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_290),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_343),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_320),
.B(n_280),
.Y(n_375)
);

AO22x2_ASAP7_75t_L g376 ( 
.A1(n_340),
.A2(n_292),
.B1(n_7),
.B2(n_8),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_354),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_298),
.B(n_247),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_294),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_353),
.B(n_6),
.Y(n_383)
);

OAI221xp5_ASAP7_75t_L g384 ( 
.A1(n_299),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_384)
);

OR2x6_ASAP7_75t_L g385 ( 
.A(n_325),
.B(n_9),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_304),
.Y(n_388)
);

OAI221xp5_ASAP7_75t_L g389 ( 
.A1(n_314),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_305),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_24),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_324),
.Y(n_393)
);

AO22x1_ASAP7_75t_L g394 ( 
.A1(n_350),
.A2(n_330),
.B1(n_345),
.B2(n_306),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

OAI221xp5_ASAP7_75t_L g397 ( 
.A1(n_314),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_319),
.B(n_274),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_335),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

AO22x2_ASAP7_75t_L g401 ( 
.A1(n_335),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_329),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_344),
.B(n_25),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_302),
.A2(n_274),
.B1(n_88),
.B2(n_90),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_334),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_334),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_323),
.A2(n_85),
.B1(n_152),
.B2(n_151),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_337),
.B(n_16),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_338),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_341),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

OAI221xp5_ASAP7_75t_L g413 ( 
.A1(n_342),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.C(n_20),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

OAI221xp5_ASAP7_75t_L g416 ( 
.A1(n_352),
.A2(n_18),
.B1(n_20),
.B2(n_26),
.C(n_28),
.Y(n_416)
);

AO22x2_ASAP7_75t_L g417 ( 
.A1(n_325),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_328),
.B(n_32),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

AO22x2_ASAP7_75t_L g421 ( 
.A1(n_327),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_320),
.B(n_37),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_322),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_322),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_374),
.B(n_320),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_363),
.B(n_351),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_360),
.B(n_351),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_360),
.B(n_323),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_400),
.B(n_300),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_SL g430 ( 
.A(n_391),
.B(n_300),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g431 ( 
.A(n_391),
.B(n_300),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_SL g432 ( 
.A(n_375),
.B(n_308),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_400),
.B(n_308),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_406),
.B(n_390),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_SL g435 ( 
.A(n_371),
.B(n_308),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_406),
.B(n_333),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_419),
.B(n_333),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_419),
.B(n_333),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_365),
.B(n_303),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_392),
.B(n_336),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_365),
.B(n_303),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_392),
.B(n_303),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_399),
.B(n_303),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_SL g444 ( 
.A(n_387),
.B(n_307),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_SL g445 ( 
.A(n_372),
.B(n_307),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_379),
.B(n_307),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_373),
.B(n_307),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_SL g448 ( 
.A(n_422),
.B(n_321),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_373),
.B(n_321),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_388),
.B(n_321),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_370),
.B(n_321),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_403),
.B(n_315),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_403),
.B(n_322),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_414),
.B(n_322),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_377),
.B(n_316),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_357),
.B(n_367),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_362),
.B(n_317),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_415),
.B(n_295),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_361),
.B(n_295),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_380),
.B(n_301),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_378),
.B(n_318),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_SL g462 ( 
.A(n_383),
.B(n_409),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_366),
.B(n_301),
.Y(n_463)
);

AND3x1_ASAP7_75t_L g464 ( 
.A(n_369),
.B(n_311),
.C(n_318),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_368),
.B(n_311),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_SL g466 ( 
.A(n_420),
.B(n_318),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_359),
.B(n_306),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_410),
.B(n_382),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_386),
.B(n_393),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_395),
.B(n_306),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_396),
.B(n_306),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_SL g472 ( 
.A(n_402),
.B(n_306),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_405),
.B(n_407),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_411),
.B(n_38),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_412),
.B(n_41),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_SL g476 ( 
.A(n_418),
.B(n_43),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_404),
.B(n_44),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_364),
.B(n_46),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_408),
.B(n_47),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_398),
.B(n_49),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_385),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_445),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_461),
.A2(n_424),
.B(n_423),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_455),
.A2(n_474),
.B(n_463),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_440),
.A2(n_358),
.B1(n_417),
.B2(n_364),
.Y(n_485)
);

AO31x2_ASAP7_75t_L g486 ( 
.A1(n_428),
.A2(n_394),
.A3(n_416),
.B(n_421),
.Y(n_486)
);

OAI22x1_ASAP7_75t_L g487 ( 
.A1(n_426),
.A2(n_385),
.B1(n_417),
.B2(n_401),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_478),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_459),
.A2(n_421),
.B(n_53),
.Y(n_489)
);

A2O1A1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_452),
.A2(n_397),
.B(n_389),
.C(n_384),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_477),
.A2(n_479),
.B(n_480),
.Y(n_491)
);

NAND3x1_ASAP7_75t_L g492 ( 
.A(n_427),
.B(n_401),
.C(n_376),
.Y(n_492)
);

A2O1A1Ixp33_ASAP7_75t_L g493 ( 
.A1(n_452),
.A2(n_413),
.B(n_376),
.C(n_381),
.Y(n_493)
);

AO32x2_ASAP7_75t_L g494 ( 
.A1(n_464),
.A2(n_153),
.A3(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_453),
.A2(n_52),
.B(n_61),
.Y(n_495)
);

OA21x2_ASAP7_75t_L g496 ( 
.A1(n_451),
.A2(n_62),
.B(n_63),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_446),
.B(n_150),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_469),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_460),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_64),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_R g501 ( 
.A(n_444),
.B(n_66),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_442),
.A2(n_67),
.B(n_68),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_430),
.A2(n_69),
.B(n_72),
.Y(n_503)
);

OA22x2_ASAP7_75t_L g504 ( 
.A1(n_425),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_434),
.B(n_149),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_432),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_465),
.A2(n_78),
.B(n_80),
.Y(n_507)
);

AO21x2_ASAP7_75t_L g508 ( 
.A1(n_457),
.A2(n_81),
.B(n_82),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_473),
.A2(n_86),
.B(n_92),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_476),
.Y(n_510)
);

A2O1A1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_448),
.A2(n_93),
.B(n_94),
.C(n_95),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_448),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_431),
.A2(n_97),
.B(n_98),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_458),
.A2(n_100),
.B(n_101),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_468),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_454),
.A2(n_107),
.B(n_108),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_437),
.A2(n_438),
.B(n_433),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_447),
.B(n_109),
.Y(n_518)
);

AO31x2_ASAP7_75t_L g519 ( 
.A1(n_466),
.A2(n_110),
.A3(n_111),
.B(n_112),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_449),
.B(n_114),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_429),
.A2(n_115),
.B(n_117),
.Y(n_521)
);

INVx2_ASAP7_75t_R g522 ( 
.A(n_435),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_450),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_436),
.A2(n_118),
.B(n_119),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_470),
.A2(n_121),
.B(n_125),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_443),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_SL g527 ( 
.A(n_475),
.B(n_126),
.C(n_128),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_471),
.A2(n_147),
.B(n_131),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_439),
.B(n_146),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_488),
.B(n_441),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_498),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_523),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_483),
.A2(n_467),
.B(n_472),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_481),
.A2(n_130),
.B1(n_133),
.B2(n_136),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_491),
.A2(n_138),
.B(n_139),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_141),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_526),
.B(n_144),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_505),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_499),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_518),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_484),
.A2(n_145),
.B(n_514),
.Y(n_541)
);

OAI22xp33_ASAP7_75t_L g542 ( 
.A1(n_487),
.A2(n_482),
.B1(n_500),
.B2(n_504),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_507),
.A2(n_509),
.B(n_516),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_529),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_492),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_525),
.A2(n_489),
.B(n_517),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_493),
.B(n_490),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_506),
.B(n_520),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_485),
.B(n_510),
.Y(n_549)
);

INVx6_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_512),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g552 ( 
.A1(n_491),
.A2(n_503),
.B(n_513),
.Y(n_552)
);

OAI21x1_ASAP7_75t_SL g553 ( 
.A1(n_528),
.A2(n_497),
.B(n_502),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_486),
.B(n_522),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_486),
.B(n_527),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_508),
.Y(n_556)
);

AOI222xp33_ASAP7_75t_L g557 ( 
.A1(n_528),
.A2(n_511),
.B1(n_494),
.B2(n_515),
.C1(n_486),
.C2(n_495),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_515),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_521),
.B(n_524),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_508),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_496),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_519),
.A2(n_483),
.B(n_484),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_519),
.A2(n_483),
.B(n_484),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_519),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_494),
.Y(n_565)
);

BUFx12f_ASAP7_75t_L g566 ( 
.A(n_494),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_488),
.B(n_374),
.Y(n_567)
);

AO21x2_ASAP7_75t_L g568 ( 
.A1(n_491),
.A2(n_363),
.B(n_483),
.Y(n_568)
);

AO21x2_ASAP7_75t_L g569 ( 
.A1(n_491),
.A2(n_363),
.B(n_483),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_488),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_498),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_567),
.B(n_547),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_571),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_571),
.B(n_532),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_554),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_570),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_550),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_554),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_564),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_531),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_564),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_549),
.B(n_565),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_562),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_570),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_561),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_540),
.B(n_538),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_563),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_568),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_551),
.Y(n_589)
);

CKINVDCx6p67_ASAP7_75t_R g590 ( 
.A(n_567),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_555),
.B(n_569),
.Y(n_591)
);

OAI21x1_ASAP7_75t_SL g592 ( 
.A1(n_553),
.A2(n_535),
.B(n_560),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_569),
.B(n_568),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_568),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_548),
.B(n_550),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_569),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_544),
.B(n_558),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_552),
.A2(n_558),
.B(n_559),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_556),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_548),
.B(n_545),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_548),
.B(n_530),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_546),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_550),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_566),
.B(n_552),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_530),
.B(n_550),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_542),
.B(n_536),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_541),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_539),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_560),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_536),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_537),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_566),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_572),
.B(n_611),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_606),
.B(n_534),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_602),
.B(n_543),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_575),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_576),
.B(n_533),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_R g619 ( 
.A(n_604),
.B(n_557),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_602),
.B(n_577),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_584),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_584),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_597),
.B(n_595),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_SL g624 ( 
.A(n_597),
.B(n_577),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_586),
.B(n_607),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_584),
.Y(n_626)
);

CKINVDCx11_ASAP7_75t_R g627 ( 
.A(n_590),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_586),
.B(n_574),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_574),
.B(n_612),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_577),
.B(n_600),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_612),
.B(n_589),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_R g632 ( 
.A(n_590),
.B(n_577),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_609),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_605),
.B(n_598),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_600),
.B(n_580),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_580),
.B(n_573),
.Y(n_636)
);

NOR2x1_ASAP7_75t_L g637 ( 
.A(n_612),
.B(n_610),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_582),
.B(n_573),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_575),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_R g640 ( 
.A(n_599),
.B(n_601),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_599),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_582),
.B(n_578),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_613),
.B(n_578),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_599),
.B(n_613),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_599),
.B(n_601),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_591),
.B(n_585),
.Y(n_646)
);

INVxp67_ASAP7_75t_SL g647 ( 
.A(n_585),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_605),
.B(n_579),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_599),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_637),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_643),
.B(n_605),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_637),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_642),
.B(n_591),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_615),
.A2(n_605),
.B1(n_592),
.B2(n_579),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_617),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_639),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_646),
.B(n_605),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_638),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_644),
.Y(n_659)
);

INVxp67_ASAP7_75t_SL g660 ( 
.A(n_647),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_631),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_623),
.B(n_599),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_634),
.B(n_581),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_645),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_614),
.B(n_610),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_616),
.B(n_596),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_636),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_636),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_634),
.B(n_616),
.Y(n_669)
);

INVxp67_ASAP7_75t_SL g670 ( 
.A(n_629),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_645),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_634),
.B(n_581),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_625),
.B(n_628),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_648),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_622),
.B(n_593),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_644),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_635),
.B(n_594),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_656),
.Y(n_678)
);

AND2x2_ASAP7_75t_SL g679 ( 
.A(n_669),
.B(n_654),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_660),
.A2(n_624),
.B(n_592),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_675),
.A2(n_618),
.B(n_630),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_666),
.B(n_657),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_669),
.B(n_641),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_655),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_674),
.A2(n_619),
.B1(n_621),
.B2(n_626),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_674),
.A2(n_620),
.B1(n_630),
.B2(n_635),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_656),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_653),
.B(n_593),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_656),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_666),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_666),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_655),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_661),
.B(n_633),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_657),
.B(n_596),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_683),
.B(n_664),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_682),
.B(n_651),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_693),
.B(n_661),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_684),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_651),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_690),
.B(n_663),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_690),
.B(n_691),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_691),
.B(n_663),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_678),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_694),
.B(n_670),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_692),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_695),
.Y(n_706)
);

AO221x2_ASAP7_75t_L g707 ( 
.A1(n_697),
.A2(n_681),
.B1(n_673),
.B2(n_679),
.C(n_665),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_R g708 ( 
.A(n_695),
.B(n_632),
.Y(n_708)
);

INVxp33_ASAP7_75t_L g709 ( 
.A(n_704),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_698),
.B(n_694),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_706),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_710),
.B(n_699),
.Y(n_712)
);

AND3x1_ASAP7_75t_L g713 ( 
.A(n_707),
.B(n_685),
.C(n_705),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_SL g714 ( 
.A1(n_707),
.A2(n_680),
.B(n_660),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_713),
.A2(n_679),
.B1(n_708),
.B2(n_672),
.Y(n_715)
);

OAI21xp5_ASAP7_75t_L g716 ( 
.A1(n_714),
.A2(n_709),
.B(n_670),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_711),
.A2(n_673),
.B(n_662),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_712),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_718),
.B(n_712),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_717),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_715),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_719),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_720),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_719),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_721),
.Y(n_725)
);

NAND4xp25_ASAP7_75t_L g726 ( 
.A(n_725),
.B(n_716),
.C(n_686),
.D(n_665),
.Y(n_726)
);

NOR3xp33_ASAP7_75t_L g727 ( 
.A(n_723),
.B(n_627),
.C(n_649),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_L g728 ( 
.A(n_723),
.B(n_652),
.C(n_650),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_722),
.B(n_652),
.C(n_650),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_SL g730 ( 
.A(n_724),
.B(n_667),
.C(n_668),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_722),
.B(n_703),
.Y(n_731)
);

NAND4xp75_ASAP7_75t_L g732 ( 
.A(n_725),
.B(n_672),
.C(n_699),
.D(n_696),
.Y(n_732)
);

NAND4xp25_ASAP7_75t_L g733 ( 
.A(n_725),
.B(n_659),
.C(n_676),
.D(n_649),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_732),
.Y(n_734)
);

NOR2x1_ASAP7_75t_L g735 ( 
.A(n_731),
.B(n_728),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_729),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_730),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_726),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_727),
.B(n_733),
.Y(n_739)
);

NOR3xp33_ASAP7_75t_L g740 ( 
.A(n_727),
.B(n_641),
.C(n_658),
.Y(n_740)
);

OAI211xp5_ASAP7_75t_SL g741 ( 
.A1(n_727),
.A2(n_688),
.B(n_653),
.C(n_668),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_734),
.A2(n_695),
.B1(n_683),
.B2(n_671),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_737),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_740),
.A2(n_683),
.B1(n_671),
.B2(n_664),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_736),
.B(n_696),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_735),
.Y(n_746)
);

XNOR2xp5_ASAP7_75t_L g747 ( 
.A(n_738),
.B(n_620),
.Y(n_747)
);

NAND3x1_ASAP7_75t_L g748 ( 
.A(n_739),
.B(n_700),
.C(n_702),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_741),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_SL g750 ( 
.A(n_746),
.B(n_640),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_SL g751 ( 
.A(n_745),
.B(n_749),
.Y(n_751)
);

XOR2xp5_ASAP7_75t_L g752 ( 
.A(n_747),
.B(n_658),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_R g753 ( 
.A(n_743),
.B(n_748),
.Y(n_753)
);

NAND2x1_ASAP7_75t_SL g754 ( 
.A(n_742),
.B(n_744),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_746),
.B(n_703),
.C(n_687),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_R g756 ( 
.A(n_746),
.B(n_659),
.Y(n_756)
);

AOI222xp33_ASAP7_75t_L g757 ( 
.A1(n_751),
.A2(n_702),
.B1(n_700),
.B2(n_701),
.C1(n_659),
.C2(n_676),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_752),
.A2(n_701),
.B1(n_664),
.B2(n_671),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_756),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_753),
.Y(n_760)
);

XNOR2x1_ASAP7_75t_L g761 ( 
.A(n_755),
.B(n_676),
.Y(n_761)
);

NOR3xp33_ASAP7_75t_L g762 ( 
.A(n_750),
.B(n_667),
.C(n_688),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_760),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_759),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_L g765 ( 
.A1(n_761),
.A2(n_754),
.B(n_762),
.Y(n_765)
);

AO22x1_ASAP7_75t_L g766 ( 
.A1(n_763),
.A2(n_758),
.B1(n_757),
.B2(n_689),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_764),
.B(n_689),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_765),
.B(n_687),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_678),
.B1(n_677),
.B2(n_608),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_769),
.B(n_767),
.C(n_766),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_770),
.A2(n_608),
.B(n_603),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_771),
.Y(n_772)
);

AOI221xp5_ASAP7_75t_L g773 ( 
.A1(n_772),
.A2(n_608),
.B1(n_583),
.B2(n_587),
.C(n_594),
.Y(n_773)
);

AOI211xp5_ASAP7_75t_L g774 ( 
.A1(n_773),
.A2(n_588),
.B(n_677),
.C(n_583),
.Y(n_774)
);


endmodule