module fake_jpeg_1556_n_74 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_16),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_26),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_28),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_27),
.Y(n_45)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_22),
.C(n_10),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_25),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_39),
.B1(n_26),
.B2(n_36),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_39),
.B(n_38),
.Y(n_48)
);

OA21x2_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_4),
.B(n_5),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_50),
.B1(n_22),
.B2(n_13),
.Y(n_58)
);

AO21x2_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_36),
.B(n_25),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_3),
.C(n_4),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_60),
.Y(n_65)
);

NOR3xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_53),
.C(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_63),
.B(n_66),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_59),
.C(n_56),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_65),
.C(n_64),
.Y(n_69)
);

AOI31xp67_ASAP7_75t_SL g70 ( 
.A1(n_69),
.A2(n_68),
.A3(n_12),
.B(n_14),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_18),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_71),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_19),
.C(n_6),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_7),
.Y(n_74)
);


endmodule