module fake_jpeg_29337_n_353 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_46),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_25),
.A2(n_8),
.B(n_15),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_54),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g54 ( 
.A(n_25),
.B(n_0),
.CON(n_54),
.SN(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_60),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_64),
.B(n_73),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_22),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_76),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_28),
.B1(n_20),
.B2(n_31),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_75),
.B1(n_28),
.B2(n_31),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_29),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_77),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_28),
.B1(n_20),
.B2(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_37),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_21),
.C(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_35),
.B1(n_39),
.B2(n_37),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_80),
.A2(n_100),
.B1(n_17),
.B2(n_27),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_83),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_30),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_33),
.Y(n_112)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_19),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_52),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_55),
.B(n_19),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_55),
.B(n_22),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_40),
.B1(n_27),
.B2(n_17),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_106),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_110),
.A2(n_127),
.B1(n_134),
.B2(n_17),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_112),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_114),
.B(n_124),
.Y(n_172)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_28),
.B1(n_23),
.B2(n_24),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_128),
.B1(n_63),
.B2(n_78),
.Y(n_148)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_75),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_136),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_23),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_122),
.B(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_71),
.B(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_77),
.B(n_40),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_27),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_26),
.B1(n_23),
.B2(n_29),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_88),
.A2(n_91),
.B1(n_72),
.B2(n_85),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_63),
.A2(n_98),
.B(n_78),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

AO22x2_ASAP7_75t_L g132 ( 
.A1(n_68),
.A2(n_29),
.B1(n_24),
.B2(n_26),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_81),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

OAI21x1_ASAP7_75t_L g196 ( 
.A1(n_142),
.A2(n_174),
.B(n_175),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_24),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_165),
.C(n_136),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_148),
.A2(n_152),
.B1(n_156),
.B2(n_129),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_68),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_150),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_94),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_94),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_153),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_61),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_87),
.B1(n_61),
.B2(n_67),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_157),
.B(n_160),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_122),
.B(n_13),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_159),
.B(n_161),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_134),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_130),
.C(n_107),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_33),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_177),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_117),
.B(n_101),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_34),
.B(n_36),
.C(n_2),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_109),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_104),
.B(n_67),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_104),
.B(n_103),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_105),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_205),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_110),
.B1(n_127),
.B2(n_97),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_185),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

INVx11_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

INVx6_ASAP7_75t_SL g233 ( 
.A(n_186),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_140),
.B1(n_138),
.B2(n_97),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_190),
.B1(n_202),
.B2(n_212),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_36),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_192),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_109),
.B1(n_34),
.B2(n_123),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_14),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_133),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_145),
.A2(n_105),
.B(n_118),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

CKINVDCx10_ASAP7_75t_R g228 ( 
.A(n_206),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_33),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_208),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_175),
.A2(n_70),
.B1(n_103),
.B2(n_66),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_211),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

BUFx16f_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_145),
.A2(n_129),
.B(n_118),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_148),
.A2(n_169),
.B1(n_154),
.B2(n_174),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_156),
.A2(n_70),
.B1(n_123),
.B2(n_102),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_213),
.A2(n_164),
.B1(n_173),
.B2(n_154),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_149),
.C(n_143),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_218),
.C(n_182),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_165),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_229),
.B1(n_232),
.B2(n_236),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_212),
.A2(n_168),
.B1(n_151),
.B2(n_155),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_207),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_200),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_147),
.B1(n_163),
.B2(n_159),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_66),
.B1(n_164),
.B2(n_171),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_191),
.Y(n_237)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_171),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_197),
.Y(n_246)
);

INVx2_ASAP7_75t_R g241 ( 
.A(n_189),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_242),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_0),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_255),
.C(n_262),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_197),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_246),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_213),
.B1(n_204),
.B2(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_181),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_227),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_221),
.A2(n_195),
.B1(n_201),
.B2(n_196),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_222),
.B1(n_219),
.B2(n_235),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_238),
.B(n_211),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_251),
.A2(n_265),
.B(n_186),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_195),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_257),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_205),
.C(n_180),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_224),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_228),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_260),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_224),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_259),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_180),
.C(n_209),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_206),
.B1(n_188),
.B2(n_210),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_220),
.B1(n_240),
.B2(n_222),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_192),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_264),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_188),
.B(n_199),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_217),
.B(n_203),
.C(n_102),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_220),
.C(n_236),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_269),
.A2(n_253),
.B1(n_256),
.B2(n_0),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_266),
.C(n_250),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_280),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_234),
.B1(n_241),
.B2(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_261),
.B1(n_276),
.B2(n_258),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_234),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_222),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_255),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_219),
.B(n_225),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_262),
.B(n_252),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_246),
.B(n_233),
.CI(n_225),
.CON(n_283),
.SN(n_283)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_248),
.Y(n_289)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_233),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_7),
.B(n_2),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_265),
.B(n_263),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_288),
.A2(n_302),
.B(n_303),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_291),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_293),
.A2(n_271),
.B1(n_281),
.B2(n_282),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_298),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_295),
.B(n_297),
.Y(n_308)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_268),
.Y(n_296)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_301),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_249),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_272),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_9),
.B(n_3),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_278),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_316),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_309),
.A2(n_298),
.B1(n_275),
.B2(n_282),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_315),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_278),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_287),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_302),
.A2(n_285),
.B(n_267),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_317),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_267),
.C(n_292),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_324),
.C(n_315),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_305),
.B(n_270),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_326),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_321),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_292),
.C(n_280),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_307),
.A2(n_303),
.B1(n_288),
.B2(n_283),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_309),
.B1(n_304),
.B2(n_310),
.Y(n_333)
);

AO221x1_ASAP7_75t_L g326 ( 
.A1(n_312),
.A2(n_301),
.B1(n_277),
.B2(n_283),
.C(n_300),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_322),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_9),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_328),
.B(n_12),
.Y(n_336)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_329),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_314),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_331),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_313),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_332),
.A2(n_333),
.A3(n_321),
.B1(n_324),
.B2(n_323),
.C1(n_318),
.C2(n_11),
.Y(n_341)
);

AOI21x1_ASAP7_75t_L g334 ( 
.A1(n_326),
.A2(n_304),
.B(n_3),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_334),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_336),
.A2(n_337),
.B1(n_14),
.B2(n_6),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_341),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_337),
.A2(n_323),
.B1(n_6),
.B2(n_7),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_335),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_331),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_344),
.A2(n_346),
.B(n_347),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_333),
.Y(n_347)
);

AOI21xp33_ASAP7_75t_L g348 ( 
.A1(n_345),
.A2(n_340),
.B(n_342),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_348),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_349),
.B1(n_347),
.B2(n_12),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_10),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_12),
.Y(n_353)
);


endmodule